module ForwardingAgeLogic(
  input         clock,
  input         reset,
  input  [23:0] io_addr_matches,
  input  [4:0]  io_youngest_st_idx,
  output        io_forwarding_val,
  output [4:0]  io_forwarding_idx
);
  wire  _T = 5'h0 >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_0 = _T ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_1 = 5'h1 >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_1 = _T_1 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_2 = 5'h2 >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_2 = _T_2 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_3 = 5'h3 >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_3 = _T_3 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_4 = 5'h4 >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_4 = _T_4 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_5 = 5'h5 >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_5 = _T_5 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_6 = 5'h6 >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_6 = _T_6 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_7 = 5'h7 >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_7 = _T_7 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_8 = 5'h8 >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_8 = _T_8 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_9 = 5'h9 >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_9 = _T_9 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_10 = 5'ha >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_10 = _T_10 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_11 = 5'hb >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_11 = _T_11 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_12 = 5'hc >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_12 = _T_12 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_13 = 5'hd >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_13 = _T_13 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_14 = 5'he >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_14 = _T_14 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_15 = 5'hf >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_15 = _T_15 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_16 = 5'h10 >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_16 = _T_16 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_17 = 5'h11 >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_17 = _T_17 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_18 = 5'h12 >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_18 = _T_18 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_19 = 5'h13 >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_19 = _T_19 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_20 = 5'h14 >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_20 = _T_20 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_21 = 5'h15 >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_21 = _T_21 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_22 = 5'h16 >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_22 = _T_22 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire  _T_23 = 5'h17 >= io_youngest_st_idx; // @[lsu.scala 1763:17]
  wire  age_mask_23 = _T_23 ? 1'h0 : 1'h1; // @[lsu.scala 1764:7 lsu.scala 1765:22 lsu.scala 1762:19]
  wire [5:0] lo_lo = {age_mask_5,age_mask_4,age_mask_3,age_mask_2,age_mask_1,age_mask_0}; // @[lsu.scala 1771:46]
  wire [11:0] lo = {age_mask_11,age_mask_10,age_mask_9,age_mask_8,age_mask_7,age_mask_6,lo_lo}; // @[lsu.scala 1771:46]
  wire [5:0] hi_lo = {age_mask_17,age_mask_16,age_mask_15,age_mask_14,age_mask_13,age_mask_12}; // @[lsu.scala 1771:46]
  wire [23:0] _T_24 = {age_mask_23,age_mask_22,age_mask_21,age_mask_20,age_mask_19,age_mask_18,hi_lo,lo}; // @[lsu.scala 1771:46]
  wire [23:0] hi_1 = io_addr_matches & _T_24; // @[lsu.scala 1771:35]
  wire [47:0] matches_ = {hi_1,io_addr_matches}; // @[Cat.scala 30:58]
  wire [1:0] _GEN_29 = matches_[2] ? 2'h2 : {{1'd0}, matches_[1]}; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [1:0] _GEN_31 = matches_[3] ? 2'h3 : _GEN_29; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [2:0] _GEN_33 = matches_[4] ? 3'h4 : {{1'd0}, _GEN_31}; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [2:0] _GEN_35 = matches_[5] ? 3'h5 : _GEN_33; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [2:0] _GEN_37 = matches_[6] ? 3'h6 : _GEN_35; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [2:0] _GEN_39 = matches_[7] ? 3'h7 : _GEN_37; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [3:0] _GEN_41 = matches_[8] ? 4'h8 : {{1'd0}, _GEN_39}; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [3:0] _GEN_43 = matches_[9] ? 4'h9 : _GEN_41; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [3:0] _GEN_45 = matches_[10] ? 4'ha : _GEN_43; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [3:0] _GEN_47 = matches_[11] ? 4'hb : _GEN_45; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [3:0] _GEN_49 = matches_[12] ? 4'hc : _GEN_47; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [3:0] _GEN_51 = matches_[13] ? 4'hd : _GEN_49; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [3:0] _GEN_53 = matches_[14] ? 4'he : _GEN_51; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [3:0] _GEN_55 = matches_[15] ? 4'hf : _GEN_53; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_57 = matches_[16] ? 5'h10 : {{1'd0}, _GEN_55}; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_59 = matches_[17] ? 5'h11 : _GEN_57; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_61 = matches_[18] ? 5'h12 : _GEN_59; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_63 = matches_[19] ? 5'h13 : _GEN_61; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_65 = matches_[20] ? 5'h14 : _GEN_63; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_67 = matches_[21] ? 5'h15 : _GEN_65; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_69 = matches_[22] ? 5'h16 : _GEN_67; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_71 = matches_[23] ? 5'h17 : _GEN_69; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_73 = matches_[24] ? 5'h0 : _GEN_71; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_75 = matches_[25] ? 5'h1 : _GEN_73; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_77 = matches_[26] ? 5'h2 : _GEN_75; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_79 = matches_[27] ? 5'h3 : _GEN_77; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_81 = matches_[28] ? 5'h4 : _GEN_79; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_83 = matches_[29] ? 5'h5 : _GEN_81; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire  _GEN_84 = matches_[30] | (matches_[29] | (matches_[28] | (matches_[27] | (matches_[26] | (matches_[25] | (
    matches_[24] | (matches_[23] | (matches_[22] | (matches_[21] | (matches_[20] | (matches_[19] | (matches_[18] | (
    matches_[17] | (matches_[16] | (matches_[15] | (matches_[14] | (matches_[13] | (matches_[12] | (matches_[11] | (
    matches_[10] | (matches_[9] | (matches_[8] | (matches_[7] | (matches_[6] | (matches_[5] | (matches_[4] | (matches_[3
    ] | (matches_[2] | (matches_[1] | matches_[0]))))))))))))))))))))))))))))); // @[lsu.scala 1782:7 lsu.scala 1783:22]
  wire [4:0] _GEN_85 = matches_[30] ? 5'h6 : _GEN_83; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_87 = matches_[31] ? 5'h7 : _GEN_85; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_89 = matches_[32] ? 5'h8 : _GEN_87; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_91 = matches_[33] ? 5'h9 : _GEN_89; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_93 = matches_[34] ? 5'ha : _GEN_91; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_95 = matches_[35] ? 5'hb : _GEN_93; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_97 = matches_[36] ? 5'hc : _GEN_95; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_99 = matches_[37] ? 5'hd : _GEN_97; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_101 = matches_[38] ? 5'he : _GEN_99; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_103 = matches_[39] ? 5'hf : _GEN_101; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_105 = matches_[40] ? 5'h10 : _GEN_103; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_107 = matches_[41] ? 5'h11 : _GEN_105; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_109 = matches_[42] ? 5'h12 : _GEN_107; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_111 = matches_[43] ? 5'h13 : _GEN_109; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_113 = matches_[44] ? 5'h14 : _GEN_111; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_115 = matches_[45] ? 5'h15 : _GEN_113; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  wire [4:0] _GEN_117 = matches_[46] ? 5'h16 : _GEN_115; // @[lsu.scala 1782:7 lsu.scala 1784:28]
  assign io_forwarding_val = matches_[47] | (matches_[46] | (matches_[45] | (matches_[44] | (matches_[43] | (matches_[42
    ] | (matches_[41] | (matches_[40] | (matches_[39] | (matches_[38] | (matches_[37] | (matches_[36] | (matches_[35] |
    (matches_[34] | (matches_[33] | (matches_[32] | (matches_[31] | _GEN_84)))))))))))))))); // @[lsu.scala 1782:7 lsu.scala 1783:22]
  assign io_forwarding_idx = matches_[47] ? 5'h17 : _GEN_117; // @[lsu.scala 1782:7 lsu.scala 1784:28]
endmodule
