module BundleBridgeNexus(
  input   clock,
  input   reset
);
endmodule
