module RenameMapTable(
  input         clock,
  input         reset,
  input  [5:0]  io_map_reqs_0_lrs1,
  input  [5:0]  io_map_reqs_0_lrs2,
  input  [5:0]  io_map_reqs_0_lrs3,
  input  [5:0]  io_map_reqs_0_ldst,
  input  [5:0]  io_map_reqs_1_lrs1,
  input  [5:0]  io_map_reqs_1_lrs2,
  input  [5:0]  io_map_reqs_1_lrs3,
  input  [5:0]  io_map_reqs_1_ldst,
  output        io_map_resps_0_prs1_valid,
  output [5:0]  io_map_resps_0_prs1_bits,
  output        io_map_resps_0_prs2_valid,
  output [5:0]  io_map_resps_0_prs2_bits,
  output        io_map_resps_0_prs3_valid,
  output [5:0]  io_map_resps_0_prs3_bits,
  output        io_map_resps_0_stale_pdst_valid,
  output [5:0]  io_map_resps_0_stale_pdst_bits,
  output        io_map_resps_1_prs1_valid,
  output [5:0]  io_map_resps_1_prs1_bits,
  output        io_map_resps_1_prs2_valid,
  output [5:0]  io_map_resps_1_prs2_bits,
  output        io_map_resps_1_prs3_valid,
  output [5:0]  io_map_resps_1_prs3_bits,
  output        io_map_resps_1_stale_pdst_valid,
  output [5:0]  io_map_resps_1_stale_pdst_bits,
  input  [5:0]  io_remap_reqs_0_ldst,
  input  [5:0]  io_remap_reqs_0_pdst,
  input         io_remap_reqs_0_valid,
  input  [5:0]  io_remap_reqs_1_ldst,
  input  [5:0]  io_remap_reqs_1_pdst,
  input         io_remap_reqs_1_valid,
  input         io_ren_br_tags_0_valid,
  input  [3:0]  io_ren_br_tags_0_bits,
  input         io_ren_br_tags_1_valid,
  input  [3:0]  io_ren_br_tags_1_bits,
  input  [11:0] io_brupdate_b1_resolve_mask,
  input  [11:0] io_brupdate_b1_mispredict_mask,
  input  [6:0]  io_brupdate_b2_uop_uopc,
  input  [31:0] io_brupdate_b2_uop_inst,
  input  [31:0] io_brupdate_b2_uop_debug_inst,
  input         io_brupdate_b2_uop_is_rvc,
  input  [39:0] io_brupdate_b2_uop_debug_pc,
  input  [2:0]  io_brupdate_b2_uop_iq_type,
  input  [9:0]  io_brupdate_b2_uop_fu_code,
  input  [3:0]  io_brupdate_b2_uop_ctrl_br_type,
  input  [1:0]  io_brupdate_b2_uop_ctrl_op1_sel,
  input  [2:0]  io_brupdate_b2_uop_ctrl_op2_sel,
  input  [2:0]  io_brupdate_b2_uop_ctrl_imm_sel,
  input  [3:0]  io_brupdate_b2_uop_ctrl_op_fcn,
  input         io_brupdate_b2_uop_ctrl_fcn_dw,
  input  [2:0]  io_brupdate_b2_uop_ctrl_csr_cmd,
  input         io_brupdate_b2_uop_ctrl_is_load,
  input         io_brupdate_b2_uop_ctrl_is_sta,
  input         io_brupdate_b2_uop_ctrl_is_std,
  input  [1:0]  io_brupdate_b2_uop_iw_state,
  input         io_brupdate_b2_uop_iw_p1_poisoned,
  input         io_brupdate_b2_uop_iw_p2_poisoned,
  input         io_brupdate_b2_uop_is_br,
  input         io_brupdate_b2_uop_is_jalr,
  input         io_brupdate_b2_uop_is_jal,
  input         io_brupdate_b2_uop_is_sfb,
  input  [11:0] io_brupdate_b2_uop_br_mask,
  input  [3:0]  io_brupdate_b2_uop_br_tag,
  input  [4:0]  io_brupdate_b2_uop_ftq_idx,
  input         io_brupdate_b2_uop_edge_inst,
  input  [5:0]  io_brupdate_b2_uop_pc_lob,
  input         io_brupdate_b2_uop_taken,
  input  [19:0] io_brupdate_b2_uop_imm_packed,
  input  [11:0] io_brupdate_b2_uop_csr_addr,
  input  [5:0]  io_brupdate_b2_uop_rob_idx,
  input  [3:0]  io_brupdate_b2_uop_ldq_idx,
  input  [3:0]  io_brupdate_b2_uop_stq_idx,
  input  [1:0]  io_brupdate_b2_uop_rxq_idx,
  input  [5:0]  io_brupdate_b2_uop_pdst,
  input  [5:0]  io_brupdate_b2_uop_prs1,
  input  [5:0]  io_brupdate_b2_uop_prs2,
  input  [5:0]  io_brupdate_b2_uop_prs3,
  input  [4:0]  io_brupdate_b2_uop_ppred,
  input         io_brupdate_b2_uop_prs1_busy,
  input         io_brupdate_b2_uop_prs2_busy,
  input         io_brupdate_b2_uop_prs3_busy,
  input         io_brupdate_b2_uop_ppred_busy,
  input  [5:0]  io_brupdate_b2_uop_stale_pdst,
  input         io_brupdate_b2_uop_exception,
  input  [63:0] io_brupdate_b2_uop_exc_cause,
  input         io_brupdate_b2_uop_bypassable,
  input  [4:0]  io_brupdate_b2_uop_mem_cmd,
  input  [1:0]  io_brupdate_b2_uop_mem_size,
  input         io_brupdate_b2_uop_mem_signed,
  input         io_brupdate_b2_uop_is_fence,
  input         io_brupdate_b2_uop_is_fencei,
  input         io_brupdate_b2_uop_is_amo,
  input         io_brupdate_b2_uop_uses_ldq,
  input         io_brupdate_b2_uop_uses_stq,
  input         io_brupdate_b2_uop_is_sys_pc2epc,
  input         io_brupdate_b2_uop_is_unique,
  input         io_brupdate_b2_uop_flush_on_commit,
  input         io_brupdate_b2_uop_ldst_is_rs1,
  input  [5:0]  io_brupdate_b2_uop_ldst,
  input  [5:0]  io_brupdate_b2_uop_lrs1,
  input  [5:0]  io_brupdate_b2_uop_lrs2,
  input  [5:0]  io_brupdate_b2_uop_lrs3,
  input         io_brupdate_b2_uop_ldst_val,
  input  [1:0]  io_brupdate_b2_uop_dst_rtype,
  input  [1:0]  io_brupdate_b2_uop_lrs1_rtype,
  input  [1:0]  io_brupdate_b2_uop_lrs2_rtype,
  input         io_brupdate_b2_uop_frs3_en,
  input         io_brupdate_b2_uop_fp_val,
  input         io_brupdate_b2_uop_fp_single,
  input         io_brupdate_b2_uop_xcpt_pf_if,
  input         io_brupdate_b2_uop_xcpt_ae_if,
  input         io_brupdate_b2_uop_xcpt_ma_if,
  input         io_brupdate_b2_uop_bp_debug_if,
  input         io_brupdate_b2_uop_bp_xcpt_if,
  input  [1:0]  io_brupdate_b2_uop_debug_fsrc,
  input  [1:0]  io_brupdate_b2_uop_debug_tsrc,
  input         io_brupdate_b2_valid,
  input         io_brupdate_b2_mispredict,
  input         io_brupdate_b2_taken,
  input  [2:0]  io_brupdate_b2_cfi_type,
  input  [1:0]  io_brupdate_b2_pc_sel,
  input  [39:0] io_brupdate_b2_jalr_target,
  input  [20:0] io_brupdate_b2_target_offset,
  input         io_rollback,
  input  [5:0]  io_commit_regs_0_ldst,
  input  [5:0]  io_commit_regs_0_pdst,
  input         io_commit_regs_0_valid,
  input  [5:0]  io_commit_regs_1_ldst,
  input  [5:0]  io_commit_regs_1_pdst,
  input         io_commit_regs_1_valid,
  input         io_flush,
  output [63:0] io_commit_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
`endif // RANDOMIZE_REG_INIT
  reg [5:0] map_table_0; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_1; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_2; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_3; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_4; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_5; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_6; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_7; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_8; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_9; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_10; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_11; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_12; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_13; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_14; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_15; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_16; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_17; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_18; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_19; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_20; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_21; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_22; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_23; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_24; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_25; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_26; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_27; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_28; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_29; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_30; // @[rename-maptable.scala 77:26]
  reg [5:0] map_table_31; // @[rename-maptable.scala 77:26]
  reg [5:0] commit_map_table_0; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_1; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_2; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_3; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_4; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_5; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_6; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_7; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_8; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_9; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_10; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_11; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_12; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_13; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_14; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_15; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_16; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_17; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_18; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_19; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_20; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_21; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_22; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_23; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_24; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_25; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_26; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_27; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_28; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_29; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_30; // @[rename-maptable.scala 78:33]
  reg [5:0] commit_map_table_31; // @[rename-maptable.scala 78:33]
  reg [5:0] br_snapshots_0_1; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_2; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_3; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_4; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_5; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_6; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_7; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_8; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_9; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_10; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_11; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_12; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_13; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_14; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_15; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_16; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_17; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_18; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_19; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_20; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_21; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_22; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_23; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_24; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_25; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_26; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_27; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_28; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_29; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_30; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_0_31; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_1; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_2; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_3; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_4; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_5; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_6; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_7; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_8; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_9; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_10; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_11; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_12; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_13; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_14; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_15; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_16; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_17; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_18; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_19; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_20; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_21; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_22; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_23; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_24; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_25; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_26; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_27; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_28; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_29; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_30; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_1_31; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_1; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_2; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_3; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_4; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_5; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_6; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_7; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_8; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_9; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_10; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_11; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_12; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_13; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_14; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_15; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_16; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_17; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_18; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_19; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_20; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_21; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_22; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_23; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_24; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_25; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_26; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_27; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_28; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_29; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_30; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_2_31; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_1; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_2; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_3; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_4; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_5; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_6; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_7; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_8; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_9; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_10; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_11; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_12; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_13; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_14; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_15; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_16; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_17; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_18; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_19; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_20; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_21; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_22; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_23; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_24; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_25; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_26; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_27; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_28; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_29; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_30; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_3_31; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_1; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_2; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_3; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_4; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_5; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_6; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_7; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_8; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_9; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_10; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_11; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_12; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_13; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_14; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_15; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_16; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_17; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_18; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_19; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_20; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_21; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_22; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_23; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_24; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_25; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_26; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_27; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_28; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_29; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_30; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_4_31; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_1; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_2; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_3; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_4; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_5; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_6; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_7; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_8; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_9; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_10; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_11; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_12; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_13; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_14; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_15; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_16; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_17; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_18; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_19; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_20; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_21; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_22; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_23; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_24; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_25; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_26; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_27; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_28; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_29; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_30; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_5_31; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_1; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_2; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_3; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_4; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_5; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_6; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_7; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_8; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_9; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_10; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_11; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_12; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_13; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_14; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_15; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_16; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_17; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_18; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_19; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_20; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_21; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_22; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_23; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_24; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_25; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_26; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_27; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_28; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_29; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_30; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_6_31; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_1; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_2; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_3; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_4; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_5; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_6; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_7; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_8; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_9; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_10; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_11; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_12; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_13; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_14; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_15; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_16; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_17; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_18; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_19; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_20; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_21; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_22; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_23; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_24; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_25; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_26; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_27; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_28; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_29; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_30; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_7_31; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_1; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_2; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_3; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_4; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_5; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_6; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_7; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_8; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_9; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_10; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_11; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_12; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_13; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_14; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_15; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_16; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_17; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_18; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_19; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_20; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_21; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_22; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_23; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_24; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_25; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_26; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_27; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_28; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_29; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_30; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_8_31; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_1; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_2; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_3; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_4; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_5; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_6; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_7; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_8; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_9; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_10; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_11; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_12; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_13; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_14; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_15; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_16; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_17; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_18; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_19; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_20; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_21; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_22; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_23; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_24; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_25; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_26; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_27; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_28; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_29; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_30; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_9_31; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_1; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_2; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_3; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_4; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_5; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_6; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_7; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_8; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_9; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_10; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_11; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_12; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_13; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_14; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_15; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_16; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_17; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_18; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_19; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_20; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_21; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_22; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_23; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_24; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_25; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_26; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_27; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_28; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_29; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_30; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_10_31; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_1; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_2; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_3; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_4; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_5; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_6; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_7; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_8; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_9; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_10; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_11; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_12; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_13; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_14; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_15; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_16; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_17; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_18; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_19; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_20; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_21; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_22; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_23; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_24; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_25; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_26; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_27; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_28; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_29; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_30; // @[rename-maptable.scala 79:25]
  reg [5:0] br_snapshots_11_31; // @[rename-maptable.scala 79:25]
  wire [63:0] _T = 64'h1 << io_remap_reqs_0_ldst; // @[OneHot.scala 58:35]
  wire [31:0] _T_2 = io_remap_reqs_0_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _GEN_2624 = {{32'd0}, _T_2}; // @[rename-maptable.scala 86:69]
  wire [63:0] remap_ldsts_oh_0 = _T & _GEN_2624; // @[rename-maptable.scala 86:69]
  wire [63:0] _T_3 = 64'h1 << io_remap_reqs_1_ldst; // @[OneHot.scala 58:35]
  wire [31:0] _T_5 = io_remap_reqs_1_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _GEN_2625 = {{32'd0}, _T_5}; // @[rename-maptable.scala 86:69]
  wire [63:0] remap_ldsts_oh_1 = _T_3 & _GEN_2625; // @[rename-maptable.scala 86:69]
  wire [63:0] _T_6 = 64'h1 << io_commit_regs_0_ldst; // @[OneHot.scala 58:35]
  wire [31:0] _T_8 = io_commit_regs_0_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _GEN_2626 = {{32'd0}, _T_8}; // @[rename-maptable.scala 89:69]
  wire [63:0] rrat_ldsts_oh_0 = _T_6 & _GEN_2626; // @[rename-maptable.scala 89:69]
  wire [63:0] _T_9 = 64'h1 << io_commit_regs_1_ldst; // @[OneHot.scala 58:35]
  wire [31:0] _T_11 = io_commit_regs_1_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _GEN_2627 = {{32'd0}, _T_11}; // @[rename-maptable.scala 89:69]
  wire [63:0] rrat_ldsts_oh_1 = _T_9 & _GEN_2627; // @[rename-maptable.scala 89:69]
  wire [5:0] _T_14 = rrat_ldsts_oh_0[0] ? io_commit_regs_0_pdst : commit_map_table_0; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_0 = rrat_ldsts_oh_1[0] ? io_commit_regs_1_pdst : _T_14; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_18 = rrat_ldsts_oh_0[1] ? io_commit_regs_0_pdst : commit_map_table_1; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_1 = rrat_ldsts_oh_1[1] ? io_commit_regs_1_pdst : _T_18; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_22 = rrat_ldsts_oh_0[2] ? io_commit_regs_0_pdst : commit_map_table_2; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_2 = rrat_ldsts_oh_1[2] ? io_commit_regs_1_pdst : _T_22; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_26 = rrat_ldsts_oh_0[3] ? io_commit_regs_0_pdst : commit_map_table_3; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_3 = rrat_ldsts_oh_1[3] ? io_commit_regs_1_pdst : _T_26; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_30 = rrat_ldsts_oh_0[4] ? io_commit_regs_0_pdst : commit_map_table_4; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_4 = rrat_ldsts_oh_1[4] ? io_commit_regs_1_pdst : _T_30; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_34 = rrat_ldsts_oh_0[5] ? io_commit_regs_0_pdst : commit_map_table_5; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_5 = rrat_ldsts_oh_1[5] ? io_commit_regs_1_pdst : _T_34; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_38 = rrat_ldsts_oh_0[6] ? io_commit_regs_0_pdst : commit_map_table_6; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_6 = rrat_ldsts_oh_1[6] ? io_commit_regs_1_pdst : _T_38; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_42 = rrat_ldsts_oh_0[7] ? io_commit_regs_0_pdst : commit_map_table_7; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_7 = rrat_ldsts_oh_1[7] ? io_commit_regs_1_pdst : _T_42; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_46 = rrat_ldsts_oh_0[8] ? io_commit_regs_0_pdst : commit_map_table_8; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_8 = rrat_ldsts_oh_1[8] ? io_commit_regs_1_pdst : _T_46; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_50 = rrat_ldsts_oh_0[9] ? io_commit_regs_0_pdst : commit_map_table_9; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_9 = rrat_ldsts_oh_1[9] ? io_commit_regs_1_pdst : _T_50; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_54 = rrat_ldsts_oh_0[10] ? io_commit_regs_0_pdst : commit_map_table_10; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_10 = rrat_ldsts_oh_1[10] ? io_commit_regs_1_pdst : _T_54; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_58 = rrat_ldsts_oh_0[11] ? io_commit_regs_0_pdst : commit_map_table_11; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_11 = rrat_ldsts_oh_1[11] ? io_commit_regs_1_pdst : _T_58; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_62 = rrat_ldsts_oh_0[12] ? io_commit_regs_0_pdst : commit_map_table_12; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_12 = rrat_ldsts_oh_1[12] ? io_commit_regs_1_pdst : _T_62; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_66 = rrat_ldsts_oh_0[13] ? io_commit_regs_0_pdst : commit_map_table_13; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_13 = rrat_ldsts_oh_1[13] ? io_commit_regs_1_pdst : _T_66; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_70 = rrat_ldsts_oh_0[14] ? io_commit_regs_0_pdst : commit_map_table_14; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_14 = rrat_ldsts_oh_1[14] ? io_commit_regs_1_pdst : _T_70; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_74 = rrat_ldsts_oh_0[15] ? io_commit_regs_0_pdst : commit_map_table_15; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_15 = rrat_ldsts_oh_1[15] ? io_commit_regs_1_pdst : _T_74; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_78 = rrat_ldsts_oh_0[16] ? io_commit_regs_0_pdst : commit_map_table_16; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_16 = rrat_ldsts_oh_1[16] ? io_commit_regs_1_pdst : _T_78; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_82 = rrat_ldsts_oh_0[17] ? io_commit_regs_0_pdst : commit_map_table_17; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_17 = rrat_ldsts_oh_1[17] ? io_commit_regs_1_pdst : _T_82; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_86 = rrat_ldsts_oh_0[18] ? io_commit_regs_0_pdst : commit_map_table_18; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_18 = rrat_ldsts_oh_1[18] ? io_commit_regs_1_pdst : _T_86; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_90 = rrat_ldsts_oh_0[19] ? io_commit_regs_0_pdst : commit_map_table_19; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_19 = rrat_ldsts_oh_1[19] ? io_commit_regs_1_pdst : _T_90; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_94 = rrat_ldsts_oh_0[20] ? io_commit_regs_0_pdst : commit_map_table_20; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_20 = rrat_ldsts_oh_1[20] ? io_commit_regs_1_pdst : _T_94; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_98 = rrat_ldsts_oh_0[21] ? io_commit_regs_0_pdst : commit_map_table_21; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_21 = rrat_ldsts_oh_1[21] ? io_commit_regs_1_pdst : _T_98; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_102 = rrat_ldsts_oh_0[22] ? io_commit_regs_0_pdst : commit_map_table_22; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_22 = rrat_ldsts_oh_1[22] ? io_commit_regs_1_pdst : _T_102; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_106 = rrat_ldsts_oh_0[23] ? io_commit_regs_0_pdst : commit_map_table_23; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_23 = rrat_ldsts_oh_1[23] ? io_commit_regs_1_pdst : _T_106; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_110 = rrat_ldsts_oh_0[24] ? io_commit_regs_0_pdst : commit_map_table_24; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_24 = rrat_ldsts_oh_1[24] ? io_commit_regs_1_pdst : _T_110; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_114 = rrat_ldsts_oh_0[25] ? io_commit_regs_0_pdst : commit_map_table_25; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_25 = rrat_ldsts_oh_1[25] ? io_commit_regs_1_pdst : _T_114; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_118 = rrat_ldsts_oh_0[26] ? io_commit_regs_0_pdst : commit_map_table_26; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_26 = rrat_ldsts_oh_1[26] ? io_commit_regs_1_pdst : _T_118; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_122 = rrat_ldsts_oh_0[27] ? io_commit_regs_0_pdst : commit_map_table_27; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_27 = rrat_ldsts_oh_1[27] ? io_commit_regs_1_pdst : _T_122; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_126 = rrat_ldsts_oh_0[28] ? io_commit_regs_0_pdst : commit_map_table_28; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_28 = rrat_ldsts_oh_1[28] ? io_commit_regs_1_pdst : _T_126; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_130 = rrat_ldsts_oh_0[29] ? io_commit_regs_0_pdst : commit_map_table_29; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_29 = rrat_ldsts_oh_1[29] ? io_commit_regs_1_pdst : _T_130; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_134 = rrat_ldsts_oh_0[30] ? io_commit_regs_0_pdst : commit_map_table_30; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_30 = rrat_ldsts_oh_1[30] ? io_commit_regs_1_pdst : _T_134; // @[rename-maptable.scala 95:75]
  wire [5:0] _T_138 = rrat_ldsts_oh_0[31] ? io_commit_regs_0_pdst : commit_map_table_31; // @[rename-maptable.scala 95:75]
  wire [5:0] t_commit_map_table_31 = rrat_ldsts_oh_1[31] ? io_commit_regs_1_pdst : _T_138; // @[rename-maptable.scala 95:75]
  wire [63:0] _T_266 = 64'h1 << t_commit_map_table_0; // @[OneHot.scala 58:35]
  wire [63:0] _T_269 = 64'h1 << t_commit_map_table_1; // @[OneHot.scala 58:35]
  wire [63:0] _T_272 = 64'h1 << t_commit_map_table_2; // @[OneHot.scala 58:35]
  wire [63:0] _T_275 = 64'h1 << t_commit_map_table_3; // @[OneHot.scala 58:35]
  wire [63:0] _T_278 = 64'h1 << t_commit_map_table_4; // @[OneHot.scala 58:35]
  wire [63:0] _T_281 = 64'h1 << t_commit_map_table_5; // @[OneHot.scala 58:35]
  wire [63:0] _T_284 = 64'h1 << t_commit_map_table_6; // @[OneHot.scala 58:35]
  wire [63:0] _T_287 = 64'h1 << t_commit_map_table_7; // @[OneHot.scala 58:35]
  wire [63:0] _T_290 = 64'h1 << t_commit_map_table_8; // @[OneHot.scala 58:35]
  wire [63:0] _T_293 = 64'h1 << t_commit_map_table_9; // @[OneHot.scala 58:35]
  wire [63:0] _T_296 = 64'h1 << t_commit_map_table_10; // @[OneHot.scala 58:35]
  wire [63:0] _T_299 = 64'h1 << t_commit_map_table_11; // @[OneHot.scala 58:35]
  wire [63:0] _T_302 = 64'h1 << t_commit_map_table_12; // @[OneHot.scala 58:35]
  wire [63:0] _T_305 = 64'h1 << t_commit_map_table_13; // @[OneHot.scala 58:35]
  wire [63:0] _T_308 = 64'h1 << t_commit_map_table_14; // @[OneHot.scala 58:35]
  wire [63:0] _T_311 = 64'h1 << t_commit_map_table_15; // @[OneHot.scala 58:35]
  wire [63:0] _T_314 = 64'h1 << t_commit_map_table_16; // @[OneHot.scala 58:35]
  wire [63:0] _T_317 = 64'h1 << t_commit_map_table_17; // @[OneHot.scala 58:35]
  wire [63:0] _T_320 = 64'h1 << t_commit_map_table_18; // @[OneHot.scala 58:35]
  wire [63:0] _T_323 = 64'h1 << t_commit_map_table_19; // @[OneHot.scala 58:35]
  wire [63:0] _T_326 = 64'h1 << t_commit_map_table_20; // @[OneHot.scala 58:35]
  wire [63:0] _T_329 = 64'h1 << t_commit_map_table_21; // @[OneHot.scala 58:35]
  wire [63:0] _T_332 = 64'h1 << t_commit_map_table_22; // @[OneHot.scala 58:35]
  wire [63:0] _T_335 = 64'h1 << t_commit_map_table_23; // @[OneHot.scala 58:35]
  wire [63:0] _T_338 = 64'h1 << t_commit_map_table_24; // @[OneHot.scala 58:35]
  wire [63:0] _T_341 = 64'h1 << t_commit_map_table_25; // @[OneHot.scala 58:35]
  wire [63:0] _T_344 = 64'h1 << t_commit_map_table_26; // @[OneHot.scala 58:35]
  wire [63:0] _T_347 = 64'h1 << t_commit_map_table_27; // @[OneHot.scala 58:35]
  wire [63:0] _T_350 = 64'h1 << t_commit_map_table_28; // @[OneHot.scala 58:35]
  wire [63:0] _T_353 = 64'h1 << t_commit_map_table_29; // @[OneHot.scala 58:35]
  wire [63:0] _T_356 = 64'h1 << t_commit_map_table_30; // @[OneHot.scala 58:35]
  wire [63:0] _T_359 = 64'h1 << t_commit_map_table_31; // @[OneHot.scala 58:35]
  wire [63:0] _T_362 = _T_266 | _T_269; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_363 = _T_362 | _T_272; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_364 = _T_363 | _T_275; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_365 = _T_364 | _T_278; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_366 = _T_365 | _T_281; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_367 = _T_366 | _T_284; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_368 = _T_367 | _T_287; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_369 = _T_368 | _T_290; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_370 = _T_369 | _T_293; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_371 = _T_370 | _T_296; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_372 = _T_371 | _T_299; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_373 = _T_372 | _T_302; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_374 = _T_373 | _T_305; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_375 = _T_374 | _T_308; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_376 = _T_375 | _T_311; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_377 = _T_376 | _T_314; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_378 = _T_377 | _T_317; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_379 = _T_378 | _T_320; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_380 = _T_379 | _T_323; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_381 = _T_380 | _T_326; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_382 = _T_381 | _T_329; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_383 = _T_382 | _T_332; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_384 = _T_383 | _T_335; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_385 = _T_384 | _T_338; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_386 = _T_385 | _T_341; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_387 = _T_386 | _T_344; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_388 = _T_387 | _T_347; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_389 = _T_388 | _T_350; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_390 = _T_389 | _T_353; // @[rename-maptable.scala 112:104]
  wire [63:0] _T_391 = _T_390 | _T_356; // @[rename-maptable.scala 112:104]
  wire [5:0] remap_table_1_1 = remap_ldsts_oh_0[1] ? io_remap_reqs_0_pdst : map_table_1; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_2 = remap_ldsts_oh_0[2] ? io_remap_reqs_0_pdst : map_table_2; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_3 = remap_ldsts_oh_0[3] ? io_remap_reqs_0_pdst : map_table_3; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_4 = remap_ldsts_oh_0[4] ? io_remap_reqs_0_pdst : map_table_4; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_5 = remap_ldsts_oh_0[5] ? io_remap_reqs_0_pdst : map_table_5; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_6 = remap_ldsts_oh_0[6] ? io_remap_reqs_0_pdst : map_table_6; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_7 = remap_ldsts_oh_0[7] ? io_remap_reqs_0_pdst : map_table_7; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_8 = remap_ldsts_oh_0[8] ? io_remap_reqs_0_pdst : map_table_8; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_9 = remap_ldsts_oh_0[9] ? io_remap_reqs_0_pdst : map_table_9; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_10 = remap_ldsts_oh_0[10] ? io_remap_reqs_0_pdst : map_table_10; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_11 = remap_ldsts_oh_0[11] ? io_remap_reqs_0_pdst : map_table_11; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_12 = remap_ldsts_oh_0[12] ? io_remap_reqs_0_pdst : map_table_12; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_13 = remap_ldsts_oh_0[13] ? io_remap_reqs_0_pdst : map_table_13; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_14 = remap_ldsts_oh_0[14] ? io_remap_reqs_0_pdst : map_table_14; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_15 = remap_ldsts_oh_0[15] ? io_remap_reqs_0_pdst : map_table_15; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_16 = remap_ldsts_oh_0[16] ? io_remap_reqs_0_pdst : map_table_16; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_17 = remap_ldsts_oh_0[17] ? io_remap_reqs_0_pdst : map_table_17; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_18 = remap_ldsts_oh_0[18] ? io_remap_reqs_0_pdst : map_table_18; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_19 = remap_ldsts_oh_0[19] ? io_remap_reqs_0_pdst : map_table_19; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_20 = remap_ldsts_oh_0[20] ? io_remap_reqs_0_pdst : map_table_20; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_21 = remap_ldsts_oh_0[21] ? io_remap_reqs_0_pdst : map_table_21; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_22 = remap_ldsts_oh_0[22] ? io_remap_reqs_0_pdst : map_table_22; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_23 = remap_ldsts_oh_0[23] ? io_remap_reqs_0_pdst : map_table_23; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_24 = remap_ldsts_oh_0[24] ? io_remap_reqs_0_pdst : map_table_24; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_25 = remap_ldsts_oh_0[25] ? io_remap_reqs_0_pdst : map_table_25; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_26 = remap_ldsts_oh_0[26] ? io_remap_reqs_0_pdst : map_table_26; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_27 = remap_ldsts_oh_0[27] ? io_remap_reqs_0_pdst : map_table_27; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_28 = remap_ldsts_oh_0[28] ? io_remap_reqs_0_pdst : map_table_28; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_29 = remap_ldsts_oh_0[29] ? io_remap_reqs_0_pdst : map_table_29; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_30 = remap_ldsts_oh_0[30] ? io_remap_reqs_0_pdst : map_table_30; // @[rename-maptable.scala 122:70]
  wire [5:0] remap_table_1_31 = remap_ldsts_oh_0[31] ? io_remap_reqs_0_pdst : map_table_31; // @[rename-maptable.scala 122:70]
  wire [5:0] _GEN_12 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_1 : br_snapshots_0_1; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_13 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_1 : br_snapshots_1_1; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_14 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_1 : br_snapshots_2_1; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_15 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_1 : br_snapshots_3_1; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_16 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_1 : br_snapshots_4_1; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_17 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_1 : br_snapshots_5_1; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_18 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_1 : br_snapshots_6_1; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_19 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_1 : br_snapshots_7_1; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_20 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_1 : br_snapshots_8_1; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_21 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_1 : br_snapshots_9_1; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_22 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_1 : br_snapshots_10_1; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_23 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_1 : br_snapshots_11_1; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_24 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_2 : br_snapshots_0_2; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_25 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_2 : br_snapshots_1_2; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_26 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_2 : br_snapshots_2_2; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_27 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_2 : br_snapshots_3_2; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_28 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_2 : br_snapshots_4_2; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_29 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_2 : br_snapshots_5_2; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_30 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_2 : br_snapshots_6_2; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_31 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_2 : br_snapshots_7_2; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_32 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_2 : br_snapshots_8_2; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_33 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_2 : br_snapshots_9_2; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_34 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_2 : br_snapshots_10_2; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_35 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_2 : br_snapshots_11_2; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_36 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_3 : br_snapshots_0_3; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_37 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_3 : br_snapshots_1_3; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_38 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_3 : br_snapshots_2_3; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_39 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_3 : br_snapshots_3_3; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_40 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_3 : br_snapshots_4_3; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_41 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_3 : br_snapshots_5_3; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_42 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_3 : br_snapshots_6_3; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_43 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_3 : br_snapshots_7_3; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_44 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_3 : br_snapshots_8_3; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_45 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_3 : br_snapshots_9_3; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_46 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_3 : br_snapshots_10_3; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_47 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_3 : br_snapshots_11_3; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_48 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_4 : br_snapshots_0_4; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_49 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_4 : br_snapshots_1_4; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_50 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_4 : br_snapshots_2_4; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_51 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_4 : br_snapshots_3_4; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_52 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_4 : br_snapshots_4_4; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_53 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_4 : br_snapshots_5_4; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_54 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_4 : br_snapshots_6_4; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_55 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_4 : br_snapshots_7_4; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_56 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_4 : br_snapshots_8_4; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_57 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_4 : br_snapshots_9_4; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_58 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_4 : br_snapshots_10_4; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_59 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_4 : br_snapshots_11_4; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_60 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_5 : br_snapshots_0_5; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_61 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_5 : br_snapshots_1_5; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_62 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_5 : br_snapshots_2_5; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_63 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_5 : br_snapshots_3_5; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_64 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_5 : br_snapshots_4_5; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_65 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_5 : br_snapshots_5_5; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_66 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_5 : br_snapshots_6_5; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_67 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_5 : br_snapshots_7_5; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_68 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_5 : br_snapshots_8_5; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_69 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_5 : br_snapshots_9_5; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_70 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_5 : br_snapshots_10_5; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_71 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_5 : br_snapshots_11_5; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_72 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_6 : br_snapshots_0_6; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_73 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_6 : br_snapshots_1_6; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_74 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_6 : br_snapshots_2_6; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_75 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_6 : br_snapshots_3_6; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_76 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_6 : br_snapshots_4_6; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_77 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_6 : br_snapshots_5_6; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_78 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_6 : br_snapshots_6_6; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_79 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_6 : br_snapshots_7_6; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_80 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_6 : br_snapshots_8_6; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_81 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_6 : br_snapshots_9_6; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_82 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_6 : br_snapshots_10_6; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_83 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_6 : br_snapshots_11_6; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_84 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_7 : br_snapshots_0_7; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_85 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_7 : br_snapshots_1_7; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_86 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_7 : br_snapshots_2_7; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_87 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_7 : br_snapshots_3_7; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_88 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_7 : br_snapshots_4_7; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_89 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_7 : br_snapshots_5_7; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_90 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_7 : br_snapshots_6_7; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_91 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_7 : br_snapshots_7_7; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_92 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_7 : br_snapshots_8_7; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_93 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_7 : br_snapshots_9_7; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_94 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_7 : br_snapshots_10_7; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_95 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_7 : br_snapshots_11_7; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_96 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_8 : br_snapshots_0_8; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_97 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_8 : br_snapshots_1_8; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_98 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_8 : br_snapshots_2_8; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_99 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_8 : br_snapshots_3_8; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_100 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_8 : br_snapshots_4_8; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_101 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_8 : br_snapshots_5_8; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_102 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_8 : br_snapshots_6_8; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_103 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_8 : br_snapshots_7_8; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_104 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_8 : br_snapshots_8_8; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_105 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_8 : br_snapshots_9_8; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_106 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_8 : br_snapshots_10_8; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_107 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_8 : br_snapshots_11_8; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_108 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_9 : br_snapshots_0_9; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_109 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_9 : br_snapshots_1_9; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_110 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_9 : br_snapshots_2_9; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_111 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_9 : br_snapshots_3_9; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_112 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_9 : br_snapshots_4_9; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_113 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_9 : br_snapshots_5_9; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_114 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_9 : br_snapshots_6_9; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_115 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_9 : br_snapshots_7_9; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_116 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_9 : br_snapshots_8_9; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_117 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_9 : br_snapshots_9_9; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_118 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_9 : br_snapshots_10_9; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_119 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_9 : br_snapshots_11_9; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_120 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_10 : br_snapshots_0_10; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_121 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_10 : br_snapshots_1_10; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_122 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_10 : br_snapshots_2_10; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_123 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_10 : br_snapshots_3_10; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_124 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_10 : br_snapshots_4_10; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_125 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_10 : br_snapshots_5_10; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_126 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_10 : br_snapshots_6_10; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_127 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_10 : br_snapshots_7_10; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_128 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_10 : br_snapshots_8_10; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_129 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_10 : br_snapshots_9_10; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_130 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_10 : br_snapshots_10_10; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_131 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_10 : br_snapshots_11_10; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_132 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_11 : br_snapshots_0_11; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_133 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_11 : br_snapshots_1_11; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_134 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_11 : br_snapshots_2_11; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_135 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_11 : br_snapshots_3_11; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_136 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_11 : br_snapshots_4_11; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_137 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_11 : br_snapshots_5_11; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_138 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_11 : br_snapshots_6_11; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_139 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_11 : br_snapshots_7_11; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_140 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_11 : br_snapshots_8_11; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_141 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_11 : br_snapshots_9_11; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_142 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_11 : br_snapshots_10_11; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_143 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_11 : br_snapshots_11_11; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_144 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_12 : br_snapshots_0_12; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_145 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_12 : br_snapshots_1_12; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_146 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_12 : br_snapshots_2_12; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_147 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_12 : br_snapshots_3_12; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_148 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_12 : br_snapshots_4_12; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_149 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_12 : br_snapshots_5_12; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_150 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_12 : br_snapshots_6_12; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_151 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_12 : br_snapshots_7_12; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_152 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_12 : br_snapshots_8_12; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_153 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_12 : br_snapshots_9_12; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_154 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_12 : br_snapshots_10_12; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_155 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_12 : br_snapshots_11_12; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_156 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_13 : br_snapshots_0_13; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_157 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_13 : br_snapshots_1_13; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_158 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_13 : br_snapshots_2_13; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_159 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_13 : br_snapshots_3_13; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_160 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_13 : br_snapshots_4_13; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_161 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_13 : br_snapshots_5_13; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_162 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_13 : br_snapshots_6_13; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_163 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_13 : br_snapshots_7_13; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_164 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_13 : br_snapshots_8_13; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_165 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_13 : br_snapshots_9_13; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_166 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_13 : br_snapshots_10_13; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_167 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_13 : br_snapshots_11_13; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_168 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_14 : br_snapshots_0_14; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_169 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_14 : br_snapshots_1_14; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_170 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_14 : br_snapshots_2_14; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_171 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_14 : br_snapshots_3_14; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_172 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_14 : br_snapshots_4_14; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_173 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_14 : br_snapshots_5_14; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_174 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_14 : br_snapshots_6_14; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_175 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_14 : br_snapshots_7_14; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_176 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_14 : br_snapshots_8_14; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_177 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_14 : br_snapshots_9_14; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_178 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_14 : br_snapshots_10_14; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_179 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_14 : br_snapshots_11_14; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_180 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_15 : br_snapshots_0_15; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_181 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_15 : br_snapshots_1_15; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_182 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_15 : br_snapshots_2_15; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_183 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_15 : br_snapshots_3_15; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_184 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_15 : br_snapshots_4_15; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_185 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_15 : br_snapshots_5_15; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_186 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_15 : br_snapshots_6_15; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_187 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_15 : br_snapshots_7_15; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_188 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_15 : br_snapshots_8_15; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_189 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_15 : br_snapshots_9_15; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_190 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_15 : br_snapshots_10_15; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_191 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_15 : br_snapshots_11_15; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_192 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_16 : br_snapshots_0_16; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_193 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_16 : br_snapshots_1_16; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_194 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_16 : br_snapshots_2_16; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_195 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_16 : br_snapshots_3_16; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_196 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_16 : br_snapshots_4_16; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_197 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_16 : br_snapshots_5_16; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_198 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_16 : br_snapshots_6_16; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_199 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_16 : br_snapshots_7_16; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_200 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_16 : br_snapshots_8_16; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_201 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_16 : br_snapshots_9_16; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_202 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_16 : br_snapshots_10_16; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_203 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_16 : br_snapshots_11_16; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_204 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_17 : br_snapshots_0_17; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_205 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_17 : br_snapshots_1_17; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_206 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_17 : br_snapshots_2_17; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_207 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_17 : br_snapshots_3_17; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_208 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_17 : br_snapshots_4_17; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_209 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_17 : br_snapshots_5_17; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_210 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_17 : br_snapshots_6_17; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_211 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_17 : br_snapshots_7_17; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_212 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_17 : br_snapshots_8_17; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_213 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_17 : br_snapshots_9_17; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_214 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_17 : br_snapshots_10_17; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_215 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_17 : br_snapshots_11_17; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_216 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_18 : br_snapshots_0_18; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_217 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_18 : br_snapshots_1_18; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_218 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_18 : br_snapshots_2_18; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_219 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_18 : br_snapshots_3_18; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_220 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_18 : br_snapshots_4_18; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_221 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_18 : br_snapshots_5_18; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_222 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_18 : br_snapshots_6_18; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_223 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_18 : br_snapshots_7_18; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_224 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_18 : br_snapshots_8_18; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_225 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_18 : br_snapshots_9_18; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_226 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_18 : br_snapshots_10_18; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_227 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_18 : br_snapshots_11_18; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_228 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_19 : br_snapshots_0_19; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_229 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_19 : br_snapshots_1_19; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_230 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_19 : br_snapshots_2_19; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_231 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_19 : br_snapshots_3_19; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_232 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_19 : br_snapshots_4_19; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_233 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_19 : br_snapshots_5_19; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_234 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_19 : br_snapshots_6_19; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_235 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_19 : br_snapshots_7_19; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_236 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_19 : br_snapshots_8_19; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_237 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_19 : br_snapshots_9_19; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_238 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_19 : br_snapshots_10_19; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_239 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_19 : br_snapshots_11_19; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_240 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_20 : br_snapshots_0_20; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_241 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_20 : br_snapshots_1_20; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_242 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_20 : br_snapshots_2_20; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_243 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_20 : br_snapshots_3_20; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_244 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_20 : br_snapshots_4_20; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_245 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_20 : br_snapshots_5_20; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_246 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_20 : br_snapshots_6_20; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_247 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_20 : br_snapshots_7_20; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_248 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_20 : br_snapshots_8_20; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_249 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_20 : br_snapshots_9_20; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_250 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_20 : br_snapshots_10_20; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_251 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_20 : br_snapshots_11_20; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_252 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_21 : br_snapshots_0_21; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_253 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_21 : br_snapshots_1_21; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_254 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_21 : br_snapshots_2_21; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_255 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_21 : br_snapshots_3_21; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_256 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_21 : br_snapshots_4_21; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_257 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_21 : br_snapshots_5_21; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_258 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_21 : br_snapshots_6_21; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_259 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_21 : br_snapshots_7_21; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_260 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_21 : br_snapshots_8_21; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_261 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_21 : br_snapshots_9_21; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_262 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_21 : br_snapshots_10_21; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_263 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_21 : br_snapshots_11_21; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_264 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_22 : br_snapshots_0_22; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_265 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_22 : br_snapshots_1_22; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_266 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_22 : br_snapshots_2_22; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_267 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_22 : br_snapshots_3_22; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_268 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_22 : br_snapshots_4_22; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_269 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_22 : br_snapshots_5_22; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_270 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_22 : br_snapshots_6_22; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_271 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_22 : br_snapshots_7_22; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_272 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_22 : br_snapshots_8_22; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_273 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_22 : br_snapshots_9_22; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_274 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_22 : br_snapshots_10_22; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_275 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_22 : br_snapshots_11_22; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_276 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_23 : br_snapshots_0_23; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_277 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_23 : br_snapshots_1_23; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_278 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_23 : br_snapshots_2_23; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_279 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_23 : br_snapshots_3_23; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_280 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_23 : br_snapshots_4_23; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_281 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_23 : br_snapshots_5_23; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_282 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_23 : br_snapshots_6_23; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_283 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_23 : br_snapshots_7_23; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_284 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_23 : br_snapshots_8_23; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_285 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_23 : br_snapshots_9_23; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_286 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_23 : br_snapshots_10_23; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_287 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_23 : br_snapshots_11_23; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_288 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_24 : br_snapshots_0_24; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_289 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_24 : br_snapshots_1_24; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_290 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_24 : br_snapshots_2_24; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_291 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_24 : br_snapshots_3_24; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_292 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_24 : br_snapshots_4_24; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_293 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_24 : br_snapshots_5_24; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_294 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_24 : br_snapshots_6_24; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_295 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_24 : br_snapshots_7_24; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_296 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_24 : br_snapshots_8_24; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_297 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_24 : br_snapshots_9_24; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_298 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_24 : br_snapshots_10_24; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_299 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_24 : br_snapshots_11_24; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_300 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_25 : br_snapshots_0_25; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_301 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_25 : br_snapshots_1_25; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_302 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_25 : br_snapshots_2_25; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_303 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_25 : br_snapshots_3_25; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_304 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_25 : br_snapshots_4_25; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_305 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_25 : br_snapshots_5_25; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_306 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_25 : br_snapshots_6_25; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_307 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_25 : br_snapshots_7_25; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_308 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_25 : br_snapshots_8_25; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_309 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_25 : br_snapshots_9_25; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_310 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_25 : br_snapshots_10_25; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_311 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_25 : br_snapshots_11_25; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_312 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_26 : br_snapshots_0_26; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_313 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_26 : br_snapshots_1_26; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_314 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_26 : br_snapshots_2_26; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_315 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_26 : br_snapshots_3_26; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_316 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_26 : br_snapshots_4_26; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_317 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_26 : br_snapshots_5_26; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_318 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_26 : br_snapshots_6_26; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_319 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_26 : br_snapshots_7_26; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_320 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_26 : br_snapshots_8_26; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_321 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_26 : br_snapshots_9_26; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_322 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_26 : br_snapshots_10_26; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_323 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_26 : br_snapshots_11_26; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_324 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_27 : br_snapshots_0_27; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_325 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_27 : br_snapshots_1_27; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_326 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_27 : br_snapshots_2_27; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_327 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_27 : br_snapshots_3_27; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_328 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_27 : br_snapshots_4_27; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_329 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_27 : br_snapshots_5_27; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_330 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_27 : br_snapshots_6_27; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_331 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_27 : br_snapshots_7_27; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_332 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_27 : br_snapshots_8_27; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_333 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_27 : br_snapshots_9_27; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_334 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_27 : br_snapshots_10_27; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_335 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_27 : br_snapshots_11_27; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_336 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_28 : br_snapshots_0_28; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_337 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_28 : br_snapshots_1_28; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_338 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_28 : br_snapshots_2_28; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_339 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_28 : br_snapshots_3_28; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_340 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_28 : br_snapshots_4_28; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_341 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_28 : br_snapshots_5_28; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_342 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_28 : br_snapshots_6_28; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_343 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_28 : br_snapshots_7_28; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_344 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_28 : br_snapshots_8_28; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_345 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_28 : br_snapshots_9_28; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_346 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_28 : br_snapshots_10_28; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_347 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_28 : br_snapshots_11_28; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_348 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_29 : br_snapshots_0_29; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_349 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_29 : br_snapshots_1_29; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_350 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_29 : br_snapshots_2_29; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_351 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_29 : br_snapshots_3_29; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_352 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_29 : br_snapshots_4_29; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_353 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_29 : br_snapshots_5_29; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_354 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_29 : br_snapshots_6_29; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_355 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_29 : br_snapshots_7_29; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_356 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_29 : br_snapshots_8_29; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_357 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_29 : br_snapshots_9_29; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_358 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_29 : br_snapshots_10_29; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_359 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_29 : br_snapshots_11_29; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_360 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_30 : br_snapshots_0_30; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_361 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_30 : br_snapshots_1_30; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_362 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_30 : br_snapshots_2_30; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_363 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_30 : br_snapshots_3_30; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_364 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_30 : br_snapshots_4_30; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_365 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_30 : br_snapshots_5_30; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_366 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_30 : br_snapshots_6_30; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_367 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_30 : br_snapshots_7_30; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_368 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_30 : br_snapshots_8_30; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_369 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_30 : br_snapshots_9_30; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_370 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_30 : br_snapshots_10_30; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_371 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_30 : br_snapshots_11_30; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_372 = 4'h0 == io_ren_br_tags_0_bits ? remap_table_1_31 : br_snapshots_0_31; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_373 = 4'h1 == io_ren_br_tags_0_bits ? remap_table_1_31 : br_snapshots_1_31; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_374 = 4'h2 == io_ren_br_tags_0_bits ? remap_table_1_31 : br_snapshots_2_31; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_375 = 4'h3 == io_ren_br_tags_0_bits ? remap_table_1_31 : br_snapshots_3_31; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_376 = 4'h4 == io_ren_br_tags_0_bits ? remap_table_1_31 : br_snapshots_4_31; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_377 = 4'h5 == io_ren_br_tags_0_bits ? remap_table_1_31 : br_snapshots_5_31; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_378 = 4'h6 == io_ren_br_tags_0_bits ? remap_table_1_31 : br_snapshots_6_31; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_379 = 4'h7 == io_ren_br_tags_0_bits ? remap_table_1_31 : br_snapshots_7_31; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_380 = 4'h8 == io_ren_br_tags_0_bits ? remap_table_1_31 : br_snapshots_8_31; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_381 = 4'h9 == io_ren_br_tags_0_bits ? remap_table_1_31 : br_snapshots_9_31; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_382 = 4'ha == io_ren_br_tags_0_bits ? remap_table_1_31 : br_snapshots_10_31; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_383 = 4'hb == io_ren_br_tags_0_bits ? remap_table_1_31 : br_snapshots_11_31; // @[rename-maptable.scala 133:44 rename-maptable.scala 133:44 rename-maptable.scala 79:25]
  wire [5:0] _GEN_396 = io_ren_br_tags_0_valid ? _GEN_12 : br_snapshots_0_1; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_397 = io_ren_br_tags_0_valid ? _GEN_13 : br_snapshots_1_1; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_398 = io_ren_br_tags_0_valid ? _GEN_14 : br_snapshots_2_1; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_399 = io_ren_br_tags_0_valid ? _GEN_15 : br_snapshots_3_1; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_400 = io_ren_br_tags_0_valid ? _GEN_16 : br_snapshots_4_1; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_401 = io_ren_br_tags_0_valid ? _GEN_17 : br_snapshots_5_1; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_402 = io_ren_br_tags_0_valid ? _GEN_18 : br_snapshots_6_1; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_403 = io_ren_br_tags_0_valid ? _GEN_19 : br_snapshots_7_1; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_404 = io_ren_br_tags_0_valid ? _GEN_20 : br_snapshots_8_1; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_405 = io_ren_br_tags_0_valid ? _GEN_21 : br_snapshots_9_1; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_406 = io_ren_br_tags_0_valid ? _GEN_22 : br_snapshots_10_1; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_407 = io_ren_br_tags_0_valid ? _GEN_23 : br_snapshots_11_1; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_408 = io_ren_br_tags_0_valid ? _GEN_24 : br_snapshots_0_2; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_409 = io_ren_br_tags_0_valid ? _GEN_25 : br_snapshots_1_2; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_410 = io_ren_br_tags_0_valid ? _GEN_26 : br_snapshots_2_2; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_411 = io_ren_br_tags_0_valid ? _GEN_27 : br_snapshots_3_2; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_412 = io_ren_br_tags_0_valid ? _GEN_28 : br_snapshots_4_2; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_413 = io_ren_br_tags_0_valid ? _GEN_29 : br_snapshots_5_2; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_414 = io_ren_br_tags_0_valid ? _GEN_30 : br_snapshots_6_2; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_415 = io_ren_br_tags_0_valid ? _GEN_31 : br_snapshots_7_2; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_416 = io_ren_br_tags_0_valid ? _GEN_32 : br_snapshots_8_2; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_417 = io_ren_br_tags_0_valid ? _GEN_33 : br_snapshots_9_2; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_418 = io_ren_br_tags_0_valid ? _GEN_34 : br_snapshots_10_2; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_419 = io_ren_br_tags_0_valid ? _GEN_35 : br_snapshots_11_2; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_420 = io_ren_br_tags_0_valid ? _GEN_36 : br_snapshots_0_3; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_421 = io_ren_br_tags_0_valid ? _GEN_37 : br_snapshots_1_3; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_422 = io_ren_br_tags_0_valid ? _GEN_38 : br_snapshots_2_3; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_423 = io_ren_br_tags_0_valid ? _GEN_39 : br_snapshots_3_3; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_424 = io_ren_br_tags_0_valid ? _GEN_40 : br_snapshots_4_3; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_425 = io_ren_br_tags_0_valid ? _GEN_41 : br_snapshots_5_3; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_426 = io_ren_br_tags_0_valid ? _GEN_42 : br_snapshots_6_3; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_427 = io_ren_br_tags_0_valid ? _GEN_43 : br_snapshots_7_3; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_428 = io_ren_br_tags_0_valid ? _GEN_44 : br_snapshots_8_3; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_429 = io_ren_br_tags_0_valid ? _GEN_45 : br_snapshots_9_3; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_430 = io_ren_br_tags_0_valid ? _GEN_46 : br_snapshots_10_3; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_431 = io_ren_br_tags_0_valid ? _GEN_47 : br_snapshots_11_3; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_432 = io_ren_br_tags_0_valid ? _GEN_48 : br_snapshots_0_4; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_433 = io_ren_br_tags_0_valid ? _GEN_49 : br_snapshots_1_4; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_434 = io_ren_br_tags_0_valid ? _GEN_50 : br_snapshots_2_4; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_435 = io_ren_br_tags_0_valid ? _GEN_51 : br_snapshots_3_4; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_436 = io_ren_br_tags_0_valid ? _GEN_52 : br_snapshots_4_4; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_437 = io_ren_br_tags_0_valid ? _GEN_53 : br_snapshots_5_4; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_438 = io_ren_br_tags_0_valid ? _GEN_54 : br_snapshots_6_4; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_439 = io_ren_br_tags_0_valid ? _GEN_55 : br_snapshots_7_4; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_440 = io_ren_br_tags_0_valid ? _GEN_56 : br_snapshots_8_4; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_441 = io_ren_br_tags_0_valid ? _GEN_57 : br_snapshots_9_4; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_442 = io_ren_br_tags_0_valid ? _GEN_58 : br_snapshots_10_4; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_443 = io_ren_br_tags_0_valid ? _GEN_59 : br_snapshots_11_4; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_444 = io_ren_br_tags_0_valid ? _GEN_60 : br_snapshots_0_5; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_445 = io_ren_br_tags_0_valid ? _GEN_61 : br_snapshots_1_5; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_446 = io_ren_br_tags_0_valid ? _GEN_62 : br_snapshots_2_5; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_447 = io_ren_br_tags_0_valid ? _GEN_63 : br_snapshots_3_5; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_448 = io_ren_br_tags_0_valid ? _GEN_64 : br_snapshots_4_5; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_449 = io_ren_br_tags_0_valid ? _GEN_65 : br_snapshots_5_5; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_450 = io_ren_br_tags_0_valid ? _GEN_66 : br_snapshots_6_5; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_451 = io_ren_br_tags_0_valid ? _GEN_67 : br_snapshots_7_5; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_452 = io_ren_br_tags_0_valid ? _GEN_68 : br_snapshots_8_5; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_453 = io_ren_br_tags_0_valid ? _GEN_69 : br_snapshots_9_5; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_454 = io_ren_br_tags_0_valid ? _GEN_70 : br_snapshots_10_5; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_455 = io_ren_br_tags_0_valid ? _GEN_71 : br_snapshots_11_5; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_456 = io_ren_br_tags_0_valid ? _GEN_72 : br_snapshots_0_6; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_457 = io_ren_br_tags_0_valid ? _GEN_73 : br_snapshots_1_6; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_458 = io_ren_br_tags_0_valid ? _GEN_74 : br_snapshots_2_6; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_459 = io_ren_br_tags_0_valid ? _GEN_75 : br_snapshots_3_6; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_460 = io_ren_br_tags_0_valid ? _GEN_76 : br_snapshots_4_6; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_461 = io_ren_br_tags_0_valid ? _GEN_77 : br_snapshots_5_6; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_462 = io_ren_br_tags_0_valid ? _GEN_78 : br_snapshots_6_6; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_463 = io_ren_br_tags_0_valid ? _GEN_79 : br_snapshots_7_6; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_464 = io_ren_br_tags_0_valid ? _GEN_80 : br_snapshots_8_6; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_465 = io_ren_br_tags_0_valid ? _GEN_81 : br_snapshots_9_6; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_466 = io_ren_br_tags_0_valid ? _GEN_82 : br_snapshots_10_6; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_467 = io_ren_br_tags_0_valid ? _GEN_83 : br_snapshots_11_6; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_468 = io_ren_br_tags_0_valid ? _GEN_84 : br_snapshots_0_7; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_469 = io_ren_br_tags_0_valid ? _GEN_85 : br_snapshots_1_7; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_470 = io_ren_br_tags_0_valid ? _GEN_86 : br_snapshots_2_7; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_471 = io_ren_br_tags_0_valid ? _GEN_87 : br_snapshots_3_7; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_472 = io_ren_br_tags_0_valid ? _GEN_88 : br_snapshots_4_7; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_473 = io_ren_br_tags_0_valid ? _GEN_89 : br_snapshots_5_7; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_474 = io_ren_br_tags_0_valid ? _GEN_90 : br_snapshots_6_7; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_475 = io_ren_br_tags_0_valid ? _GEN_91 : br_snapshots_7_7; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_476 = io_ren_br_tags_0_valid ? _GEN_92 : br_snapshots_8_7; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_477 = io_ren_br_tags_0_valid ? _GEN_93 : br_snapshots_9_7; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_478 = io_ren_br_tags_0_valid ? _GEN_94 : br_snapshots_10_7; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_479 = io_ren_br_tags_0_valid ? _GEN_95 : br_snapshots_11_7; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_480 = io_ren_br_tags_0_valid ? _GEN_96 : br_snapshots_0_8; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_481 = io_ren_br_tags_0_valid ? _GEN_97 : br_snapshots_1_8; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_482 = io_ren_br_tags_0_valid ? _GEN_98 : br_snapshots_2_8; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_483 = io_ren_br_tags_0_valid ? _GEN_99 : br_snapshots_3_8; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_484 = io_ren_br_tags_0_valid ? _GEN_100 : br_snapshots_4_8; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_485 = io_ren_br_tags_0_valid ? _GEN_101 : br_snapshots_5_8; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_486 = io_ren_br_tags_0_valid ? _GEN_102 : br_snapshots_6_8; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_487 = io_ren_br_tags_0_valid ? _GEN_103 : br_snapshots_7_8; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_488 = io_ren_br_tags_0_valid ? _GEN_104 : br_snapshots_8_8; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_489 = io_ren_br_tags_0_valid ? _GEN_105 : br_snapshots_9_8; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_490 = io_ren_br_tags_0_valid ? _GEN_106 : br_snapshots_10_8; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_491 = io_ren_br_tags_0_valid ? _GEN_107 : br_snapshots_11_8; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_492 = io_ren_br_tags_0_valid ? _GEN_108 : br_snapshots_0_9; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_493 = io_ren_br_tags_0_valid ? _GEN_109 : br_snapshots_1_9; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_494 = io_ren_br_tags_0_valid ? _GEN_110 : br_snapshots_2_9; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_495 = io_ren_br_tags_0_valid ? _GEN_111 : br_snapshots_3_9; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_496 = io_ren_br_tags_0_valid ? _GEN_112 : br_snapshots_4_9; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_497 = io_ren_br_tags_0_valid ? _GEN_113 : br_snapshots_5_9; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_498 = io_ren_br_tags_0_valid ? _GEN_114 : br_snapshots_6_9; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_499 = io_ren_br_tags_0_valid ? _GEN_115 : br_snapshots_7_9; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_500 = io_ren_br_tags_0_valid ? _GEN_116 : br_snapshots_8_9; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_501 = io_ren_br_tags_0_valid ? _GEN_117 : br_snapshots_9_9; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_502 = io_ren_br_tags_0_valid ? _GEN_118 : br_snapshots_10_9; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_503 = io_ren_br_tags_0_valid ? _GEN_119 : br_snapshots_11_9; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_504 = io_ren_br_tags_0_valid ? _GEN_120 : br_snapshots_0_10; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_505 = io_ren_br_tags_0_valid ? _GEN_121 : br_snapshots_1_10; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_506 = io_ren_br_tags_0_valid ? _GEN_122 : br_snapshots_2_10; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_507 = io_ren_br_tags_0_valid ? _GEN_123 : br_snapshots_3_10; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_508 = io_ren_br_tags_0_valid ? _GEN_124 : br_snapshots_4_10; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_509 = io_ren_br_tags_0_valid ? _GEN_125 : br_snapshots_5_10; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_510 = io_ren_br_tags_0_valid ? _GEN_126 : br_snapshots_6_10; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_511 = io_ren_br_tags_0_valid ? _GEN_127 : br_snapshots_7_10; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_512 = io_ren_br_tags_0_valid ? _GEN_128 : br_snapshots_8_10; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_513 = io_ren_br_tags_0_valid ? _GEN_129 : br_snapshots_9_10; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_514 = io_ren_br_tags_0_valid ? _GEN_130 : br_snapshots_10_10; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_515 = io_ren_br_tags_0_valid ? _GEN_131 : br_snapshots_11_10; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_516 = io_ren_br_tags_0_valid ? _GEN_132 : br_snapshots_0_11; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_517 = io_ren_br_tags_0_valid ? _GEN_133 : br_snapshots_1_11; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_518 = io_ren_br_tags_0_valid ? _GEN_134 : br_snapshots_2_11; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_519 = io_ren_br_tags_0_valid ? _GEN_135 : br_snapshots_3_11; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_520 = io_ren_br_tags_0_valid ? _GEN_136 : br_snapshots_4_11; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_521 = io_ren_br_tags_0_valid ? _GEN_137 : br_snapshots_5_11; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_522 = io_ren_br_tags_0_valid ? _GEN_138 : br_snapshots_6_11; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_523 = io_ren_br_tags_0_valid ? _GEN_139 : br_snapshots_7_11; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_524 = io_ren_br_tags_0_valid ? _GEN_140 : br_snapshots_8_11; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_525 = io_ren_br_tags_0_valid ? _GEN_141 : br_snapshots_9_11; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_526 = io_ren_br_tags_0_valid ? _GEN_142 : br_snapshots_10_11; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_527 = io_ren_br_tags_0_valid ? _GEN_143 : br_snapshots_11_11; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_528 = io_ren_br_tags_0_valid ? _GEN_144 : br_snapshots_0_12; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_529 = io_ren_br_tags_0_valid ? _GEN_145 : br_snapshots_1_12; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_530 = io_ren_br_tags_0_valid ? _GEN_146 : br_snapshots_2_12; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_531 = io_ren_br_tags_0_valid ? _GEN_147 : br_snapshots_3_12; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_532 = io_ren_br_tags_0_valid ? _GEN_148 : br_snapshots_4_12; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_533 = io_ren_br_tags_0_valid ? _GEN_149 : br_snapshots_5_12; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_534 = io_ren_br_tags_0_valid ? _GEN_150 : br_snapshots_6_12; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_535 = io_ren_br_tags_0_valid ? _GEN_151 : br_snapshots_7_12; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_536 = io_ren_br_tags_0_valid ? _GEN_152 : br_snapshots_8_12; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_537 = io_ren_br_tags_0_valid ? _GEN_153 : br_snapshots_9_12; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_538 = io_ren_br_tags_0_valid ? _GEN_154 : br_snapshots_10_12; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_539 = io_ren_br_tags_0_valid ? _GEN_155 : br_snapshots_11_12; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_540 = io_ren_br_tags_0_valid ? _GEN_156 : br_snapshots_0_13; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_541 = io_ren_br_tags_0_valid ? _GEN_157 : br_snapshots_1_13; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_542 = io_ren_br_tags_0_valid ? _GEN_158 : br_snapshots_2_13; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_543 = io_ren_br_tags_0_valid ? _GEN_159 : br_snapshots_3_13; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_544 = io_ren_br_tags_0_valid ? _GEN_160 : br_snapshots_4_13; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_545 = io_ren_br_tags_0_valid ? _GEN_161 : br_snapshots_5_13; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_546 = io_ren_br_tags_0_valid ? _GEN_162 : br_snapshots_6_13; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_547 = io_ren_br_tags_0_valid ? _GEN_163 : br_snapshots_7_13; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_548 = io_ren_br_tags_0_valid ? _GEN_164 : br_snapshots_8_13; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_549 = io_ren_br_tags_0_valid ? _GEN_165 : br_snapshots_9_13; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_550 = io_ren_br_tags_0_valid ? _GEN_166 : br_snapshots_10_13; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_551 = io_ren_br_tags_0_valid ? _GEN_167 : br_snapshots_11_13; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_552 = io_ren_br_tags_0_valid ? _GEN_168 : br_snapshots_0_14; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_553 = io_ren_br_tags_0_valid ? _GEN_169 : br_snapshots_1_14; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_554 = io_ren_br_tags_0_valid ? _GEN_170 : br_snapshots_2_14; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_555 = io_ren_br_tags_0_valid ? _GEN_171 : br_snapshots_3_14; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_556 = io_ren_br_tags_0_valid ? _GEN_172 : br_snapshots_4_14; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_557 = io_ren_br_tags_0_valid ? _GEN_173 : br_snapshots_5_14; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_558 = io_ren_br_tags_0_valid ? _GEN_174 : br_snapshots_6_14; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_559 = io_ren_br_tags_0_valid ? _GEN_175 : br_snapshots_7_14; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_560 = io_ren_br_tags_0_valid ? _GEN_176 : br_snapshots_8_14; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_561 = io_ren_br_tags_0_valid ? _GEN_177 : br_snapshots_9_14; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_562 = io_ren_br_tags_0_valid ? _GEN_178 : br_snapshots_10_14; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_563 = io_ren_br_tags_0_valid ? _GEN_179 : br_snapshots_11_14; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_564 = io_ren_br_tags_0_valid ? _GEN_180 : br_snapshots_0_15; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_565 = io_ren_br_tags_0_valid ? _GEN_181 : br_snapshots_1_15; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_566 = io_ren_br_tags_0_valid ? _GEN_182 : br_snapshots_2_15; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_567 = io_ren_br_tags_0_valid ? _GEN_183 : br_snapshots_3_15; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_568 = io_ren_br_tags_0_valid ? _GEN_184 : br_snapshots_4_15; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_569 = io_ren_br_tags_0_valid ? _GEN_185 : br_snapshots_5_15; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_570 = io_ren_br_tags_0_valid ? _GEN_186 : br_snapshots_6_15; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_571 = io_ren_br_tags_0_valid ? _GEN_187 : br_snapshots_7_15; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_572 = io_ren_br_tags_0_valid ? _GEN_188 : br_snapshots_8_15; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_573 = io_ren_br_tags_0_valid ? _GEN_189 : br_snapshots_9_15; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_574 = io_ren_br_tags_0_valid ? _GEN_190 : br_snapshots_10_15; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_575 = io_ren_br_tags_0_valid ? _GEN_191 : br_snapshots_11_15; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_576 = io_ren_br_tags_0_valid ? _GEN_192 : br_snapshots_0_16; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_577 = io_ren_br_tags_0_valid ? _GEN_193 : br_snapshots_1_16; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_578 = io_ren_br_tags_0_valid ? _GEN_194 : br_snapshots_2_16; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_579 = io_ren_br_tags_0_valid ? _GEN_195 : br_snapshots_3_16; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_580 = io_ren_br_tags_0_valid ? _GEN_196 : br_snapshots_4_16; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_581 = io_ren_br_tags_0_valid ? _GEN_197 : br_snapshots_5_16; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_582 = io_ren_br_tags_0_valid ? _GEN_198 : br_snapshots_6_16; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_583 = io_ren_br_tags_0_valid ? _GEN_199 : br_snapshots_7_16; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_584 = io_ren_br_tags_0_valid ? _GEN_200 : br_snapshots_8_16; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_585 = io_ren_br_tags_0_valid ? _GEN_201 : br_snapshots_9_16; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_586 = io_ren_br_tags_0_valid ? _GEN_202 : br_snapshots_10_16; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_587 = io_ren_br_tags_0_valid ? _GEN_203 : br_snapshots_11_16; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_588 = io_ren_br_tags_0_valid ? _GEN_204 : br_snapshots_0_17; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_589 = io_ren_br_tags_0_valid ? _GEN_205 : br_snapshots_1_17; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_590 = io_ren_br_tags_0_valid ? _GEN_206 : br_snapshots_2_17; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_591 = io_ren_br_tags_0_valid ? _GEN_207 : br_snapshots_3_17; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_592 = io_ren_br_tags_0_valid ? _GEN_208 : br_snapshots_4_17; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_593 = io_ren_br_tags_0_valid ? _GEN_209 : br_snapshots_5_17; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_594 = io_ren_br_tags_0_valid ? _GEN_210 : br_snapshots_6_17; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_595 = io_ren_br_tags_0_valid ? _GEN_211 : br_snapshots_7_17; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_596 = io_ren_br_tags_0_valid ? _GEN_212 : br_snapshots_8_17; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_597 = io_ren_br_tags_0_valid ? _GEN_213 : br_snapshots_9_17; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_598 = io_ren_br_tags_0_valid ? _GEN_214 : br_snapshots_10_17; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_599 = io_ren_br_tags_0_valid ? _GEN_215 : br_snapshots_11_17; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_600 = io_ren_br_tags_0_valid ? _GEN_216 : br_snapshots_0_18; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_601 = io_ren_br_tags_0_valid ? _GEN_217 : br_snapshots_1_18; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_602 = io_ren_br_tags_0_valid ? _GEN_218 : br_snapshots_2_18; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_603 = io_ren_br_tags_0_valid ? _GEN_219 : br_snapshots_3_18; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_604 = io_ren_br_tags_0_valid ? _GEN_220 : br_snapshots_4_18; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_605 = io_ren_br_tags_0_valid ? _GEN_221 : br_snapshots_5_18; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_606 = io_ren_br_tags_0_valid ? _GEN_222 : br_snapshots_6_18; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_607 = io_ren_br_tags_0_valid ? _GEN_223 : br_snapshots_7_18; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_608 = io_ren_br_tags_0_valid ? _GEN_224 : br_snapshots_8_18; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_609 = io_ren_br_tags_0_valid ? _GEN_225 : br_snapshots_9_18; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_610 = io_ren_br_tags_0_valid ? _GEN_226 : br_snapshots_10_18; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_611 = io_ren_br_tags_0_valid ? _GEN_227 : br_snapshots_11_18; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_612 = io_ren_br_tags_0_valid ? _GEN_228 : br_snapshots_0_19; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_613 = io_ren_br_tags_0_valid ? _GEN_229 : br_snapshots_1_19; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_614 = io_ren_br_tags_0_valid ? _GEN_230 : br_snapshots_2_19; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_615 = io_ren_br_tags_0_valid ? _GEN_231 : br_snapshots_3_19; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_616 = io_ren_br_tags_0_valid ? _GEN_232 : br_snapshots_4_19; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_617 = io_ren_br_tags_0_valid ? _GEN_233 : br_snapshots_5_19; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_618 = io_ren_br_tags_0_valid ? _GEN_234 : br_snapshots_6_19; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_619 = io_ren_br_tags_0_valid ? _GEN_235 : br_snapshots_7_19; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_620 = io_ren_br_tags_0_valid ? _GEN_236 : br_snapshots_8_19; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_621 = io_ren_br_tags_0_valid ? _GEN_237 : br_snapshots_9_19; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_622 = io_ren_br_tags_0_valid ? _GEN_238 : br_snapshots_10_19; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_623 = io_ren_br_tags_0_valid ? _GEN_239 : br_snapshots_11_19; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_624 = io_ren_br_tags_0_valid ? _GEN_240 : br_snapshots_0_20; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_625 = io_ren_br_tags_0_valid ? _GEN_241 : br_snapshots_1_20; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_626 = io_ren_br_tags_0_valid ? _GEN_242 : br_snapshots_2_20; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_627 = io_ren_br_tags_0_valid ? _GEN_243 : br_snapshots_3_20; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_628 = io_ren_br_tags_0_valid ? _GEN_244 : br_snapshots_4_20; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_629 = io_ren_br_tags_0_valid ? _GEN_245 : br_snapshots_5_20; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_630 = io_ren_br_tags_0_valid ? _GEN_246 : br_snapshots_6_20; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_631 = io_ren_br_tags_0_valid ? _GEN_247 : br_snapshots_7_20; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_632 = io_ren_br_tags_0_valid ? _GEN_248 : br_snapshots_8_20; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_633 = io_ren_br_tags_0_valid ? _GEN_249 : br_snapshots_9_20; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_634 = io_ren_br_tags_0_valid ? _GEN_250 : br_snapshots_10_20; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_635 = io_ren_br_tags_0_valid ? _GEN_251 : br_snapshots_11_20; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_636 = io_ren_br_tags_0_valid ? _GEN_252 : br_snapshots_0_21; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_637 = io_ren_br_tags_0_valid ? _GEN_253 : br_snapshots_1_21; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_638 = io_ren_br_tags_0_valid ? _GEN_254 : br_snapshots_2_21; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_639 = io_ren_br_tags_0_valid ? _GEN_255 : br_snapshots_3_21; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_640 = io_ren_br_tags_0_valid ? _GEN_256 : br_snapshots_4_21; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_641 = io_ren_br_tags_0_valid ? _GEN_257 : br_snapshots_5_21; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_642 = io_ren_br_tags_0_valid ? _GEN_258 : br_snapshots_6_21; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_643 = io_ren_br_tags_0_valid ? _GEN_259 : br_snapshots_7_21; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_644 = io_ren_br_tags_0_valid ? _GEN_260 : br_snapshots_8_21; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_645 = io_ren_br_tags_0_valid ? _GEN_261 : br_snapshots_9_21; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_646 = io_ren_br_tags_0_valid ? _GEN_262 : br_snapshots_10_21; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_647 = io_ren_br_tags_0_valid ? _GEN_263 : br_snapshots_11_21; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_648 = io_ren_br_tags_0_valid ? _GEN_264 : br_snapshots_0_22; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_649 = io_ren_br_tags_0_valid ? _GEN_265 : br_snapshots_1_22; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_650 = io_ren_br_tags_0_valid ? _GEN_266 : br_snapshots_2_22; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_651 = io_ren_br_tags_0_valid ? _GEN_267 : br_snapshots_3_22; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_652 = io_ren_br_tags_0_valid ? _GEN_268 : br_snapshots_4_22; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_653 = io_ren_br_tags_0_valid ? _GEN_269 : br_snapshots_5_22; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_654 = io_ren_br_tags_0_valid ? _GEN_270 : br_snapshots_6_22; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_655 = io_ren_br_tags_0_valid ? _GEN_271 : br_snapshots_7_22; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_656 = io_ren_br_tags_0_valid ? _GEN_272 : br_snapshots_8_22; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_657 = io_ren_br_tags_0_valid ? _GEN_273 : br_snapshots_9_22; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_658 = io_ren_br_tags_0_valid ? _GEN_274 : br_snapshots_10_22; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_659 = io_ren_br_tags_0_valid ? _GEN_275 : br_snapshots_11_22; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_660 = io_ren_br_tags_0_valid ? _GEN_276 : br_snapshots_0_23; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_661 = io_ren_br_tags_0_valid ? _GEN_277 : br_snapshots_1_23; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_662 = io_ren_br_tags_0_valid ? _GEN_278 : br_snapshots_2_23; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_663 = io_ren_br_tags_0_valid ? _GEN_279 : br_snapshots_3_23; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_664 = io_ren_br_tags_0_valid ? _GEN_280 : br_snapshots_4_23; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_665 = io_ren_br_tags_0_valid ? _GEN_281 : br_snapshots_5_23; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_666 = io_ren_br_tags_0_valid ? _GEN_282 : br_snapshots_6_23; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_667 = io_ren_br_tags_0_valid ? _GEN_283 : br_snapshots_7_23; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_668 = io_ren_br_tags_0_valid ? _GEN_284 : br_snapshots_8_23; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_669 = io_ren_br_tags_0_valid ? _GEN_285 : br_snapshots_9_23; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_670 = io_ren_br_tags_0_valid ? _GEN_286 : br_snapshots_10_23; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_671 = io_ren_br_tags_0_valid ? _GEN_287 : br_snapshots_11_23; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_672 = io_ren_br_tags_0_valid ? _GEN_288 : br_snapshots_0_24; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_673 = io_ren_br_tags_0_valid ? _GEN_289 : br_snapshots_1_24; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_674 = io_ren_br_tags_0_valid ? _GEN_290 : br_snapshots_2_24; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_675 = io_ren_br_tags_0_valid ? _GEN_291 : br_snapshots_3_24; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_676 = io_ren_br_tags_0_valid ? _GEN_292 : br_snapshots_4_24; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_677 = io_ren_br_tags_0_valid ? _GEN_293 : br_snapshots_5_24; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_678 = io_ren_br_tags_0_valid ? _GEN_294 : br_snapshots_6_24; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_679 = io_ren_br_tags_0_valid ? _GEN_295 : br_snapshots_7_24; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_680 = io_ren_br_tags_0_valid ? _GEN_296 : br_snapshots_8_24; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_681 = io_ren_br_tags_0_valid ? _GEN_297 : br_snapshots_9_24; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_682 = io_ren_br_tags_0_valid ? _GEN_298 : br_snapshots_10_24; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_683 = io_ren_br_tags_0_valid ? _GEN_299 : br_snapshots_11_24; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_684 = io_ren_br_tags_0_valid ? _GEN_300 : br_snapshots_0_25; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_685 = io_ren_br_tags_0_valid ? _GEN_301 : br_snapshots_1_25; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_686 = io_ren_br_tags_0_valid ? _GEN_302 : br_snapshots_2_25; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_687 = io_ren_br_tags_0_valid ? _GEN_303 : br_snapshots_3_25; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_688 = io_ren_br_tags_0_valid ? _GEN_304 : br_snapshots_4_25; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_689 = io_ren_br_tags_0_valid ? _GEN_305 : br_snapshots_5_25; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_690 = io_ren_br_tags_0_valid ? _GEN_306 : br_snapshots_6_25; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_691 = io_ren_br_tags_0_valid ? _GEN_307 : br_snapshots_7_25; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_692 = io_ren_br_tags_0_valid ? _GEN_308 : br_snapshots_8_25; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_693 = io_ren_br_tags_0_valid ? _GEN_309 : br_snapshots_9_25; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_694 = io_ren_br_tags_0_valid ? _GEN_310 : br_snapshots_10_25; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_695 = io_ren_br_tags_0_valid ? _GEN_311 : br_snapshots_11_25; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_696 = io_ren_br_tags_0_valid ? _GEN_312 : br_snapshots_0_26; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_697 = io_ren_br_tags_0_valid ? _GEN_313 : br_snapshots_1_26; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_698 = io_ren_br_tags_0_valid ? _GEN_314 : br_snapshots_2_26; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_699 = io_ren_br_tags_0_valid ? _GEN_315 : br_snapshots_3_26; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_700 = io_ren_br_tags_0_valid ? _GEN_316 : br_snapshots_4_26; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_701 = io_ren_br_tags_0_valid ? _GEN_317 : br_snapshots_5_26; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_702 = io_ren_br_tags_0_valid ? _GEN_318 : br_snapshots_6_26; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_703 = io_ren_br_tags_0_valid ? _GEN_319 : br_snapshots_7_26; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_704 = io_ren_br_tags_0_valid ? _GEN_320 : br_snapshots_8_26; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_705 = io_ren_br_tags_0_valid ? _GEN_321 : br_snapshots_9_26; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_706 = io_ren_br_tags_0_valid ? _GEN_322 : br_snapshots_10_26; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_707 = io_ren_br_tags_0_valid ? _GEN_323 : br_snapshots_11_26; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_708 = io_ren_br_tags_0_valid ? _GEN_324 : br_snapshots_0_27; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_709 = io_ren_br_tags_0_valid ? _GEN_325 : br_snapshots_1_27; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_710 = io_ren_br_tags_0_valid ? _GEN_326 : br_snapshots_2_27; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_711 = io_ren_br_tags_0_valid ? _GEN_327 : br_snapshots_3_27; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_712 = io_ren_br_tags_0_valid ? _GEN_328 : br_snapshots_4_27; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_713 = io_ren_br_tags_0_valid ? _GEN_329 : br_snapshots_5_27; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_714 = io_ren_br_tags_0_valid ? _GEN_330 : br_snapshots_6_27; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_715 = io_ren_br_tags_0_valid ? _GEN_331 : br_snapshots_7_27; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_716 = io_ren_br_tags_0_valid ? _GEN_332 : br_snapshots_8_27; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_717 = io_ren_br_tags_0_valid ? _GEN_333 : br_snapshots_9_27; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_718 = io_ren_br_tags_0_valid ? _GEN_334 : br_snapshots_10_27; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_719 = io_ren_br_tags_0_valid ? _GEN_335 : br_snapshots_11_27; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_720 = io_ren_br_tags_0_valid ? _GEN_336 : br_snapshots_0_28; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_721 = io_ren_br_tags_0_valid ? _GEN_337 : br_snapshots_1_28; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_722 = io_ren_br_tags_0_valid ? _GEN_338 : br_snapshots_2_28; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_723 = io_ren_br_tags_0_valid ? _GEN_339 : br_snapshots_3_28; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_724 = io_ren_br_tags_0_valid ? _GEN_340 : br_snapshots_4_28; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_725 = io_ren_br_tags_0_valid ? _GEN_341 : br_snapshots_5_28; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_726 = io_ren_br_tags_0_valid ? _GEN_342 : br_snapshots_6_28; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_727 = io_ren_br_tags_0_valid ? _GEN_343 : br_snapshots_7_28; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_728 = io_ren_br_tags_0_valid ? _GEN_344 : br_snapshots_8_28; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_729 = io_ren_br_tags_0_valid ? _GEN_345 : br_snapshots_9_28; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_730 = io_ren_br_tags_0_valid ? _GEN_346 : br_snapshots_10_28; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_731 = io_ren_br_tags_0_valid ? _GEN_347 : br_snapshots_11_28; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_732 = io_ren_br_tags_0_valid ? _GEN_348 : br_snapshots_0_29; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_733 = io_ren_br_tags_0_valid ? _GEN_349 : br_snapshots_1_29; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_734 = io_ren_br_tags_0_valid ? _GEN_350 : br_snapshots_2_29; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_735 = io_ren_br_tags_0_valid ? _GEN_351 : br_snapshots_3_29; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_736 = io_ren_br_tags_0_valid ? _GEN_352 : br_snapshots_4_29; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_737 = io_ren_br_tags_0_valid ? _GEN_353 : br_snapshots_5_29; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_738 = io_ren_br_tags_0_valid ? _GEN_354 : br_snapshots_6_29; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_739 = io_ren_br_tags_0_valid ? _GEN_355 : br_snapshots_7_29; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_740 = io_ren_br_tags_0_valid ? _GEN_356 : br_snapshots_8_29; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_741 = io_ren_br_tags_0_valid ? _GEN_357 : br_snapshots_9_29; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_742 = io_ren_br_tags_0_valid ? _GEN_358 : br_snapshots_10_29; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_743 = io_ren_br_tags_0_valid ? _GEN_359 : br_snapshots_11_29; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_744 = io_ren_br_tags_0_valid ? _GEN_360 : br_snapshots_0_30; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_745 = io_ren_br_tags_0_valid ? _GEN_361 : br_snapshots_1_30; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_746 = io_ren_br_tags_0_valid ? _GEN_362 : br_snapshots_2_30; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_747 = io_ren_br_tags_0_valid ? _GEN_363 : br_snapshots_3_30; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_748 = io_ren_br_tags_0_valid ? _GEN_364 : br_snapshots_4_30; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_749 = io_ren_br_tags_0_valid ? _GEN_365 : br_snapshots_5_30; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_750 = io_ren_br_tags_0_valid ? _GEN_366 : br_snapshots_6_30; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_751 = io_ren_br_tags_0_valid ? _GEN_367 : br_snapshots_7_30; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_752 = io_ren_br_tags_0_valid ? _GEN_368 : br_snapshots_8_30; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_753 = io_ren_br_tags_0_valid ? _GEN_369 : br_snapshots_9_30; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_754 = io_ren_br_tags_0_valid ? _GEN_370 : br_snapshots_10_30; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_755 = io_ren_br_tags_0_valid ? _GEN_371 : br_snapshots_11_30; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_756 = io_ren_br_tags_0_valid ? _GEN_372 : br_snapshots_0_31; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_757 = io_ren_br_tags_0_valid ? _GEN_373 : br_snapshots_1_31; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_758 = io_ren_br_tags_0_valid ? _GEN_374 : br_snapshots_2_31; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_759 = io_ren_br_tags_0_valid ? _GEN_375 : br_snapshots_3_31; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_760 = io_ren_br_tags_0_valid ? _GEN_376 : br_snapshots_4_31; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_761 = io_ren_br_tags_0_valid ? _GEN_377 : br_snapshots_5_31; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_762 = io_ren_br_tags_0_valid ? _GEN_378 : br_snapshots_6_31; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_763 = io_ren_br_tags_0_valid ? _GEN_379 : br_snapshots_7_31; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_764 = io_ren_br_tags_0_valid ? _GEN_380 : br_snapshots_8_31; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_765 = io_ren_br_tags_0_valid ? _GEN_381 : br_snapshots_9_31; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_766 = io_ren_br_tags_0_valid ? _GEN_382 : br_snapshots_10_31; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_767 = io_ren_br_tags_0_valid ? _GEN_383 : br_snapshots_11_31; // @[rename-maptable.scala 132:36 rename-maptable.scala 79:25]
  wire [5:0] _GEN_1549 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_1 : br_snapshots_0_1; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1550 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_1 : _GEN_1549; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1551 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_1 : _GEN_1550; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1552 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_1 : _GEN_1551; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1553 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_1 : _GEN_1552; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1554 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_1 : _GEN_1553; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1555 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_1 : _GEN_1554; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1556 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_1 : _GEN_1555; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1557 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_1 : _GEN_1556; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1558 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_1 : _GEN_1557; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1561 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_2 : br_snapshots_0_2; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1562 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_2 : _GEN_1561; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1563 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_2 : _GEN_1562; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1564 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_2 : _GEN_1563; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1565 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_2 : _GEN_1564; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1566 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_2 : _GEN_1565; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1567 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_2 : _GEN_1566; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1568 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_2 : _GEN_1567; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1569 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_2 : _GEN_1568; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1570 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_2 : _GEN_1569; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1573 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_3 : br_snapshots_0_3; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1574 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_3 : _GEN_1573; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1575 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_3 : _GEN_1574; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1576 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_3 : _GEN_1575; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1577 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_3 : _GEN_1576; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1578 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_3 : _GEN_1577; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1579 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_3 : _GEN_1578; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1580 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_3 : _GEN_1579; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1581 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_3 : _GEN_1580; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1582 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_3 : _GEN_1581; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1585 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_4 : br_snapshots_0_4; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1586 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_4 : _GEN_1585; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1587 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_4 : _GEN_1586; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1588 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_4 : _GEN_1587; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1589 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_4 : _GEN_1588; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1590 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_4 : _GEN_1589; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1591 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_4 : _GEN_1590; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1592 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_4 : _GEN_1591; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1593 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_4 : _GEN_1592; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1594 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_4 : _GEN_1593; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1597 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_5 : br_snapshots_0_5; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1598 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_5 : _GEN_1597; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1599 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_5 : _GEN_1598; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1600 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_5 : _GEN_1599; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1601 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_5 : _GEN_1600; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1602 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_5 : _GEN_1601; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1603 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_5 : _GEN_1602; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1604 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_5 : _GEN_1603; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1605 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_5 : _GEN_1604; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1606 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_5 : _GEN_1605; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1609 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_6 : br_snapshots_0_6; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1610 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_6 : _GEN_1609; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1611 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_6 : _GEN_1610; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1612 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_6 : _GEN_1611; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1613 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_6 : _GEN_1612; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1614 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_6 : _GEN_1613; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1615 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_6 : _GEN_1614; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1616 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_6 : _GEN_1615; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1617 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_6 : _GEN_1616; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1618 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_6 : _GEN_1617; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1621 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_7 : br_snapshots_0_7; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1622 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_7 : _GEN_1621; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1623 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_7 : _GEN_1622; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1624 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_7 : _GEN_1623; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1625 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_7 : _GEN_1624; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1626 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_7 : _GEN_1625; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1627 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_7 : _GEN_1626; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1628 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_7 : _GEN_1627; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1629 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_7 : _GEN_1628; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1630 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_7 : _GEN_1629; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1633 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_8 : br_snapshots_0_8; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1634 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_8 : _GEN_1633; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1635 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_8 : _GEN_1634; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1636 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_8 : _GEN_1635; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1637 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_8 : _GEN_1636; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1638 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_8 : _GEN_1637; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1639 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_8 : _GEN_1638; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1640 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_8 : _GEN_1639; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1641 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_8 : _GEN_1640; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1642 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_8 : _GEN_1641; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1645 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_9 : br_snapshots_0_9; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1646 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_9 : _GEN_1645; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1647 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_9 : _GEN_1646; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1648 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_9 : _GEN_1647; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1649 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_9 : _GEN_1648; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1650 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_9 : _GEN_1649; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1651 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_9 : _GEN_1650; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1652 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_9 : _GEN_1651; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1653 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_9 : _GEN_1652; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1654 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_9 : _GEN_1653; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1657 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_10 : br_snapshots_0_10; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1658 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_10 : _GEN_1657; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1659 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_10 : _GEN_1658; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1660 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_10 : _GEN_1659; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1661 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_10 : _GEN_1660; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1662 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_10 : _GEN_1661; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1663 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_10 : _GEN_1662; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1664 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_10 : _GEN_1663; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1665 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_10 : _GEN_1664; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1666 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_10 : _GEN_1665; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1669 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_11 : br_snapshots_0_11; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1670 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_11 : _GEN_1669; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1671 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_11 : _GEN_1670; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1672 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_11 : _GEN_1671; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1673 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_11 : _GEN_1672; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1674 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_11 : _GEN_1673; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1675 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_11 : _GEN_1674; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1676 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_11 : _GEN_1675; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1677 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_11 : _GEN_1676; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1678 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_11 : _GEN_1677; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1681 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_12 : br_snapshots_0_12; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1682 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_12 : _GEN_1681; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1683 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_12 : _GEN_1682; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1684 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_12 : _GEN_1683; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1685 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_12 : _GEN_1684; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1686 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_12 : _GEN_1685; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1687 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_12 : _GEN_1686; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1688 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_12 : _GEN_1687; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1689 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_12 : _GEN_1688; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1690 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_12 : _GEN_1689; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1693 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_13 : br_snapshots_0_13; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1694 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_13 : _GEN_1693; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1695 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_13 : _GEN_1694; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1696 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_13 : _GEN_1695; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1697 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_13 : _GEN_1696; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1698 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_13 : _GEN_1697; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1699 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_13 : _GEN_1698; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1700 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_13 : _GEN_1699; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1701 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_13 : _GEN_1700; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1702 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_13 : _GEN_1701; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1705 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_14 : br_snapshots_0_14; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1706 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_14 : _GEN_1705; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1707 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_14 : _GEN_1706; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1708 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_14 : _GEN_1707; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1709 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_14 : _GEN_1708; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1710 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_14 : _GEN_1709; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1711 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_14 : _GEN_1710; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1712 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_14 : _GEN_1711; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1713 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_14 : _GEN_1712; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1714 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_14 : _GEN_1713; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1717 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_15 : br_snapshots_0_15; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1718 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_15 : _GEN_1717; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1719 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_15 : _GEN_1718; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1720 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_15 : _GEN_1719; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1721 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_15 : _GEN_1720; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1722 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_15 : _GEN_1721; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1723 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_15 : _GEN_1722; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1724 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_15 : _GEN_1723; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1725 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_15 : _GEN_1724; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1726 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_15 : _GEN_1725; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1729 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_16 : br_snapshots_0_16; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1730 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_16 : _GEN_1729; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1731 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_16 : _GEN_1730; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1732 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_16 : _GEN_1731; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1733 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_16 : _GEN_1732; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1734 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_16 : _GEN_1733; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1735 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_16 : _GEN_1734; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1736 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_16 : _GEN_1735; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1737 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_16 : _GEN_1736; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1738 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_16 : _GEN_1737; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1741 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_17 : br_snapshots_0_17; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1742 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_17 : _GEN_1741; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1743 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_17 : _GEN_1742; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1744 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_17 : _GEN_1743; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1745 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_17 : _GEN_1744; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1746 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_17 : _GEN_1745; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1747 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_17 : _GEN_1746; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1748 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_17 : _GEN_1747; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1749 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_17 : _GEN_1748; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1750 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_17 : _GEN_1749; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1753 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_18 : br_snapshots_0_18; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1754 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_18 : _GEN_1753; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1755 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_18 : _GEN_1754; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1756 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_18 : _GEN_1755; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1757 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_18 : _GEN_1756; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1758 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_18 : _GEN_1757; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1759 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_18 : _GEN_1758; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1760 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_18 : _GEN_1759; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1761 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_18 : _GEN_1760; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1762 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_18 : _GEN_1761; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1765 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_19 : br_snapshots_0_19; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1766 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_19 : _GEN_1765; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1767 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_19 : _GEN_1766; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1768 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_19 : _GEN_1767; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1769 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_19 : _GEN_1768; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1770 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_19 : _GEN_1769; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1771 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_19 : _GEN_1770; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1772 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_19 : _GEN_1771; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1773 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_19 : _GEN_1772; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1774 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_19 : _GEN_1773; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1777 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_20 : br_snapshots_0_20; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1778 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_20 : _GEN_1777; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1779 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_20 : _GEN_1778; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1780 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_20 : _GEN_1779; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1781 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_20 : _GEN_1780; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1782 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_20 : _GEN_1781; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1783 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_20 : _GEN_1782; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1784 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_20 : _GEN_1783; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1785 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_20 : _GEN_1784; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1786 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_20 : _GEN_1785; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1789 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_21 : br_snapshots_0_21; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1790 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_21 : _GEN_1789; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1791 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_21 : _GEN_1790; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1792 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_21 : _GEN_1791; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1793 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_21 : _GEN_1792; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1794 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_21 : _GEN_1793; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1795 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_21 : _GEN_1794; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1796 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_21 : _GEN_1795; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1797 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_21 : _GEN_1796; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1798 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_21 : _GEN_1797; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1801 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_22 : br_snapshots_0_22; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1802 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_22 : _GEN_1801; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1803 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_22 : _GEN_1802; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1804 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_22 : _GEN_1803; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1805 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_22 : _GEN_1804; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1806 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_22 : _GEN_1805; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1807 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_22 : _GEN_1806; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1808 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_22 : _GEN_1807; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1809 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_22 : _GEN_1808; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1810 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_22 : _GEN_1809; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1813 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_23 : br_snapshots_0_23; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1814 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_23 : _GEN_1813; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1815 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_23 : _GEN_1814; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1816 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_23 : _GEN_1815; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1817 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_23 : _GEN_1816; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1818 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_23 : _GEN_1817; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1819 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_23 : _GEN_1818; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1820 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_23 : _GEN_1819; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1821 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_23 : _GEN_1820; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1822 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_23 : _GEN_1821; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1825 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_24 : br_snapshots_0_24; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1826 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_24 : _GEN_1825; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1827 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_24 : _GEN_1826; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1828 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_24 : _GEN_1827; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1829 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_24 : _GEN_1828; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1830 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_24 : _GEN_1829; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1831 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_24 : _GEN_1830; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1832 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_24 : _GEN_1831; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1833 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_24 : _GEN_1832; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1834 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_24 : _GEN_1833; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1837 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_25 : br_snapshots_0_25; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1838 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_25 : _GEN_1837; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1839 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_25 : _GEN_1838; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1840 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_25 : _GEN_1839; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1841 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_25 : _GEN_1840; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1842 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_25 : _GEN_1841; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1843 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_25 : _GEN_1842; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1844 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_25 : _GEN_1843; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1845 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_25 : _GEN_1844; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1846 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_25 : _GEN_1845; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1849 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_26 : br_snapshots_0_26; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1850 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_26 : _GEN_1849; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1851 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_26 : _GEN_1850; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1852 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_26 : _GEN_1851; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1853 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_26 : _GEN_1852; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1854 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_26 : _GEN_1853; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1855 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_26 : _GEN_1854; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1856 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_26 : _GEN_1855; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1857 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_26 : _GEN_1856; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1858 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_26 : _GEN_1857; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1861 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_27 : br_snapshots_0_27; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1862 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_27 : _GEN_1861; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1863 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_27 : _GEN_1862; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1864 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_27 : _GEN_1863; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1865 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_27 : _GEN_1864; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1866 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_27 : _GEN_1865; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1867 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_27 : _GEN_1866; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1868 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_27 : _GEN_1867; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1869 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_27 : _GEN_1868; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1870 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_27 : _GEN_1869; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1873 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_28 : br_snapshots_0_28; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1874 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_28 : _GEN_1873; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1875 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_28 : _GEN_1874; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1876 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_28 : _GEN_1875; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1877 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_28 : _GEN_1876; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1878 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_28 : _GEN_1877; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1879 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_28 : _GEN_1878; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1880 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_28 : _GEN_1879; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1881 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_28 : _GEN_1880; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1882 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_28 : _GEN_1881; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1885 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_29 : br_snapshots_0_29; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1886 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_29 : _GEN_1885; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1887 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_29 : _GEN_1886; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1888 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_29 : _GEN_1887; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1889 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_29 : _GEN_1888; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1890 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_29 : _GEN_1889; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1891 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_29 : _GEN_1890; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1892 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_29 : _GEN_1891; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1893 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_29 : _GEN_1892; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1894 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_29 : _GEN_1893; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1897 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_30 : br_snapshots_0_30; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1898 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_30 : _GEN_1897; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1899 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_30 : _GEN_1898; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1900 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_30 : _GEN_1899; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1901 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_30 : _GEN_1900; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1902 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_30 : _GEN_1901; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1903 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_30 : _GEN_1902; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1904 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_30 : _GEN_1903; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1905 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_30 : _GEN_1904; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1906 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_30 : _GEN_1905; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1909 = 4'h1 == io_brupdate_b2_uop_br_tag ? br_snapshots_1_31 : br_snapshots_0_31; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1910 = 4'h2 == io_brupdate_b2_uop_br_tag ? br_snapshots_2_31 : _GEN_1909; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1911 = 4'h3 == io_brupdate_b2_uop_br_tag ? br_snapshots_3_31 : _GEN_1910; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1912 = 4'h4 == io_brupdate_b2_uop_br_tag ? br_snapshots_4_31 : _GEN_1911; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1913 = 4'h5 == io_brupdate_b2_uop_br_tag ? br_snapshots_5_31 : _GEN_1912; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1914 = 4'h6 == io_brupdate_b2_uop_br_tag ? br_snapshots_6_31 : _GEN_1913; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1915 = 4'h7 == io_brupdate_b2_uop_br_tag ? br_snapshots_7_31 : _GEN_1914; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1916 = 4'h8 == io_brupdate_b2_uop_br_tag ? br_snapshots_8_31 : _GEN_1915; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1917 = 4'h9 == io_brupdate_b2_uop_br_tag ? br_snapshots_9_31 : _GEN_1916; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_1918 = 4'ha == io_brupdate_b2_uop_br_tag ? br_snapshots_10_31 : _GEN_1917; // @[rename-maptable.scala 148:15 rename-maptable.scala 148:15]
  wire [5:0] _GEN_2369 = 5'h1 == io_map_reqs_0_lrs1[4:0] ? map_table_1 : map_table_0; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2370 = 5'h2 == io_map_reqs_0_lrs1[4:0] ? map_table_2 : _GEN_2369; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2371 = 5'h3 == io_map_reqs_0_lrs1[4:0] ? map_table_3 : _GEN_2370; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2372 = 5'h4 == io_map_reqs_0_lrs1[4:0] ? map_table_4 : _GEN_2371; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2373 = 5'h5 == io_map_reqs_0_lrs1[4:0] ? map_table_5 : _GEN_2372; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2374 = 5'h6 == io_map_reqs_0_lrs1[4:0] ? map_table_6 : _GEN_2373; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2375 = 5'h7 == io_map_reqs_0_lrs1[4:0] ? map_table_7 : _GEN_2374; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2376 = 5'h8 == io_map_reqs_0_lrs1[4:0] ? map_table_8 : _GEN_2375; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2377 = 5'h9 == io_map_reqs_0_lrs1[4:0] ? map_table_9 : _GEN_2376; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2378 = 5'ha == io_map_reqs_0_lrs1[4:0] ? map_table_10 : _GEN_2377; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2379 = 5'hb == io_map_reqs_0_lrs1[4:0] ? map_table_11 : _GEN_2378; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2380 = 5'hc == io_map_reqs_0_lrs1[4:0] ? map_table_12 : _GEN_2379; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2381 = 5'hd == io_map_reqs_0_lrs1[4:0] ? map_table_13 : _GEN_2380; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2382 = 5'he == io_map_reqs_0_lrs1[4:0] ? map_table_14 : _GEN_2381; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2383 = 5'hf == io_map_reqs_0_lrs1[4:0] ? map_table_15 : _GEN_2382; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2384 = 5'h10 == io_map_reqs_0_lrs1[4:0] ? map_table_16 : _GEN_2383; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2385 = 5'h11 == io_map_reqs_0_lrs1[4:0] ? map_table_17 : _GEN_2384; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2386 = 5'h12 == io_map_reqs_0_lrs1[4:0] ? map_table_18 : _GEN_2385; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2387 = 5'h13 == io_map_reqs_0_lrs1[4:0] ? map_table_19 : _GEN_2386; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2388 = 5'h14 == io_map_reqs_0_lrs1[4:0] ? map_table_20 : _GEN_2387; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2389 = 5'h15 == io_map_reqs_0_lrs1[4:0] ? map_table_21 : _GEN_2388; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2390 = 5'h16 == io_map_reqs_0_lrs1[4:0] ? map_table_22 : _GEN_2389; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2391 = 5'h17 == io_map_reqs_0_lrs1[4:0] ? map_table_23 : _GEN_2390; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2392 = 5'h18 == io_map_reqs_0_lrs1[4:0] ? map_table_24 : _GEN_2391; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2393 = 5'h19 == io_map_reqs_0_lrs1[4:0] ? map_table_25 : _GEN_2392; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2394 = 5'h1a == io_map_reqs_0_lrs1[4:0] ? map_table_26 : _GEN_2393; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2395 = 5'h1b == io_map_reqs_0_lrs1[4:0] ? map_table_27 : _GEN_2394; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2396 = 5'h1c == io_map_reqs_0_lrs1[4:0] ? map_table_28 : _GEN_2395; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2397 = 5'h1d == io_map_reqs_0_lrs1[4:0] ? map_table_29 : _GEN_2396; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2398 = 5'h1e == io_map_reqs_0_lrs1[4:0] ? map_table_30 : _GEN_2397; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  wire [5:0] _GEN_2401 = 5'h1 == io_map_reqs_0_lrs2[4:0] ? map_table_1 : map_table_0; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2402 = 5'h2 == io_map_reqs_0_lrs2[4:0] ? map_table_2 : _GEN_2401; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2403 = 5'h3 == io_map_reqs_0_lrs2[4:0] ? map_table_3 : _GEN_2402; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2404 = 5'h4 == io_map_reqs_0_lrs2[4:0] ? map_table_4 : _GEN_2403; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2405 = 5'h5 == io_map_reqs_0_lrs2[4:0] ? map_table_5 : _GEN_2404; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2406 = 5'h6 == io_map_reqs_0_lrs2[4:0] ? map_table_6 : _GEN_2405; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2407 = 5'h7 == io_map_reqs_0_lrs2[4:0] ? map_table_7 : _GEN_2406; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2408 = 5'h8 == io_map_reqs_0_lrs2[4:0] ? map_table_8 : _GEN_2407; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2409 = 5'h9 == io_map_reqs_0_lrs2[4:0] ? map_table_9 : _GEN_2408; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2410 = 5'ha == io_map_reqs_0_lrs2[4:0] ? map_table_10 : _GEN_2409; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2411 = 5'hb == io_map_reqs_0_lrs2[4:0] ? map_table_11 : _GEN_2410; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2412 = 5'hc == io_map_reqs_0_lrs2[4:0] ? map_table_12 : _GEN_2411; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2413 = 5'hd == io_map_reqs_0_lrs2[4:0] ? map_table_13 : _GEN_2412; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2414 = 5'he == io_map_reqs_0_lrs2[4:0] ? map_table_14 : _GEN_2413; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2415 = 5'hf == io_map_reqs_0_lrs2[4:0] ? map_table_15 : _GEN_2414; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2416 = 5'h10 == io_map_reqs_0_lrs2[4:0] ? map_table_16 : _GEN_2415; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2417 = 5'h11 == io_map_reqs_0_lrs2[4:0] ? map_table_17 : _GEN_2416; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2418 = 5'h12 == io_map_reqs_0_lrs2[4:0] ? map_table_18 : _GEN_2417; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2419 = 5'h13 == io_map_reqs_0_lrs2[4:0] ? map_table_19 : _GEN_2418; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2420 = 5'h14 == io_map_reqs_0_lrs2[4:0] ? map_table_20 : _GEN_2419; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2421 = 5'h15 == io_map_reqs_0_lrs2[4:0] ? map_table_21 : _GEN_2420; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2422 = 5'h16 == io_map_reqs_0_lrs2[4:0] ? map_table_22 : _GEN_2421; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2423 = 5'h17 == io_map_reqs_0_lrs2[4:0] ? map_table_23 : _GEN_2422; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2424 = 5'h18 == io_map_reqs_0_lrs2[4:0] ? map_table_24 : _GEN_2423; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2425 = 5'h19 == io_map_reqs_0_lrs2[4:0] ? map_table_25 : _GEN_2424; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2426 = 5'h1a == io_map_reqs_0_lrs2[4:0] ? map_table_26 : _GEN_2425; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2427 = 5'h1b == io_map_reqs_0_lrs2[4:0] ? map_table_27 : _GEN_2426; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2428 = 5'h1c == io_map_reqs_0_lrs2[4:0] ? map_table_28 : _GEN_2427; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2429 = 5'h1d == io_map_reqs_0_lrs2[4:0] ? map_table_29 : _GEN_2428; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2430 = 5'h1e == io_map_reqs_0_lrs2[4:0] ? map_table_30 : _GEN_2429; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  wire [5:0] _GEN_2465 = 5'h1 == io_map_reqs_0_ldst[4:0] ? map_table_1 : map_table_0; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2466 = 5'h2 == io_map_reqs_0_ldst[4:0] ? map_table_2 : _GEN_2465; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2467 = 5'h3 == io_map_reqs_0_ldst[4:0] ? map_table_3 : _GEN_2466; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2468 = 5'h4 == io_map_reqs_0_ldst[4:0] ? map_table_4 : _GEN_2467; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2469 = 5'h5 == io_map_reqs_0_ldst[4:0] ? map_table_5 : _GEN_2468; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2470 = 5'h6 == io_map_reqs_0_ldst[4:0] ? map_table_6 : _GEN_2469; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2471 = 5'h7 == io_map_reqs_0_ldst[4:0] ? map_table_7 : _GEN_2470; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2472 = 5'h8 == io_map_reqs_0_ldst[4:0] ? map_table_8 : _GEN_2471; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2473 = 5'h9 == io_map_reqs_0_ldst[4:0] ? map_table_9 : _GEN_2472; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2474 = 5'ha == io_map_reqs_0_ldst[4:0] ? map_table_10 : _GEN_2473; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2475 = 5'hb == io_map_reqs_0_ldst[4:0] ? map_table_11 : _GEN_2474; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2476 = 5'hc == io_map_reqs_0_ldst[4:0] ? map_table_12 : _GEN_2475; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2477 = 5'hd == io_map_reqs_0_ldst[4:0] ? map_table_13 : _GEN_2476; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2478 = 5'he == io_map_reqs_0_ldst[4:0] ? map_table_14 : _GEN_2477; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2479 = 5'hf == io_map_reqs_0_ldst[4:0] ? map_table_15 : _GEN_2478; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2480 = 5'h10 == io_map_reqs_0_ldst[4:0] ? map_table_16 : _GEN_2479; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2481 = 5'h11 == io_map_reqs_0_ldst[4:0] ? map_table_17 : _GEN_2480; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2482 = 5'h12 == io_map_reqs_0_ldst[4:0] ? map_table_18 : _GEN_2481; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2483 = 5'h13 == io_map_reqs_0_ldst[4:0] ? map_table_19 : _GEN_2482; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2484 = 5'h14 == io_map_reqs_0_ldst[4:0] ? map_table_20 : _GEN_2483; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2485 = 5'h15 == io_map_reqs_0_ldst[4:0] ? map_table_21 : _GEN_2484; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2486 = 5'h16 == io_map_reqs_0_ldst[4:0] ? map_table_22 : _GEN_2485; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2487 = 5'h17 == io_map_reqs_0_ldst[4:0] ? map_table_23 : _GEN_2486; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2488 = 5'h18 == io_map_reqs_0_ldst[4:0] ? map_table_24 : _GEN_2487; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2489 = 5'h19 == io_map_reqs_0_ldst[4:0] ? map_table_25 : _GEN_2488; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2490 = 5'h1a == io_map_reqs_0_ldst[4:0] ? map_table_26 : _GEN_2489; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2491 = 5'h1b == io_map_reqs_0_ldst[4:0] ? map_table_27 : _GEN_2490; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2492 = 5'h1c == io_map_reqs_0_ldst[4:0] ? map_table_28 : _GEN_2491; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2493 = 5'h1d == io_map_reqs_0_ldst[4:0] ? map_table_29 : _GEN_2492; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2494 = 5'h1e == io_map_reqs_0_ldst[4:0] ? map_table_30 : _GEN_2493; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  wire [5:0] _GEN_2497 = 5'h1 == io_map_reqs_1_lrs1[4:0] ? map_table_1 : map_table_0; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2498 = 5'h2 == io_map_reqs_1_lrs1[4:0] ? map_table_2 : _GEN_2497; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2499 = 5'h3 == io_map_reqs_1_lrs1[4:0] ? map_table_3 : _GEN_2498; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2500 = 5'h4 == io_map_reqs_1_lrs1[4:0] ? map_table_4 : _GEN_2499; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2501 = 5'h5 == io_map_reqs_1_lrs1[4:0] ? map_table_5 : _GEN_2500; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2502 = 5'h6 == io_map_reqs_1_lrs1[4:0] ? map_table_6 : _GEN_2501; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2503 = 5'h7 == io_map_reqs_1_lrs1[4:0] ? map_table_7 : _GEN_2502; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2504 = 5'h8 == io_map_reqs_1_lrs1[4:0] ? map_table_8 : _GEN_2503; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2505 = 5'h9 == io_map_reqs_1_lrs1[4:0] ? map_table_9 : _GEN_2504; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2506 = 5'ha == io_map_reqs_1_lrs1[4:0] ? map_table_10 : _GEN_2505; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2507 = 5'hb == io_map_reqs_1_lrs1[4:0] ? map_table_11 : _GEN_2506; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2508 = 5'hc == io_map_reqs_1_lrs1[4:0] ? map_table_12 : _GEN_2507; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2509 = 5'hd == io_map_reqs_1_lrs1[4:0] ? map_table_13 : _GEN_2508; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2510 = 5'he == io_map_reqs_1_lrs1[4:0] ? map_table_14 : _GEN_2509; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2511 = 5'hf == io_map_reqs_1_lrs1[4:0] ? map_table_15 : _GEN_2510; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2512 = 5'h10 == io_map_reqs_1_lrs1[4:0] ? map_table_16 : _GEN_2511; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2513 = 5'h11 == io_map_reqs_1_lrs1[4:0] ? map_table_17 : _GEN_2512; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2514 = 5'h12 == io_map_reqs_1_lrs1[4:0] ? map_table_18 : _GEN_2513; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2515 = 5'h13 == io_map_reqs_1_lrs1[4:0] ? map_table_19 : _GEN_2514; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2516 = 5'h14 == io_map_reqs_1_lrs1[4:0] ? map_table_20 : _GEN_2515; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2517 = 5'h15 == io_map_reqs_1_lrs1[4:0] ? map_table_21 : _GEN_2516; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2518 = 5'h16 == io_map_reqs_1_lrs1[4:0] ? map_table_22 : _GEN_2517; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2519 = 5'h17 == io_map_reqs_1_lrs1[4:0] ? map_table_23 : _GEN_2518; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2520 = 5'h18 == io_map_reqs_1_lrs1[4:0] ? map_table_24 : _GEN_2519; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2521 = 5'h19 == io_map_reqs_1_lrs1[4:0] ? map_table_25 : _GEN_2520; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2522 = 5'h1a == io_map_reqs_1_lrs1[4:0] ? map_table_26 : _GEN_2521; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2523 = 5'h1b == io_map_reqs_1_lrs1[4:0] ? map_table_27 : _GEN_2522; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2524 = 5'h1c == io_map_reqs_1_lrs1[4:0] ? map_table_28 : _GEN_2523; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2525 = 5'h1d == io_map_reqs_1_lrs1[4:0] ? map_table_29 : _GEN_2524; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2526 = 5'h1e == io_map_reqs_1_lrs1[4:0] ? map_table_30 : _GEN_2525; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  wire [5:0] _GEN_2529 = 5'h1 == io_map_reqs_1_lrs2[4:0] ? map_table_1 : map_table_0; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2530 = 5'h2 == io_map_reqs_1_lrs2[4:0] ? map_table_2 : _GEN_2529; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2531 = 5'h3 == io_map_reqs_1_lrs2[4:0] ? map_table_3 : _GEN_2530; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2532 = 5'h4 == io_map_reqs_1_lrs2[4:0] ? map_table_4 : _GEN_2531; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2533 = 5'h5 == io_map_reqs_1_lrs2[4:0] ? map_table_5 : _GEN_2532; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2534 = 5'h6 == io_map_reqs_1_lrs2[4:0] ? map_table_6 : _GEN_2533; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2535 = 5'h7 == io_map_reqs_1_lrs2[4:0] ? map_table_7 : _GEN_2534; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2536 = 5'h8 == io_map_reqs_1_lrs2[4:0] ? map_table_8 : _GEN_2535; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2537 = 5'h9 == io_map_reqs_1_lrs2[4:0] ? map_table_9 : _GEN_2536; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2538 = 5'ha == io_map_reqs_1_lrs2[4:0] ? map_table_10 : _GEN_2537; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2539 = 5'hb == io_map_reqs_1_lrs2[4:0] ? map_table_11 : _GEN_2538; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2540 = 5'hc == io_map_reqs_1_lrs2[4:0] ? map_table_12 : _GEN_2539; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2541 = 5'hd == io_map_reqs_1_lrs2[4:0] ? map_table_13 : _GEN_2540; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2542 = 5'he == io_map_reqs_1_lrs2[4:0] ? map_table_14 : _GEN_2541; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2543 = 5'hf == io_map_reqs_1_lrs2[4:0] ? map_table_15 : _GEN_2542; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2544 = 5'h10 == io_map_reqs_1_lrs2[4:0] ? map_table_16 : _GEN_2543; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2545 = 5'h11 == io_map_reqs_1_lrs2[4:0] ? map_table_17 : _GEN_2544; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2546 = 5'h12 == io_map_reqs_1_lrs2[4:0] ? map_table_18 : _GEN_2545; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2547 = 5'h13 == io_map_reqs_1_lrs2[4:0] ? map_table_19 : _GEN_2546; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2548 = 5'h14 == io_map_reqs_1_lrs2[4:0] ? map_table_20 : _GEN_2547; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2549 = 5'h15 == io_map_reqs_1_lrs2[4:0] ? map_table_21 : _GEN_2548; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2550 = 5'h16 == io_map_reqs_1_lrs2[4:0] ? map_table_22 : _GEN_2549; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2551 = 5'h17 == io_map_reqs_1_lrs2[4:0] ? map_table_23 : _GEN_2550; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2552 = 5'h18 == io_map_reqs_1_lrs2[4:0] ? map_table_24 : _GEN_2551; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2553 = 5'h19 == io_map_reqs_1_lrs2[4:0] ? map_table_25 : _GEN_2552; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2554 = 5'h1a == io_map_reqs_1_lrs2[4:0] ? map_table_26 : _GEN_2553; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2555 = 5'h1b == io_map_reqs_1_lrs2[4:0] ? map_table_27 : _GEN_2554; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2556 = 5'h1c == io_map_reqs_1_lrs2[4:0] ? map_table_28 : _GEN_2555; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2557 = 5'h1d == io_map_reqs_1_lrs2[4:0] ? map_table_29 : _GEN_2556; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2558 = 5'h1e == io_map_reqs_1_lrs2[4:0] ? map_table_30 : _GEN_2557; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  wire [5:0] _GEN_2593 = 5'h1 == io_map_reqs_1_ldst[4:0] ? map_table_1 : map_table_0; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2594 = 5'h2 == io_map_reqs_1_ldst[4:0] ? map_table_2 : _GEN_2593; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2595 = 5'h3 == io_map_reqs_1_ldst[4:0] ? map_table_3 : _GEN_2594; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2596 = 5'h4 == io_map_reqs_1_ldst[4:0] ? map_table_4 : _GEN_2595; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2597 = 5'h5 == io_map_reqs_1_ldst[4:0] ? map_table_5 : _GEN_2596; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2598 = 5'h6 == io_map_reqs_1_ldst[4:0] ? map_table_6 : _GEN_2597; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2599 = 5'h7 == io_map_reqs_1_ldst[4:0] ? map_table_7 : _GEN_2598; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2600 = 5'h8 == io_map_reqs_1_ldst[4:0] ? map_table_8 : _GEN_2599; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2601 = 5'h9 == io_map_reqs_1_ldst[4:0] ? map_table_9 : _GEN_2600; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2602 = 5'ha == io_map_reqs_1_ldst[4:0] ? map_table_10 : _GEN_2601; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2603 = 5'hb == io_map_reqs_1_ldst[4:0] ? map_table_11 : _GEN_2602; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2604 = 5'hc == io_map_reqs_1_ldst[4:0] ? map_table_12 : _GEN_2603; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2605 = 5'hd == io_map_reqs_1_ldst[4:0] ? map_table_13 : _GEN_2604; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2606 = 5'he == io_map_reqs_1_ldst[4:0] ? map_table_14 : _GEN_2605; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2607 = 5'hf == io_map_reqs_1_ldst[4:0] ? map_table_15 : _GEN_2606; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2608 = 5'h10 == io_map_reqs_1_ldst[4:0] ? map_table_16 : _GEN_2607; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2609 = 5'h11 == io_map_reqs_1_ldst[4:0] ? map_table_17 : _GEN_2608; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2610 = 5'h12 == io_map_reqs_1_ldst[4:0] ? map_table_18 : _GEN_2609; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2611 = 5'h13 == io_map_reqs_1_ldst[4:0] ? map_table_19 : _GEN_2610; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2612 = 5'h14 == io_map_reqs_1_ldst[4:0] ? map_table_20 : _GEN_2611; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2613 = 5'h15 == io_map_reqs_1_ldst[4:0] ? map_table_21 : _GEN_2612; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2614 = 5'h16 == io_map_reqs_1_ldst[4:0] ? map_table_22 : _GEN_2613; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2615 = 5'h17 == io_map_reqs_1_ldst[4:0] ? map_table_23 : _GEN_2614; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2616 = 5'h18 == io_map_reqs_1_ldst[4:0] ? map_table_24 : _GEN_2615; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2617 = 5'h19 == io_map_reqs_1_ldst[4:0] ? map_table_25 : _GEN_2616; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2618 = 5'h1a == io_map_reqs_1_ldst[4:0] ? map_table_26 : _GEN_2617; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2619 = 5'h1b == io_map_reqs_1_ldst[4:0] ? map_table_27 : _GEN_2618; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2620 = 5'h1c == io_map_reqs_1_ldst[4:0] ? map_table_28 : _GEN_2619; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2621 = 5'h1d == io_map_reqs_1_ldst[4:0] ? map_table_29 : _GEN_2620; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire [5:0] _GEN_2622 = 5'h1e == io_map_reqs_1_ldst[4:0] ? map_table_30 : _GEN_2621; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  wire  _T_565 = map_table_15 == io_remap_reqs_0_pdst; // @[rename-maptable.scala 176:38]
  wire  _T_597 = map_table_0 == io_remap_reqs_0_pdst | map_table_1 == io_remap_reqs_0_pdst | map_table_2 ==
    io_remap_reqs_0_pdst | map_table_3 == io_remap_reqs_0_pdst | map_table_4 == io_remap_reqs_0_pdst | map_table_5 ==
    io_remap_reqs_0_pdst | map_table_6 == io_remap_reqs_0_pdst | map_table_7 == io_remap_reqs_0_pdst | map_table_8 ==
    io_remap_reqs_0_pdst | map_table_9 == io_remap_reqs_0_pdst | map_table_10 == io_remap_reqs_0_pdst | map_table_11 ==
    io_remap_reqs_0_pdst | map_table_12 == io_remap_reqs_0_pdst | map_table_13 == io_remap_reqs_0_pdst | map_table_14
     == io_remap_reqs_0_pdst | _T_565; // @[rename-maptable.scala 176:38]
  wire  _T_612 = _T_597 | map_table_16 == io_remap_reqs_0_pdst | map_table_17 == io_remap_reqs_0_pdst | map_table_18 ==
    io_remap_reqs_0_pdst | map_table_19 == io_remap_reqs_0_pdst | map_table_20 == io_remap_reqs_0_pdst | map_table_21
     == io_remap_reqs_0_pdst | map_table_22 == io_remap_reqs_0_pdst | map_table_23 == io_remap_reqs_0_pdst |
    map_table_24 == io_remap_reqs_0_pdst | map_table_25 == io_remap_reqs_0_pdst | map_table_26 == io_remap_reqs_0_pdst
     | map_table_27 == io_remap_reqs_0_pdst | map_table_28 == io_remap_reqs_0_pdst | map_table_29 ==
    io_remap_reqs_0_pdst | map_table_30 == io_remap_reqs_0_pdst; // @[rename-maptable.scala 176:38]
  wire  _T_638 = map_table_15 == io_remap_reqs_1_pdst; // @[rename-maptable.scala 176:38]
  wire  _T_670 = map_table_0 == io_remap_reqs_1_pdst | map_table_1 == io_remap_reqs_1_pdst | map_table_2 ==
    io_remap_reqs_1_pdst | map_table_3 == io_remap_reqs_1_pdst | map_table_4 == io_remap_reqs_1_pdst | map_table_5 ==
    io_remap_reqs_1_pdst | map_table_6 == io_remap_reqs_1_pdst | map_table_7 == io_remap_reqs_1_pdst | map_table_8 ==
    io_remap_reqs_1_pdst | map_table_9 == io_remap_reqs_1_pdst | map_table_10 == io_remap_reqs_1_pdst | map_table_11 ==
    io_remap_reqs_1_pdst | map_table_12 == io_remap_reqs_1_pdst | map_table_13 == io_remap_reqs_1_pdst | map_table_14
     == io_remap_reqs_1_pdst | _T_638; // @[rename-maptable.scala 176:38]
  wire  _T_685 = _T_670 | map_table_16 == io_remap_reqs_1_pdst | map_table_17 == io_remap_reqs_1_pdst | map_table_18 ==
    io_remap_reqs_1_pdst | map_table_19 == io_remap_reqs_1_pdst | map_table_20 == io_remap_reqs_1_pdst | map_table_21
     == io_remap_reqs_1_pdst | map_table_22 == io_remap_reqs_1_pdst | map_table_23 == io_remap_reqs_1_pdst |
    map_table_24 == io_remap_reqs_1_pdst | map_table_25 == io_remap_reqs_1_pdst | map_table_26 == io_remap_reqs_1_pdst
     | map_table_27 == io_remap_reqs_1_pdst | map_table_28 == io_remap_reqs_1_pdst | map_table_29 ==
    io_remap_reqs_1_pdst | map_table_30 == io_remap_reqs_1_pdst; // @[rename-maptable.scala 176:38]
  assign io_map_resps_0_prs1_valid = ~io_flush; // @[rename-maptable.scala 156:35]
  assign io_map_resps_0_prs1_bits = 5'h1f == io_map_reqs_0_lrs1[4:0] ? map_table_31 : _GEN_2398; // @[rename-maptable.scala 161:37 rename-maptable.scala 161:37]
  assign io_map_resps_0_prs2_valid = ~io_flush; // @[rename-maptable.scala 157:35]
  assign io_map_resps_0_prs2_bits = 5'h1f == io_map_reqs_0_lrs2[4:0] ? map_table_31 : _GEN_2430; // @[rename-maptable.scala 163:36 rename-maptable.scala 163:36]
  assign io_map_resps_0_prs3_valid = 1'h0;
  assign io_map_resps_0_prs3_bits = 6'h0;
  assign io_map_resps_0_stale_pdst_valid = ~io_flush; // @[rename-maptable.scala 159:41]
  assign io_map_resps_0_stale_pdst_bits = 5'h1f == io_map_reqs_0_ldst[4:0] ? map_table_31 : _GEN_2494; // @[rename-maptable.scala 167:37 rename-maptable.scala 167:37]
  assign io_map_resps_1_prs1_valid = ~io_flush; // @[rename-maptable.scala 156:35]
  assign io_map_resps_1_prs1_bits = 5'h1f == io_map_reqs_1_lrs1[4:0] ? map_table_31 : _GEN_2526; // @[rename-maptable.scala 162:10 rename-maptable.scala 162:10]
  assign io_map_resps_1_prs2_valid = ~io_flush; // @[rename-maptable.scala 157:35]
  assign io_map_resps_1_prs2_bits = 5'h1f == io_map_reqs_1_lrs2[4:0] ? map_table_31 : _GEN_2558; // @[rename-maptable.scala 164:10 rename-maptable.scala 164:10]
  assign io_map_resps_1_prs3_valid = 1'h0;
  assign io_map_resps_1_prs3_bits = 6'h0;
  assign io_map_resps_1_stale_pdst_valid = ~io_flush; // @[rename-maptable.scala 159:41]
  assign io_map_resps_1_stale_pdst_bits = 5'h1f == io_map_reqs_1_ldst[4:0] ? map_table_31 : _GEN_2622; // @[rename-maptable.scala 168:10 rename-maptable.scala 168:10]
  assign io_commit_bits = _T_391 | _T_359; // @[rename-maptable.scala 112:104]
  always @(posedge clock) begin
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_0 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_0 <= commit_map_table_0; // @[rename-maptable.scala 139:20]
    end else begin
      map_table_0 <= 6'h0;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_1 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_1 <= commit_map_table_1; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_1 <= br_snapshots_11_1; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_1 <= _GEN_1558;
      end
    end else if (remap_ldsts_oh_1[1]) begin // @[rename-maptable.scala 122:70]
      map_table_1 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_1 <= remap_table_1_1;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_2 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_2 <= commit_map_table_2; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_2 <= br_snapshots_11_2; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_2 <= _GEN_1570;
      end
    end else if (remap_ldsts_oh_1[2]) begin // @[rename-maptable.scala 122:70]
      map_table_2 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_2 <= remap_table_1_2;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_3 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_3 <= commit_map_table_3; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_3 <= br_snapshots_11_3; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_3 <= _GEN_1582;
      end
    end else if (remap_ldsts_oh_1[3]) begin // @[rename-maptable.scala 122:70]
      map_table_3 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_3 <= remap_table_1_3;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_4 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_4 <= commit_map_table_4; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_4 <= br_snapshots_11_4; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_4 <= _GEN_1594;
      end
    end else if (remap_ldsts_oh_1[4]) begin // @[rename-maptable.scala 122:70]
      map_table_4 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_4 <= remap_table_1_4;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_5 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_5 <= commit_map_table_5; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_5 <= br_snapshots_11_5; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_5 <= _GEN_1606;
      end
    end else if (remap_ldsts_oh_1[5]) begin // @[rename-maptable.scala 122:70]
      map_table_5 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_5 <= remap_table_1_5;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_6 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_6 <= commit_map_table_6; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_6 <= br_snapshots_11_6; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_6 <= _GEN_1618;
      end
    end else if (remap_ldsts_oh_1[6]) begin // @[rename-maptable.scala 122:70]
      map_table_6 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_6 <= remap_table_1_6;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_7 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_7 <= commit_map_table_7; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_7 <= br_snapshots_11_7; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_7 <= _GEN_1630;
      end
    end else if (remap_ldsts_oh_1[7]) begin // @[rename-maptable.scala 122:70]
      map_table_7 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_7 <= remap_table_1_7;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_8 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_8 <= commit_map_table_8; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_8 <= br_snapshots_11_8; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_8 <= _GEN_1642;
      end
    end else if (remap_ldsts_oh_1[8]) begin // @[rename-maptable.scala 122:70]
      map_table_8 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_8 <= remap_table_1_8;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_9 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_9 <= commit_map_table_9; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_9 <= br_snapshots_11_9; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_9 <= _GEN_1654;
      end
    end else if (remap_ldsts_oh_1[9]) begin // @[rename-maptable.scala 122:70]
      map_table_9 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_9 <= remap_table_1_9;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_10 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_10 <= commit_map_table_10; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_10 <= br_snapshots_11_10; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_10 <= _GEN_1666;
      end
    end else if (remap_ldsts_oh_1[10]) begin // @[rename-maptable.scala 122:70]
      map_table_10 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_10 <= remap_table_1_10;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_11 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_11 <= commit_map_table_11; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_11 <= br_snapshots_11_11; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_11 <= _GEN_1678;
      end
    end else if (remap_ldsts_oh_1[11]) begin // @[rename-maptable.scala 122:70]
      map_table_11 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_11 <= remap_table_1_11;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_12 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_12 <= commit_map_table_12; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_12 <= br_snapshots_11_12; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_12 <= _GEN_1690;
      end
    end else if (remap_ldsts_oh_1[12]) begin // @[rename-maptable.scala 122:70]
      map_table_12 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_12 <= remap_table_1_12;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_13 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_13 <= commit_map_table_13; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_13 <= br_snapshots_11_13; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_13 <= _GEN_1702;
      end
    end else if (remap_ldsts_oh_1[13]) begin // @[rename-maptable.scala 122:70]
      map_table_13 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_13 <= remap_table_1_13;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_14 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_14 <= commit_map_table_14; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_14 <= br_snapshots_11_14; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_14 <= _GEN_1714;
      end
    end else if (remap_ldsts_oh_1[14]) begin // @[rename-maptable.scala 122:70]
      map_table_14 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_14 <= remap_table_1_14;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_15 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_15 <= commit_map_table_15; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_15 <= br_snapshots_11_15; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_15 <= _GEN_1726;
      end
    end else if (remap_ldsts_oh_1[15]) begin // @[rename-maptable.scala 122:70]
      map_table_15 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_15 <= remap_table_1_15;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_16 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_16 <= commit_map_table_16; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_16 <= br_snapshots_11_16; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_16 <= _GEN_1738;
      end
    end else if (remap_ldsts_oh_1[16]) begin // @[rename-maptable.scala 122:70]
      map_table_16 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_16 <= remap_table_1_16;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_17 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_17 <= commit_map_table_17; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_17 <= br_snapshots_11_17; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_17 <= _GEN_1750;
      end
    end else if (remap_ldsts_oh_1[17]) begin // @[rename-maptable.scala 122:70]
      map_table_17 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_17 <= remap_table_1_17;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_18 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_18 <= commit_map_table_18; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_18 <= br_snapshots_11_18; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_18 <= _GEN_1762;
      end
    end else if (remap_ldsts_oh_1[18]) begin // @[rename-maptable.scala 122:70]
      map_table_18 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_18 <= remap_table_1_18;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_19 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_19 <= commit_map_table_19; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_19 <= br_snapshots_11_19; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_19 <= _GEN_1774;
      end
    end else if (remap_ldsts_oh_1[19]) begin // @[rename-maptable.scala 122:70]
      map_table_19 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_19 <= remap_table_1_19;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_20 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_20 <= commit_map_table_20; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_20 <= br_snapshots_11_20; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_20 <= _GEN_1786;
      end
    end else if (remap_ldsts_oh_1[20]) begin // @[rename-maptable.scala 122:70]
      map_table_20 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_20 <= remap_table_1_20;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_21 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_21 <= commit_map_table_21; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_21 <= br_snapshots_11_21; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_21 <= _GEN_1798;
      end
    end else if (remap_ldsts_oh_1[21]) begin // @[rename-maptable.scala 122:70]
      map_table_21 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_21 <= remap_table_1_21;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_22 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_22 <= commit_map_table_22; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_22 <= br_snapshots_11_22; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_22 <= _GEN_1810;
      end
    end else if (remap_ldsts_oh_1[22]) begin // @[rename-maptable.scala 122:70]
      map_table_22 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_22 <= remap_table_1_22;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_23 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_23 <= commit_map_table_23; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_23 <= br_snapshots_11_23; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_23 <= _GEN_1822;
      end
    end else if (remap_ldsts_oh_1[23]) begin // @[rename-maptable.scala 122:70]
      map_table_23 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_23 <= remap_table_1_23;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_24 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_24 <= commit_map_table_24; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_24 <= br_snapshots_11_24; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_24 <= _GEN_1834;
      end
    end else if (remap_ldsts_oh_1[24]) begin // @[rename-maptable.scala 122:70]
      map_table_24 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_24 <= remap_table_1_24;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_25 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_25 <= commit_map_table_25; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_25 <= br_snapshots_11_25; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_25 <= _GEN_1846;
      end
    end else if (remap_ldsts_oh_1[25]) begin // @[rename-maptable.scala 122:70]
      map_table_25 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_25 <= remap_table_1_25;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_26 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_26 <= commit_map_table_26; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_26 <= br_snapshots_11_26; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_26 <= _GEN_1858;
      end
    end else if (remap_ldsts_oh_1[26]) begin // @[rename-maptable.scala 122:70]
      map_table_26 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_26 <= remap_table_1_26;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_27 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_27 <= commit_map_table_27; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_27 <= br_snapshots_11_27; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_27 <= _GEN_1870;
      end
    end else if (remap_ldsts_oh_1[27]) begin // @[rename-maptable.scala 122:70]
      map_table_27 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_27 <= remap_table_1_27;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_28 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_28 <= commit_map_table_28; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_28 <= br_snapshots_11_28; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_28 <= _GEN_1882;
      end
    end else if (remap_ldsts_oh_1[28]) begin // @[rename-maptable.scala 122:70]
      map_table_28 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_28 <= remap_table_1_28;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_29 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_29 <= commit_map_table_29; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_29 <= br_snapshots_11_29; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_29 <= _GEN_1894;
      end
    end else if (remap_ldsts_oh_1[29]) begin // @[rename-maptable.scala 122:70]
      map_table_29 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_29 <= remap_table_1_29;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_30 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_30 <= commit_map_table_30; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_30 <= br_snapshots_11_30; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_30 <= _GEN_1906;
      end
    end else if (remap_ldsts_oh_1[30]) begin // @[rename-maptable.scala 122:70]
      map_table_30 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_30 <= remap_table_1_30;
    end
    if (reset) begin // @[rename-maptable.scala 77:26]
      map_table_31 <= 6'h0; // @[rename-maptable.scala 77:26]
    end else if (io_flush) begin // @[rename-maptable.scala 137:19]
      map_table_31 <= commit_map_table_31; // @[rename-maptable.scala 139:20]
    end else if (io_brupdate_b2_mispredict) begin // @[rename-maptable.scala 146:42]
      if (4'hb == io_brupdate_b2_uop_br_tag) begin // @[rename-maptable.scala 148:15]
        map_table_31 <= br_snapshots_11_31; // @[rename-maptable.scala 148:15]
      end else begin
        map_table_31 <= _GEN_1918;
      end
    end else if (remap_ldsts_oh_1[31]) begin // @[rename-maptable.scala 122:70]
      map_table_31 <= io_remap_reqs_1_pdst;
    end else begin
      map_table_31 <= remap_table_1_31;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_0 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[0]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_0 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[0]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_0 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_1 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[1]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_1 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[1]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_1 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_2 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[2]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_2 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[2]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_2 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_3 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[3]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_3 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[3]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_3 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_4 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[4]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_4 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[4]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_4 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_5 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[5]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_5 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[5]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_5 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_6 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[6]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_6 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[6]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_6 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_7 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[7]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_7 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[7]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_7 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_8 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[8]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_8 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[8]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_8 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_9 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[9]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_9 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[9]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_9 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_10 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[10]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_10 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[10]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_10 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_11 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[11]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_11 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[11]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_11 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_12 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[12]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_12 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[12]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_12 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_13 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[13]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_13 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[13]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_13 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_14 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[14]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_14 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[14]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_14 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_15 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[15]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_15 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[15]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_15 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_16 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[16]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_16 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[16]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_16 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_17 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[17]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_17 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[17]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_17 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_18 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[18]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_18 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[18]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_18 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_19 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[19]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_19 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[19]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_19 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_20 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[20]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_20 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[20]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_20 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_21 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[21]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_21 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[21]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_21 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_22 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[22]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_22 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[22]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_22 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_23 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[23]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_23 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[23]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_23 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_24 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[24]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_24 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[24]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_24 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_25 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[25]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_25 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[25]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_25 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_26 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[26]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_26 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[26]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_26 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_27 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[27]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_27 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[27]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_27 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_28 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[28]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_28 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[28]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_28 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_29 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[29]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_29 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[29]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_29 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_30 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[30]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_30 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[30]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_30 <= io_commit_regs_0_pdst;
    end
    if (reset) begin // @[rename-maptable.scala 78:33]
      commit_map_table_31 <= 6'h0; // @[rename-maptable.scala 78:33]
    end else if (rrat_ldsts_oh_1[31]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_31 <= io_commit_regs_1_pdst;
    end else if (rrat_ldsts_oh_0[31]) begin // @[rename-maptable.scala 95:75]
      commit_map_table_31 <= io_commit_regs_0_pdst;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_1 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[1]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_1 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_1 <= remap_table_1_1;
        end
      end else begin
        br_snapshots_0_1 <= _GEN_396;
      end
    end else begin
      br_snapshots_0_1 <= _GEN_396;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_2 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[2]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_2 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_2 <= remap_table_1_2;
        end
      end else begin
        br_snapshots_0_2 <= _GEN_408;
      end
    end else begin
      br_snapshots_0_2 <= _GEN_408;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_3 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[3]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_3 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_3 <= remap_table_1_3;
        end
      end else begin
        br_snapshots_0_3 <= _GEN_420;
      end
    end else begin
      br_snapshots_0_3 <= _GEN_420;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_4 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[4]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_4 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_4 <= remap_table_1_4;
        end
      end else begin
        br_snapshots_0_4 <= _GEN_432;
      end
    end else begin
      br_snapshots_0_4 <= _GEN_432;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_5 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[5]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_5 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_5 <= remap_table_1_5;
        end
      end else begin
        br_snapshots_0_5 <= _GEN_444;
      end
    end else begin
      br_snapshots_0_5 <= _GEN_444;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_6 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[6]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_6 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_6 <= remap_table_1_6;
        end
      end else begin
        br_snapshots_0_6 <= _GEN_456;
      end
    end else begin
      br_snapshots_0_6 <= _GEN_456;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_7 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[7]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_7 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_7 <= remap_table_1_7;
        end
      end else begin
        br_snapshots_0_7 <= _GEN_468;
      end
    end else begin
      br_snapshots_0_7 <= _GEN_468;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_8 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[8]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_8 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_8 <= remap_table_1_8;
        end
      end else begin
        br_snapshots_0_8 <= _GEN_480;
      end
    end else begin
      br_snapshots_0_8 <= _GEN_480;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_9 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[9]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_9 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_9 <= remap_table_1_9;
        end
      end else begin
        br_snapshots_0_9 <= _GEN_492;
      end
    end else begin
      br_snapshots_0_9 <= _GEN_492;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_10 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[10]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_10 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_10 <= remap_table_1_10;
        end
      end else begin
        br_snapshots_0_10 <= _GEN_504;
      end
    end else begin
      br_snapshots_0_10 <= _GEN_504;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_11 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[11]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_11 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_11 <= remap_table_1_11;
        end
      end else begin
        br_snapshots_0_11 <= _GEN_516;
      end
    end else begin
      br_snapshots_0_11 <= _GEN_516;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_12 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[12]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_12 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_12 <= remap_table_1_12;
        end
      end else begin
        br_snapshots_0_12 <= _GEN_528;
      end
    end else begin
      br_snapshots_0_12 <= _GEN_528;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_13 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[13]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_13 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_13 <= remap_table_1_13;
        end
      end else begin
        br_snapshots_0_13 <= _GEN_540;
      end
    end else begin
      br_snapshots_0_13 <= _GEN_540;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_14 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[14]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_14 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_14 <= remap_table_1_14;
        end
      end else begin
        br_snapshots_0_14 <= _GEN_552;
      end
    end else begin
      br_snapshots_0_14 <= _GEN_552;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_15 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[15]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_15 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_15 <= remap_table_1_15;
        end
      end else begin
        br_snapshots_0_15 <= _GEN_564;
      end
    end else begin
      br_snapshots_0_15 <= _GEN_564;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_16 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[16]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_16 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_16 <= remap_table_1_16;
        end
      end else begin
        br_snapshots_0_16 <= _GEN_576;
      end
    end else begin
      br_snapshots_0_16 <= _GEN_576;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_17 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[17]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_17 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_17 <= remap_table_1_17;
        end
      end else begin
        br_snapshots_0_17 <= _GEN_588;
      end
    end else begin
      br_snapshots_0_17 <= _GEN_588;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_18 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[18]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_18 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_18 <= remap_table_1_18;
        end
      end else begin
        br_snapshots_0_18 <= _GEN_600;
      end
    end else begin
      br_snapshots_0_18 <= _GEN_600;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_19 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[19]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_19 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_19 <= remap_table_1_19;
        end
      end else begin
        br_snapshots_0_19 <= _GEN_612;
      end
    end else begin
      br_snapshots_0_19 <= _GEN_612;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_20 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[20]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_20 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_20 <= remap_table_1_20;
        end
      end else begin
        br_snapshots_0_20 <= _GEN_624;
      end
    end else begin
      br_snapshots_0_20 <= _GEN_624;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_21 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[21]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_21 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_21 <= remap_table_1_21;
        end
      end else begin
        br_snapshots_0_21 <= _GEN_636;
      end
    end else begin
      br_snapshots_0_21 <= _GEN_636;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_22 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[22]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_22 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_22 <= remap_table_1_22;
        end
      end else begin
        br_snapshots_0_22 <= _GEN_648;
      end
    end else begin
      br_snapshots_0_22 <= _GEN_648;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_23 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[23]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_23 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_23 <= remap_table_1_23;
        end
      end else begin
        br_snapshots_0_23 <= _GEN_660;
      end
    end else begin
      br_snapshots_0_23 <= _GEN_660;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_24 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[24]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_24 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_24 <= remap_table_1_24;
        end
      end else begin
        br_snapshots_0_24 <= _GEN_672;
      end
    end else begin
      br_snapshots_0_24 <= _GEN_672;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_25 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[25]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_25 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_25 <= remap_table_1_25;
        end
      end else begin
        br_snapshots_0_25 <= _GEN_684;
      end
    end else begin
      br_snapshots_0_25 <= _GEN_684;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_26 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[26]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_26 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_26 <= remap_table_1_26;
        end
      end else begin
        br_snapshots_0_26 <= _GEN_696;
      end
    end else begin
      br_snapshots_0_26 <= _GEN_696;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_27 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[27]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_27 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_27 <= remap_table_1_27;
        end
      end else begin
        br_snapshots_0_27 <= _GEN_708;
      end
    end else begin
      br_snapshots_0_27 <= _GEN_708;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_28 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[28]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_28 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_28 <= remap_table_1_28;
        end
      end else begin
        br_snapshots_0_28 <= _GEN_720;
      end
    end else begin
      br_snapshots_0_28 <= _GEN_720;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_29 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[29]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_29 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_29 <= remap_table_1_29;
        end
      end else begin
        br_snapshots_0_29 <= _GEN_732;
      end
    end else begin
      br_snapshots_0_29 <= _GEN_732;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_30 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[30]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_30 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_30 <= remap_table_1_30;
        end
      end else begin
        br_snapshots_0_30 <= _GEN_744;
      end
    end else begin
      br_snapshots_0_30 <= _GEN_744;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_0_31 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h0 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[31]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_0_31 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_0_31 <= remap_table_1_31;
        end
      end else begin
        br_snapshots_0_31 <= _GEN_756;
      end
    end else begin
      br_snapshots_0_31 <= _GEN_756;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_1 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[1]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_1 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_1 <= remap_table_1_1;
        end
      end else begin
        br_snapshots_1_1 <= _GEN_397;
      end
    end else begin
      br_snapshots_1_1 <= _GEN_397;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_2 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[2]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_2 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_2 <= remap_table_1_2;
        end
      end else begin
        br_snapshots_1_2 <= _GEN_409;
      end
    end else begin
      br_snapshots_1_2 <= _GEN_409;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_3 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[3]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_3 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_3 <= remap_table_1_3;
        end
      end else begin
        br_snapshots_1_3 <= _GEN_421;
      end
    end else begin
      br_snapshots_1_3 <= _GEN_421;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_4 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[4]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_4 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_4 <= remap_table_1_4;
        end
      end else begin
        br_snapshots_1_4 <= _GEN_433;
      end
    end else begin
      br_snapshots_1_4 <= _GEN_433;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_5 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[5]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_5 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_5 <= remap_table_1_5;
        end
      end else begin
        br_snapshots_1_5 <= _GEN_445;
      end
    end else begin
      br_snapshots_1_5 <= _GEN_445;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_6 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[6]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_6 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_6 <= remap_table_1_6;
        end
      end else begin
        br_snapshots_1_6 <= _GEN_457;
      end
    end else begin
      br_snapshots_1_6 <= _GEN_457;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_7 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[7]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_7 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_7 <= remap_table_1_7;
        end
      end else begin
        br_snapshots_1_7 <= _GEN_469;
      end
    end else begin
      br_snapshots_1_7 <= _GEN_469;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_8 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[8]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_8 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_8 <= remap_table_1_8;
        end
      end else begin
        br_snapshots_1_8 <= _GEN_481;
      end
    end else begin
      br_snapshots_1_8 <= _GEN_481;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_9 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[9]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_9 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_9 <= remap_table_1_9;
        end
      end else begin
        br_snapshots_1_9 <= _GEN_493;
      end
    end else begin
      br_snapshots_1_9 <= _GEN_493;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_10 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[10]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_10 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_10 <= remap_table_1_10;
        end
      end else begin
        br_snapshots_1_10 <= _GEN_505;
      end
    end else begin
      br_snapshots_1_10 <= _GEN_505;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_11 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[11]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_11 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_11 <= remap_table_1_11;
        end
      end else begin
        br_snapshots_1_11 <= _GEN_517;
      end
    end else begin
      br_snapshots_1_11 <= _GEN_517;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_12 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[12]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_12 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_12 <= remap_table_1_12;
        end
      end else begin
        br_snapshots_1_12 <= _GEN_529;
      end
    end else begin
      br_snapshots_1_12 <= _GEN_529;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_13 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[13]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_13 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_13 <= remap_table_1_13;
        end
      end else begin
        br_snapshots_1_13 <= _GEN_541;
      end
    end else begin
      br_snapshots_1_13 <= _GEN_541;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_14 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[14]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_14 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_14 <= remap_table_1_14;
        end
      end else begin
        br_snapshots_1_14 <= _GEN_553;
      end
    end else begin
      br_snapshots_1_14 <= _GEN_553;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_15 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[15]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_15 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_15 <= remap_table_1_15;
        end
      end else begin
        br_snapshots_1_15 <= _GEN_565;
      end
    end else begin
      br_snapshots_1_15 <= _GEN_565;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_16 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[16]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_16 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_16 <= remap_table_1_16;
        end
      end else begin
        br_snapshots_1_16 <= _GEN_577;
      end
    end else begin
      br_snapshots_1_16 <= _GEN_577;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_17 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[17]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_17 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_17 <= remap_table_1_17;
        end
      end else begin
        br_snapshots_1_17 <= _GEN_589;
      end
    end else begin
      br_snapshots_1_17 <= _GEN_589;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_18 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[18]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_18 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_18 <= remap_table_1_18;
        end
      end else begin
        br_snapshots_1_18 <= _GEN_601;
      end
    end else begin
      br_snapshots_1_18 <= _GEN_601;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_19 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[19]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_19 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_19 <= remap_table_1_19;
        end
      end else begin
        br_snapshots_1_19 <= _GEN_613;
      end
    end else begin
      br_snapshots_1_19 <= _GEN_613;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_20 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[20]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_20 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_20 <= remap_table_1_20;
        end
      end else begin
        br_snapshots_1_20 <= _GEN_625;
      end
    end else begin
      br_snapshots_1_20 <= _GEN_625;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_21 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[21]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_21 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_21 <= remap_table_1_21;
        end
      end else begin
        br_snapshots_1_21 <= _GEN_637;
      end
    end else begin
      br_snapshots_1_21 <= _GEN_637;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_22 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[22]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_22 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_22 <= remap_table_1_22;
        end
      end else begin
        br_snapshots_1_22 <= _GEN_649;
      end
    end else begin
      br_snapshots_1_22 <= _GEN_649;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_23 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[23]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_23 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_23 <= remap_table_1_23;
        end
      end else begin
        br_snapshots_1_23 <= _GEN_661;
      end
    end else begin
      br_snapshots_1_23 <= _GEN_661;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_24 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[24]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_24 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_24 <= remap_table_1_24;
        end
      end else begin
        br_snapshots_1_24 <= _GEN_673;
      end
    end else begin
      br_snapshots_1_24 <= _GEN_673;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_25 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[25]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_25 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_25 <= remap_table_1_25;
        end
      end else begin
        br_snapshots_1_25 <= _GEN_685;
      end
    end else begin
      br_snapshots_1_25 <= _GEN_685;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_26 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[26]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_26 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_26 <= remap_table_1_26;
        end
      end else begin
        br_snapshots_1_26 <= _GEN_697;
      end
    end else begin
      br_snapshots_1_26 <= _GEN_697;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_27 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[27]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_27 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_27 <= remap_table_1_27;
        end
      end else begin
        br_snapshots_1_27 <= _GEN_709;
      end
    end else begin
      br_snapshots_1_27 <= _GEN_709;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_28 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[28]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_28 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_28 <= remap_table_1_28;
        end
      end else begin
        br_snapshots_1_28 <= _GEN_721;
      end
    end else begin
      br_snapshots_1_28 <= _GEN_721;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_29 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[29]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_29 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_29 <= remap_table_1_29;
        end
      end else begin
        br_snapshots_1_29 <= _GEN_733;
      end
    end else begin
      br_snapshots_1_29 <= _GEN_733;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_30 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[30]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_30 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_30 <= remap_table_1_30;
        end
      end else begin
        br_snapshots_1_30 <= _GEN_745;
      end
    end else begin
      br_snapshots_1_30 <= _GEN_745;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_1_31 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h1 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[31]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_1_31 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_1_31 <= remap_table_1_31;
        end
      end else begin
        br_snapshots_1_31 <= _GEN_757;
      end
    end else begin
      br_snapshots_1_31 <= _GEN_757;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_1 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[1]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_1 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_1 <= remap_table_1_1;
        end
      end else begin
        br_snapshots_2_1 <= _GEN_398;
      end
    end else begin
      br_snapshots_2_1 <= _GEN_398;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_2 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[2]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_2 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_2 <= remap_table_1_2;
        end
      end else begin
        br_snapshots_2_2 <= _GEN_410;
      end
    end else begin
      br_snapshots_2_2 <= _GEN_410;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_3 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[3]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_3 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_3 <= remap_table_1_3;
        end
      end else begin
        br_snapshots_2_3 <= _GEN_422;
      end
    end else begin
      br_snapshots_2_3 <= _GEN_422;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_4 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[4]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_4 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_4 <= remap_table_1_4;
        end
      end else begin
        br_snapshots_2_4 <= _GEN_434;
      end
    end else begin
      br_snapshots_2_4 <= _GEN_434;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_5 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[5]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_5 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_5 <= remap_table_1_5;
        end
      end else begin
        br_snapshots_2_5 <= _GEN_446;
      end
    end else begin
      br_snapshots_2_5 <= _GEN_446;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_6 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[6]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_6 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_6 <= remap_table_1_6;
        end
      end else begin
        br_snapshots_2_6 <= _GEN_458;
      end
    end else begin
      br_snapshots_2_6 <= _GEN_458;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_7 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[7]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_7 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_7 <= remap_table_1_7;
        end
      end else begin
        br_snapshots_2_7 <= _GEN_470;
      end
    end else begin
      br_snapshots_2_7 <= _GEN_470;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_8 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[8]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_8 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_8 <= remap_table_1_8;
        end
      end else begin
        br_snapshots_2_8 <= _GEN_482;
      end
    end else begin
      br_snapshots_2_8 <= _GEN_482;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_9 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[9]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_9 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_9 <= remap_table_1_9;
        end
      end else begin
        br_snapshots_2_9 <= _GEN_494;
      end
    end else begin
      br_snapshots_2_9 <= _GEN_494;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_10 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[10]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_10 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_10 <= remap_table_1_10;
        end
      end else begin
        br_snapshots_2_10 <= _GEN_506;
      end
    end else begin
      br_snapshots_2_10 <= _GEN_506;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_11 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[11]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_11 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_11 <= remap_table_1_11;
        end
      end else begin
        br_snapshots_2_11 <= _GEN_518;
      end
    end else begin
      br_snapshots_2_11 <= _GEN_518;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_12 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[12]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_12 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_12 <= remap_table_1_12;
        end
      end else begin
        br_snapshots_2_12 <= _GEN_530;
      end
    end else begin
      br_snapshots_2_12 <= _GEN_530;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_13 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[13]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_13 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_13 <= remap_table_1_13;
        end
      end else begin
        br_snapshots_2_13 <= _GEN_542;
      end
    end else begin
      br_snapshots_2_13 <= _GEN_542;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_14 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[14]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_14 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_14 <= remap_table_1_14;
        end
      end else begin
        br_snapshots_2_14 <= _GEN_554;
      end
    end else begin
      br_snapshots_2_14 <= _GEN_554;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_15 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[15]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_15 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_15 <= remap_table_1_15;
        end
      end else begin
        br_snapshots_2_15 <= _GEN_566;
      end
    end else begin
      br_snapshots_2_15 <= _GEN_566;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_16 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[16]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_16 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_16 <= remap_table_1_16;
        end
      end else begin
        br_snapshots_2_16 <= _GEN_578;
      end
    end else begin
      br_snapshots_2_16 <= _GEN_578;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_17 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[17]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_17 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_17 <= remap_table_1_17;
        end
      end else begin
        br_snapshots_2_17 <= _GEN_590;
      end
    end else begin
      br_snapshots_2_17 <= _GEN_590;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_18 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[18]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_18 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_18 <= remap_table_1_18;
        end
      end else begin
        br_snapshots_2_18 <= _GEN_602;
      end
    end else begin
      br_snapshots_2_18 <= _GEN_602;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_19 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[19]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_19 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_19 <= remap_table_1_19;
        end
      end else begin
        br_snapshots_2_19 <= _GEN_614;
      end
    end else begin
      br_snapshots_2_19 <= _GEN_614;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_20 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[20]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_20 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_20 <= remap_table_1_20;
        end
      end else begin
        br_snapshots_2_20 <= _GEN_626;
      end
    end else begin
      br_snapshots_2_20 <= _GEN_626;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_21 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[21]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_21 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_21 <= remap_table_1_21;
        end
      end else begin
        br_snapshots_2_21 <= _GEN_638;
      end
    end else begin
      br_snapshots_2_21 <= _GEN_638;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_22 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[22]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_22 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_22 <= remap_table_1_22;
        end
      end else begin
        br_snapshots_2_22 <= _GEN_650;
      end
    end else begin
      br_snapshots_2_22 <= _GEN_650;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_23 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[23]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_23 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_23 <= remap_table_1_23;
        end
      end else begin
        br_snapshots_2_23 <= _GEN_662;
      end
    end else begin
      br_snapshots_2_23 <= _GEN_662;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_24 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[24]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_24 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_24 <= remap_table_1_24;
        end
      end else begin
        br_snapshots_2_24 <= _GEN_674;
      end
    end else begin
      br_snapshots_2_24 <= _GEN_674;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_25 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[25]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_25 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_25 <= remap_table_1_25;
        end
      end else begin
        br_snapshots_2_25 <= _GEN_686;
      end
    end else begin
      br_snapshots_2_25 <= _GEN_686;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_26 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[26]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_26 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_26 <= remap_table_1_26;
        end
      end else begin
        br_snapshots_2_26 <= _GEN_698;
      end
    end else begin
      br_snapshots_2_26 <= _GEN_698;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_27 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[27]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_27 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_27 <= remap_table_1_27;
        end
      end else begin
        br_snapshots_2_27 <= _GEN_710;
      end
    end else begin
      br_snapshots_2_27 <= _GEN_710;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_28 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[28]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_28 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_28 <= remap_table_1_28;
        end
      end else begin
        br_snapshots_2_28 <= _GEN_722;
      end
    end else begin
      br_snapshots_2_28 <= _GEN_722;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_29 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[29]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_29 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_29 <= remap_table_1_29;
        end
      end else begin
        br_snapshots_2_29 <= _GEN_734;
      end
    end else begin
      br_snapshots_2_29 <= _GEN_734;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_30 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[30]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_30 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_30 <= remap_table_1_30;
        end
      end else begin
        br_snapshots_2_30 <= _GEN_746;
      end
    end else begin
      br_snapshots_2_30 <= _GEN_746;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_2_31 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h2 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[31]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_2_31 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_2_31 <= remap_table_1_31;
        end
      end else begin
        br_snapshots_2_31 <= _GEN_758;
      end
    end else begin
      br_snapshots_2_31 <= _GEN_758;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_1 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[1]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_1 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_1 <= remap_table_1_1;
        end
      end else begin
        br_snapshots_3_1 <= _GEN_399;
      end
    end else begin
      br_snapshots_3_1 <= _GEN_399;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_2 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[2]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_2 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_2 <= remap_table_1_2;
        end
      end else begin
        br_snapshots_3_2 <= _GEN_411;
      end
    end else begin
      br_snapshots_3_2 <= _GEN_411;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_3 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[3]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_3 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_3 <= remap_table_1_3;
        end
      end else begin
        br_snapshots_3_3 <= _GEN_423;
      end
    end else begin
      br_snapshots_3_3 <= _GEN_423;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_4 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[4]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_4 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_4 <= remap_table_1_4;
        end
      end else begin
        br_snapshots_3_4 <= _GEN_435;
      end
    end else begin
      br_snapshots_3_4 <= _GEN_435;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_5 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[5]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_5 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_5 <= remap_table_1_5;
        end
      end else begin
        br_snapshots_3_5 <= _GEN_447;
      end
    end else begin
      br_snapshots_3_5 <= _GEN_447;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_6 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[6]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_6 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_6 <= remap_table_1_6;
        end
      end else begin
        br_snapshots_3_6 <= _GEN_459;
      end
    end else begin
      br_snapshots_3_6 <= _GEN_459;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_7 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[7]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_7 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_7 <= remap_table_1_7;
        end
      end else begin
        br_snapshots_3_7 <= _GEN_471;
      end
    end else begin
      br_snapshots_3_7 <= _GEN_471;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_8 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[8]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_8 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_8 <= remap_table_1_8;
        end
      end else begin
        br_snapshots_3_8 <= _GEN_483;
      end
    end else begin
      br_snapshots_3_8 <= _GEN_483;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_9 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[9]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_9 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_9 <= remap_table_1_9;
        end
      end else begin
        br_snapshots_3_9 <= _GEN_495;
      end
    end else begin
      br_snapshots_3_9 <= _GEN_495;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_10 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[10]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_10 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_10 <= remap_table_1_10;
        end
      end else begin
        br_snapshots_3_10 <= _GEN_507;
      end
    end else begin
      br_snapshots_3_10 <= _GEN_507;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_11 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[11]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_11 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_11 <= remap_table_1_11;
        end
      end else begin
        br_snapshots_3_11 <= _GEN_519;
      end
    end else begin
      br_snapshots_3_11 <= _GEN_519;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_12 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[12]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_12 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_12 <= remap_table_1_12;
        end
      end else begin
        br_snapshots_3_12 <= _GEN_531;
      end
    end else begin
      br_snapshots_3_12 <= _GEN_531;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_13 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[13]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_13 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_13 <= remap_table_1_13;
        end
      end else begin
        br_snapshots_3_13 <= _GEN_543;
      end
    end else begin
      br_snapshots_3_13 <= _GEN_543;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_14 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[14]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_14 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_14 <= remap_table_1_14;
        end
      end else begin
        br_snapshots_3_14 <= _GEN_555;
      end
    end else begin
      br_snapshots_3_14 <= _GEN_555;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_15 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[15]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_15 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_15 <= remap_table_1_15;
        end
      end else begin
        br_snapshots_3_15 <= _GEN_567;
      end
    end else begin
      br_snapshots_3_15 <= _GEN_567;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_16 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[16]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_16 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_16 <= remap_table_1_16;
        end
      end else begin
        br_snapshots_3_16 <= _GEN_579;
      end
    end else begin
      br_snapshots_3_16 <= _GEN_579;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_17 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[17]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_17 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_17 <= remap_table_1_17;
        end
      end else begin
        br_snapshots_3_17 <= _GEN_591;
      end
    end else begin
      br_snapshots_3_17 <= _GEN_591;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_18 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[18]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_18 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_18 <= remap_table_1_18;
        end
      end else begin
        br_snapshots_3_18 <= _GEN_603;
      end
    end else begin
      br_snapshots_3_18 <= _GEN_603;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_19 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[19]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_19 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_19 <= remap_table_1_19;
        end
      end else begin
        br_snapshots_3_19 <= _GEN_615;
      end
    end else begin
      br_snapshots_3_19 <= _GEN_615;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_20 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[20]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_20 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_20 <= remap_table_1_20;
        end
      end else begin
        br_snapshots_3_20 <= _GEN_627;
      end
    end else begin
      br_snapshots_3_20 <= _GEN_627;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_21 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[21]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_21 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_21 <= remap_table_1_21;
        end
      end else begin
        br_snapshots_3_21 <= _GEN_639;
      end
    end else begin
      br_snapshots_3_21 <= _GEN_639;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_22 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[22]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_22 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_22 <= remap_table_1_22;
        end
      end else begin
        br_snapshots_3_22 <= _GEN_651;
      end
    end else begin
      br_snapshots_3_22 <= _GEN_651;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_23 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[23]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_23 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_23 <= remap_table_1_23;
        end
      end else begin
        br_snapshots_3_23 <= _GEN_663;
      end
    end else begin
      br_snapshots_3_23 <= _GEN_663;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_24 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[24]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_24 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_24 <= remap_table_1_24;
        end
      end else begin
        br_snapshots_3_24 <= _GEN_675;
      end
    end else begin
      br_snapshots_3_24 <= _GEN_675;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_25 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[25]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_25 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_25 <= remap_table_1_25;
        end
      end else begin
        br_snapshots_3_25 <= _GEN_687;
      end
    end else begin
      br_snapshots_3_25 <= _GEN_687;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_26 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[26]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_26 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_26 <= remap_table_1_26;
        end
      end else begin
        br_snapshots_3_26 <= _GEN_699;
      end
    end else begin
      br_snapshots_3_26 <= _GEN_699;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_27 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[27]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_27 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_27 <= remap_table_1_27;
        end
      end else begin
        br_snapshots_3_27 <= _GEN_711;
      end
    end else begin
      br_snapshots_3_27 <= _GEN_711;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_28 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[28]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_28 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_28 <= remap_table_1_28;
        end
      end else begin
        br_snapshots_3_28 <= _GEN_723;
      end
    end else begin
      br_snapshots_3_28 <= _GEN_723;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_29 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[29]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_29 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_29 <= remap_table_1_29;
        end
      end else begin
        br_snapshots_3_29 <= _GEN_735;
      end
    end else begin
      br_snapshots_3_29 <= _GEN_735;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_30 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[30]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_30 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_30 <= remap_table_1_30;
        end
      end else begin
        br_snapshots_3_30 <= _GEN_747;
      end
    end else begin
      br_snapshots_3_30 <= _GEN_747;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_3_31 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h3 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[31]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_3_31 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_3_31 <= remap_table_1_31;
        end
      end else begin
        br_snapshots_3_31 <= _GEN_759;
      end
    end else begin
      br_snapshots_3_31 <= _GEN_759;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_1 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[1]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_1 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_1 <= remap_table_1_1;
        end
      end else begin
        br_snapshots_4_1 <= _GEN_400;
      end
    end else begin
      br_snapshots_4_1 <= _GEN_400;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_2 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[2]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_2 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_2 <= remap_table_1_2;
        end
      end else begin
        br_snapshots_4_2 <= _GEN_412;
      end
    end else begin
      br_snapshots_4_2 <= _GEN_412;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_3 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[3]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_3 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_3 <= remap_table_1_3;
        end
      end else begin
        br_snapshots_4_3 <= _GEN_424;
      end
    end else begin
      br_snapshots_4_3 <= _GEN_424;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_4 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[4]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_4 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_4 <= remap_table_1_4;
        end
      end else begin
        br_snapshots_4_4 <= _GEN_436;
      end
    end else begin
      br_snapshots_4_4 <= _GEN_436;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_5 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[5]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_5 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_5 <= remap_table_1_5;
        end
      end else begin
        br_snapshots_4_5 <= _GEN_448;
      end
    end else begin
      br_snapshots_4_5 <= _GEN_448;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_6 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[6]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_6 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_6 <= remap_table_1_6;
        end
      end else begin
        br_snapshots_4_6 <= _GEN_460;
      end
    end else begin
      br_snapshots_4_6 <= _GEN_460;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_7 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[7]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_7 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_7 <= remap_table_1_7;
        end
      end else begin
        br_snapshots_4_7 <= _GEN_472;
      end
    end else begin
      br_snapshots_4_7 <= _GEN_472;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_8 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[8]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_8 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_8 <= remap_table_1_8;
        end
      end else begin
        br_snapshots_4_8 <= _GEN_484;
      end
    end else begin
      br_snapshots_4_8 <= _GEN_484;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_9 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[9]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_9 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_9 <= remap_table_1_9;
        end
      end else begin
        br_snapshots_4_9 <= _GEN_496;
      end
    end else begin
      br_snapshots_4_9 <= _GEN_496;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_10 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[10]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_10 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_10 <= remap_table_1_10;
        end
      end else begin
        br_snapshots_4_10 <= _GEN_508;
      end
    end else begin
      br_snapshots_4_10 <= _GEN_508;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_11 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[11]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_11 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_11 <= remap_table_1_11;
        end
      end else begin
        br_snapshots_4_11 <= _GEN_520;
      end
    end else begin
      br_snapshots_4_11 <= _GEN_520;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_12 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[12]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_12 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_12 <= remap_table_1_12;
        end
      end else begin
        br_snapshots_4_12 <= _GEN_532;
      end
    end else begin
      br_snapshots_4_12 <= _GEN_532;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_13 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[13]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_13 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_13 <= remap_table_1_13;
        end
      end else begin
        br_snapshots_4_13 <= _GEN_544;
      end
    end else begin
      br_snapshots_4_13 <= _GEN_544;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_14 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[14]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_14 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_14 <= remap_table_1_14;
        end
      end else begin
        br_snapshots_4_14 <= _GEN_556;
      end
    end else begin
      br_snapshots_4_14 <= _GEN_556;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_15 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[15]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_15 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_15 <= remap_table_1_15;
        end
      end else begin
        br_snapshots_4_15 <= _GEN_568;
      end
    end else begin
      br_snapshots_4_15 <= _GEN_568;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_16 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[16]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_16 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_16 <= remap_table_1_16;
        end
      end else begin
        br_snapshots_4_16 <= _GEN_580;
      end
    end else begin
      br_snapshots_4_16 <= _GEN_580;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_17 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[17]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_17 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_17 <= remap_table_1_17;
        end
      end else begin
        br_snapshots_4_17 <= _GEN_592;
      end
    end else begin
      br_snapshots_4_17 <= _GEN_592;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_18 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[18]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_18 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_18 <= remap_table_1_18;
        end
      end else begin
        br_snapshots_4_18 <= _GEN_604;
      end
    end else begin
      br_snapshots_4_18 <= _GEN_604;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_19 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[19]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_19 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_19 <= remap_table_1_19;
        end
      end else begin
        br_snapshots_4_19 <= _GEN_616;
      end
    end else begin
      br_snapshots_4_19 <= _GEN_616;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_20 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[20]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_20 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_20 <= remap_table_1_20;
        end
      end else begin
        br_snapshots_4_20 <= _GEN_628;
      end
    end else begin
      br_snapshots_4_20 <= _GEN_628;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_21 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[21]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_21 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_21 <= remap_table_1_21;
        end
      end else begin
        br_snapshots_4_21 <= _GEN_640;
      end
    end else begin
      br_snapshots_4_21 <= _GEN_640;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_22 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[22]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_22 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_22 <= remap_table_1_22;
        end
      end else begin
        br_snapshots_4_22 <= _GEN_652;
      end
    end else begin
      br_snapshots_4_22 <= _GEN_652;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_23 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[23]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_23 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_23 <= remap_table_1_23;
        end
      end else begin
        br_snapshots_4_23 <= _GEN_664;
      end
    end else begin
      br_snapshots_4_23 <= _GEN_664;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_24 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[24]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_24 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_24 <= remap_table_1_24;
        end
      end else begin
        br_snapshots_4_24 <= _GEN_676;
      end
    end else begin
      br_snapshots_4_24 <= _GEN_676;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_25 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[25]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_25 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_25 <= remap_table_1_25;
        end
      end else begin
        br_snapshots_4_25 <= _GEN_688;
      end
    end else begin
      br_snapshots_4_25 <= _GEN_688;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_26 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[26]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_26 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_26 <= remap_table_1_26;
        end
      end else begin
        br_snapshots_4_26 <= _GEN_700;
      end
    end else begin
      br_snapshots_4_26 <= _GEN_700;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_27 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[27]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_27 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_27 <= remap_table_1_27;
        end
      end else begin
        br_snapshots_4_27 <= _GEN_712;
      end
    end else begin
      br_snapshots_4_27 <= _GEN_712;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_28 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[28]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_28 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_28 <= remap_table_1_28;
        end
      end else begin
        br_snapshots_4_28 <= _GEN_724;
      end
    end else begin
      br_snapshots_4_28 <= _GEN_724;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_29 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[29]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_29 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_29 <= remap_table_1_29;
        end
      end else begin
        br_snapshots_4_29 <= _GEN_736;
      end
    end else begin
      br_snapshots_4_29 <= _GEN_736;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_30 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[30]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_30 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_30 <= remap_table_1_30;
        end
      end else begin
        br_snapshots_4_30 <= _GEN_748;
      end
    end else begin
      br_snapshots_4_30 <= _GEN_748;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_4_31 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h4 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[31]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_4_31 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_4_31 <= remap_table_1_31;
        end
      end else begin
        br_snapshots_4_31 <= _GEN_760;
      end
    end else begin
      br_snapshots_4_31 <= _GEN_760;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_1 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[1]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_1 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_1 <= remap_table_1_1;
        end
      end else begin
        br_snapshots_5_1 <= _GEN_401;
      end
    end else begin
      br_snapshots_5_1 <= _GEN_401;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_2 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[2]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_2 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_2 <= remap_table_1_2;
        end
      end else begin
        br_snapshots_5_2 <= _GEN_413;
      end
    end else begin
      br_snapshots_5_2 <= _GEN_413;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_3 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[3]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_3 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_3 <= remap_table_1_3;
        end
      end else begin
        br_snapshots_5_3 <= _GEN_425;
      end
    end else begin
      br_snapshots_5_3 <= _GEN_425;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_4 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[4]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_4 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_4 <= remap_table_1_4;
        end
      end else begin
        br_snapshots_5_4 <= _GEN_437;
      end
    end else begin
      br_snapshots_5_4 <= _GEN_437;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_5 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[5]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_5 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_5 <= remap_table_1_5;
        end
      end else begin
        br_snapshots_5_5 <= _GEN_449;
      end
    end else begin
      br_snapshots_5_5 <= _GEN_449;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_6 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[6]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_6 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_6 <= remap_table_1_6;
        end
      end else begin
        br_snapshots_5_6 <= _GEN_461;
      end
    end else begin
      br_snapshots_5_6 <= _GEN_461;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_7 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[7]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_7 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_7 <= remap_table_1_7;
        end
      end else begin
        br_snapshots_5_7 <= _GEN_473;
      end
    end else begin
      br_snapshots_5_7 <= _GEN_473;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_8 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[8]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_8 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_8 <= remap_table_1_8;
        end
      end else begin
        br_snapshots_5_8 <= _GEN_485;
      end
    end else begin
      br_snapshots_5_8 <= _GEN_485;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_9 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[9]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_9 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_9 <= remap_table_1_9;
        end
      end else begin
        br_snapshots_5_9 <= _GEN_497;
      end
    end else begin
      br_snapshots_5_9 <= _GEN_497;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_10 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[10]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_10 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_10 <= remap_table_1_10;
        end
      end else begin
        br_snapshots_5_10 <= _GEN_509;
      end
    end else begin
      br_snapshots_5_10 <= _GEN_509;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_11 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[11]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_11 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_11 <= remap_table_1_11;
        end
      end else begin
        br_snapshots_5_11 <= _GEN_521;
      end
    end else begin
      br_snapshots_5_11 <= _GEN_521;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_12 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[12]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_12 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_12 <= remap_table_1_12;
        end
      end else begin
        br_snapshots_5_12 <= _GEN_533;
      end
    end else begin
      br_snapshots_5_12 <= _GEN_533;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_13 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[13]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_13 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_13 <= remap_table_1_13;
        end
      end else begin
        br_snapshots_5_13 <= _GEN_545;
      end
    end else begin
      br_snapshots_5_13 <= _GEN_545;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_14 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[14]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_14 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_14 <= remap_table_1_14;
        end
      end else begin
        br_snapshots_5_14 <= _GEN_557;
      end
    end else begin
      br_snapshots_5_14 <= _GEN_557;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_15 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[15]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_15 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_15 <= remap_table_1_15;
        end
      end else begin
        br_snapshots_5_15 <= _GEN_569;
      end
    end else begin
      br_snapshots_5_15 <= _GEN_569;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_16 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[16]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_16 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_16 <= remap_table_1_16;
        end
      end else begin
        br_snapshots_5_16 <= _GEN_581;
      end
    end else begin
      br_snapshots_5_16 <= _GEN_581;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_17 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[17]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_17 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_17 <= remap_table_1_17;
        end
      end else begin
        br_snapshots_5_17 <= _GEN_593;
      end
    end else begin
      br_snapshots_5_17 <= _GEN_593;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_18 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[18]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_18 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_18 <= remap_table_1_18;
        end
      end else begin
        br_snapshots_5_18 <= _GEN_605;
      end
    end else begin
      br_snapshots_5_18 <= _GEN_605;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_19 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[19]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_19 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_19 <= remap_table_1_19;
        end
      end else begin
        br_snapshots_5_19 <= _GEN_617;
      end
    end else begin
      br_snapshots_5_19 <= _GEN_617;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_20 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[20]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_20 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_20 <= remap_table_1_20;
        end
      end else begin
        br_snapshots_5_20 <= _GEN_629;
      end
    end else begin
      br_snapshots_5_20 <= _GEN_629;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_21 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[21]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_21 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_21 <= remap_table_1_21;
        end
      end else begin
        br_snapshots_5_21 <= _GEN_641;
      end
    end else begin
      br_snapshots_5_21 <= _GEN_641;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_22 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[22]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_22 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_22 <= remap_table_1_22;
        end
      end else begin
        br_snapshots_5_22 <= _GEN_653;
      end
    end else begin
      br_snapshots_5_22 <= _GEN_653;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_23 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[23]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_23 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_23 <= remap_table_1_23;
        end
      end else begin
        br_snapshots_5_23 <= _GEN_665;
      end
    end else begin
      br_snapshots_5_23 <= _GEN_665;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_24 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[24]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_24 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_24 <= remap_table_1_24;
        end
      end else begin
        br_snapshots_5_24 <= _GEN_677;
      end
    end else begin
      br_snapshots_5_24 <= _GEN_677;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_25 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[25]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_25 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_25 <= remap_table_1_25;
        end
      end else begin
        br_snapshots_5_25 <= _GEN_689;
      end
    end else begin
      br_snapshots_5_25 <= _GEN_689;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_26 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[26]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_26 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_26 <= remap_table_1_26;
        end
      end else begin
        br_snapshots_5_26 <= _GEN_701;
      end
    end else begin
      br_snapshots_5_26 <= _GEN_701;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_27 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[27]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_27 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_27 <= remap_table_1_27;
        end
      end else begin
        br_snapshots_5_27 <= _GEN_713;
      end
    end else begin
      br_snapshots_5_27 <= _GEN_713;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_28 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[28]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_28 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_28 <= remap_table_1_28;
        end
      end else begin
        br_snapshots_5_28 <= _GEN_725;
      end
    end else begin
      br_snapshots_5_28 <= _GEN_725;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_29 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[29]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_29 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_29 <= remap_table_1_29;
        end
      end else begin
        br_snapshots_5_29 <= _GEN_737;
      end
    end else begin
      br_snapshots_5_29 <= _GEN_737;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_30 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[30]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_30 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_30 <= remap_table_1_30;
        end
      end else begin
        br_snapshots_5_30 <= _GEN_749;
      end
    end else begin
      br_snapshots_5_30 <= _GEN_749;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_5_31 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h5 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[31]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_5_31 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_5_31 <= remap_table_1_31;
        end
      end else begin
        br_snapshots_5_31 <= _GEN_761;
      end
    end else begin
      br_snapshots_5_31 <= _GEN_761;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_1 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[1]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_1 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_1 <= remap_table_1_1;
        end
      end else begin
        br_snapshots_6_1 <= _GEN_402;
      end
    end else begin
      br_snapshots_6_1 <= _GEN_402;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_2 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[2]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_2 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_2 <= remap_table_1_2;
        end
      end else begin
        br_snapshots_6_2 <= _GEN_414;
      end
    end else begin
      br_snapshots_6_2 <= _GEN_414;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_3 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[3]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_3 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_3 <= remap_table_1_3;
        end
      end else begin
        br_snapshots_6_3 <= _GEN_426;
      end
    end else begin
      br_snapshots_6_3 <= _GEN_426;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_4 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[4]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_4 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_4 <= remap_table_1_4;
        end
      end else begin
        br_snapshots_6_4 <= _GEN_438;
      end
    end else begin
      br_snapshots_6_4 <= _GEN_438;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_5 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[5]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_5 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_5 <= remap_table_1_5;
        end
      end else begin
        br_snapshots_6_5 <= _GEN_450;
      end
    end else begin
      br_snapshots_6_5 <= _GEN_450;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_6 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[6]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_6 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_6 <= remap_table_1_6;
        end
      end else begin
        br_snapshots_6_6 <= _GEN_462;
      end
    end else begin
      br_snapshots_6_6 <= _GEN_462;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_7 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[7]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_7 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_7 <= remap_table_1_7;
        end
      end else begin
        br_snapshots_6_7 <= _GEN_474;
      end
    end else begin
      br_snapshots_6_7 <= _GEN_474;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_8 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[8]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_8 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_8 <= remap_table_1_8;
        end
      end else begin
        br_snapshots_6_8 <= _GEN_486;
      end
    end else begin
      br_snapshots_6_8 <= _GEN_486;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_9 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[9]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_9 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_9 <= remap_table_1_9;
        end
      end else begin
        br_snapshots_6_9 <= _GEN_498;
      end
    end else begin
      br_snapshots_6_9 <= _GEN_498;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_10 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[10]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_10 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_10 <= remap_table_1_10;
        end
      end else begin
        br_snapshots_6_10 <= _GEN_510;
      end
    end else begin
      br_snapshots_6_10 <= _GEN_510;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_11 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[11]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_11 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_11 <= remap_table_1_11;
        end
      end else begin
        br_snapshots_6_11 <= _GEN_522;
      end
    end else begin
      br_snapshots_6_11 <= _GEN_522;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_12 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[12]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_12 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_12 <= remap_table_1_12;
        end
      end else begin
        br_snapshots_6_12 <= _GEN_534;
      end
    end else begin
      br_snapshots_6_12 <= _GEN_534;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_13 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[13]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_13 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_13 <= remap_table_1_13;
        end
      end else begin
        br_snapshots_6_13 <= _GEN_546;
      end
    end else begin
      br_snapshots_6_13 <= _GEN_546;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_14 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[14]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_14 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_14 <= remap_table_1_14;
        end
      end else begin
        br_snapshots_6_14 <= _GEN_558;
      end
    end else begin
      br_snapshots_6_14 <= _GEN_558;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_15 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[15]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_15 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_15 <= remap_table_1_15;
        end
      end else begin
        br_snapshots_6_15 <= _GEN_570;
      end
    end else begin
      br_snapshots_6_15 <= _GEN_570;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_16 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[16]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_16 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_16 <= remap_table_1_16;
        end
      end else begin
        br_snapshots_6_16 <= _GEN_582;
      end
    end else begin
      br_snapshots_6_16 <= _GEN_582;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_17 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[17]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_17 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_17 <= remap_table_1_17;
        end
      end else begin
        br_snapshots_6_17 <= _GEN_594;
      end
    end else begin
      br_snapshots_6_17 <= _GEN_594;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_18 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[18]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_18 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_18 <= remap_table_1_18;
        end
      end else begin
        br_snapshots_6_18 <= _GEN_606;
      end
    end else begin
      br_snapshots_6_18 <= _GEN_606;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_19 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[19]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_19 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_19 <= remap_table_1_19;
        end
      end else begin
        br_snapshots_6_19 <= _GEN_618;
      end
    end else begin
      br_snapshots_6_19 <= _GEN_618;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_20 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[20]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_20 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_20 <= remap_table_1_20;
        end
      end else begin
        br_snapshots_6_20 <= _GEN_630;
      end
    end else begin
      br_snapshots_6_20 <= _GEN_630;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_21 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[21]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_21 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_21 <= remap_table_1_21;
        end
      end else begin
        br_snapshots_6_21 <= _GEN_642;
      end
    end else begin
      br_snapshots_6_21 <= _GEN_642;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_22 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[22]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_22 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_22 <= remap_table_1_22;
        end
      end else begin
        br_snapshots_6_22 <= _GEN_654;
      end
    end else begin
      br_snapshots_6_22 <= _GEN_654;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_23 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[23]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_23 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_23 <= remap_table_1_23;
        end
      end else begin
        br_snapshots_6_23 <= _GEN_666;
      end
    end else begin
      br_snapshots_6_23 <= _GEN_666;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_24 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[24]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_24 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_24 <= remap_table_1_24;
        end
      end else begin
        br_snapshots_6_24 <= _GEN_678;
      end
    end else begin
      br_snapshots_6_24 <= _GEN_678;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_25 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[25]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_25 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_25 <= remap_table_1_25;
        end
      end else begin
        br_snapshots_6_25 <= _GEN_690;
      end
    end else begin
      br_snapshots_6_25 <= _GEN_690;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_26 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[26]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_26 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_26 <= remap_table_1_26;
        end
      end else begin
        br_snapshots_6_26 <= _GEN_702;
      end
    end else begin
      br_snapshots_6_26 <= _GEN_702;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_27 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[27]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_27 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_27 <= remap_table_1_27;
        end
      end else begin
        br_snapshots_6_27 <= _GEN_714;
      end
    end else begin
      br_snapshots_6_27 <= _GEN_714;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_28 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[28]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_28 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_28 <= remap_table_1_28;
        end
      end else begin
        br_snapshots_6_28 <= _GEN_726;
      end
    end else begin
      br_snapshots_6_28 <= _GEN_726;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_29 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[29]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_29 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_29 <= remap_table_1_29;
        end
      end else begin
        br_snapshots_6_29 <= _GEN_738;
      end
    end else begin
      br_snapshots_6_29 <= _GEN_738;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_30 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[30]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_30 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_30 <= remap_table_1_30;
        end
      end else begin
        br_snapshots_6_30 <= _GEN_750;
      end
    end else begin
      br_snapshots_6_30 <= _GEN_750;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_6_31 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h6 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[31]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_6_31 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_6_31 <= remap_table_1_31;
        end
      end else begin
        br_snapshots_6_31 <= _GEN_762;
      end
    end else begin
      br_snapshots_6_31 <= _GEN_762;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_1 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[1]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_1 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_1 <= remap_table_1_1;
        end
      end else begin
        br_snapshots_7_1 <= _GEN_403;
      end
    end else begin
      br_snapshots_7_1 <= _GEN_403;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_2 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[2]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_2 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_2 <= remap_table_1_2;
        end
      end else begin
        br_snapshots_7_2 <= _GEN_415;
      end
    end else begin
      br_snapshots_7_2 <= _GEN_415;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_3 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[3]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_3 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_3 <= remap_table_1_3;
        end
      end else begin
        br_snapshots_7_3 <= _GEN_427;
      end
    end else begin
      br_snapshots_7_3 <= _GEN_427;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_4 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[4]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_4 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_4 <= remap_table_1_4;
        end
      end else begin
        br_snapshots_7_4 <= _GEN_439;
      end
    end else begin
      br_snapshots_7_4 <= _GEN_439;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_5 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[5]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_5 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_5 <= remap_table_1_5;
        end
      end else begin
        br_snapshots_7_5 <= _GEN_451;
      end
    end else begin
      br_snapshots_7_5 <= _GEN_451;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_6 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[6]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_6 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_6 <= remap_table_1_6;
        end
      end else begin
        br_snapshots_7_6 <= _GEN_463;
      end
    end else begin
      br_snapshots_7_6 <= _GEN_463;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_7 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[7]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_7 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_7 <= remap_table_1_7;
        end
      end else begin
        br_snapshots_7_7 <= _GEN_475;
      end
    end else begin
      br_snapshots_7_7 <= _GEN_475;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_8 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[8]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_8 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_8 <= remap_table_1_8;
        end
      end else begin
        br_snapshots_7_8 <= _GEN_487;
      end
    end else begin
      br_snapshots_7_8 <= _GEN_487;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_9 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[9]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_9 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_9 <= remap_table_1_9;
        end
      end else begin
        br_snapshots_7_9 <= _GEN_499;
      end
    end else begin
      br_snapshots_7_9 <= _GEN_499;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_10 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[10]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_10 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_10 <= remap_table_1_10;
        end
      end else begin
        br_snapshots_7_10 <= _GEN_511;
      end
    end else begin
      br_snapshots_7_10 <= _GEN_511;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_11 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[11]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_11 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_11 <= remap_table_1_11;
        end
      end else begin
        br_snapshots_7_11 <= _GEN_523;
      end
    end else begin
      br_snapshots_7_11 <= _GEN_523;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_12 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[12]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_12 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_12 <= remap_table_1_12;
        end
      end else begin
        br_snapshots_7_12 <= _GEN_535;
      end
    end else begin
      br_snapshots_7_12 <= _GEN_535;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_13 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[13]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_13 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_13 <= remap_table_1_13;
        end
      end else begin
        br_snapshots_7_13 <= _GEN_547;
      end
    end else begin
      br_snapshots_7_13 <= _GEN_547;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_14 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[14]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_14 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_14 <= remap_table_1_14;
        end
      end else begin
        br_snapshots_7_14 <= _GEN_559;
      end
    end else begin
      br_snapshots_7_14 <= _GEN_559;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_15 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[15]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_15 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_15 <= remap_table_1_15;
        end
      end else begin
        br_snapshots_7_15 <= _GEN_571;
      end
    end else begin
      br_snapshots_7_15 <= _GEN_571;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_16 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[16]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_16 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_16 <= remap_table_1_16;
        end
      end else begin
        br_snapshots_7_16 <= _GEN_583;
      end
    end else begin
      br_snapshots_7_16 <= _GEN_583;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_17 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[17]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_17 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_17 <= remap_table_1_17;
        end
      end else begin
        br_snapshots_7_17 <= _GEN_595;
      end
    end else begin
      br_snapshots_7_17 <= _GEN_595;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_18 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[18]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_18 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_18 <= remap_table_1_18;
        end
      end else begin
        br_snapshots_7_18 <= _GEN_607;
      end
    end else begin
      br_snapshots_7_18 <= _GEN_607;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_19 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[19]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_19 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_19 <= remap_table_1_19;
        end
      end else begin
        br_snapshots_7_19 <= _GEN_619;
      end
    end else begin
      br_snapshots_7_19 <= _GEN_619;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_20 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[20]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_20 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_20 <= remap_table_1_20;
        end
      end else begin
        br_snapshots_7_20 <= _GEN_631;
      end
    end else begin
      br_snapshots_7_20 <= _GEN_631;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_21 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[21]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_21 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_21 <= remap_table_1_21;
        end
      end else begin
        br_snapshots_7_21 <= _GEN_643;
      end
    end else begin
      br_snapshots_7_21 <= _GEN_643;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_22 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[22]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_22 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_22 <= remap_table_1_22;
        end
      end else begin
        br_snapshots_7_22 <= _GEN_655;
      end
    end else begin
      br_snapshots_7_22 <= _GEN_655;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_23 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[23]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_23 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_23 <= remap_table_1_23;
        end
      end else begin
        br_snapshots_7_23 <= _GEN_667;
      end
    end else begin
      br_snapshots_7_23 <= _GEN_667;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_24 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[24]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_24 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_24 <= remap_table_1_24;
        end
      end else begin
        br_snapshots_7_24 <= _GEN_679;
      end
    end else begin
      br_snapshots_7_24 <= _GEN_679;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_25 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[25]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_25 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_25 <= remap_table_1_25;
        end
      end else begin
        br_snapshots_7_25 <= _GEN_691;
      end
    end else begin
      br_snapshots_7_25 <= _GEN_691;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_26 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[26]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_26 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_26 <= remap_table_1_26;
        end
      end else begin
        br_snapshots_7_26 <= _GEN_703;
      end
    end else begin
      br_snapshots_7_26 <= _GEN_703;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_27 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[27]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_27 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_27 <= remap_table_1_27;
        end
      end else begin
        br_snapshots_7_27 <= _GEN_715;
      end
    end else begin
      br_snapshots_7_27 <= _GEN_715;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_28 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[28]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_28 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_28 <= remap_table_1_28;
        end
      end else begin
        br_snapshots_7_28 <= _GEN_727;
      end
    end else begin
      br_snapshots_7_28 <= _GEN_727;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_29 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[29]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_29 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_29 <= remap_table_1_29;
        end
      end else begin
        br_snapshots_7_29 <= _GEN_739;
      end
    end else begin
      br_snapshots_7_29 <= _GEN_739;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_30 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[30]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_30 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_30 <= remap_table_1_30;
        end
      end else begin
        br_snapshots_7_30 <= _GEN_751;
      end
    end else begin
      br_snapshots_7_30 <= _GEN_751;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_7_31 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h7 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[31]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_7_31 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_7_31 <= remap_table_1_31;
        end
      end else begin
        br_snapshots_7_31 <= _GEN_763;
      end
    end else begin
      br_snapshots_7_31 <= _GEN_763;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_1 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[1]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_1 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_1 <= remap_table_1_1;
        end
      end else begin
        br_snapshots_8_1 <= _GEN_404;
      end
    end else begin
      br_snapshots_8_1 <= _GEN_404;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_2 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[2]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_2 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_2 <= remap_table_1_2;
        end
      end else begin
        br_snapshots_8_2 <= _GEN_416;
      end
    end else begin
      br_snapshots_8_2 <= _GEN_416;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_3 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[3]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_3 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_3 <= remap_table_1_3;
        end
      end else begin
        br_snapshots_8_3 <= _GEN_428;
      end
    end else begin
      br_snapshots_8_3 <= _GEN_428;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_4 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[4]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_4 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_4 <= remap_table_1_4;
        end
      end else begin
        br_snapshots_8_4 <= _GEN_440;
      end
    end else begin
      br_snapshots_8_4 <= _GEN_440;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_5 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[5]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_5 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_5 <= remap_table_1_5;
        end
      end else begin
        br_snapshots_8_5 <= _GEN_452;
      end
    end else begin
      br_snapshots_8_5 <= _GEN_452;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_6 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[6]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_6 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_6 <= remap_table_1_6;
        end
      end else begin
        br_snapshots_8_6 <= _GEN_464;
      end
    end else begin
      br_snapshots_8_6 <= _GEN_464;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_7 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[7]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_7 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_7 <= remap_table_1_7;
        end
      end else begin
        br_snapshots_8_7 <= _GEN_476;
      end
    end else begin
      br_snapshots_8_7 <= _GEN_476;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_8 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[8]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_8 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_8 <= remap_table_1_8;
        end
      end else begin
        br_snapshots_8_8 <= _GEN_488;
      end
    end else begin
      br_snapshots_8_8 <= _GEN_488;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_9 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[9]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_9 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_9 <= remap_table_1_9;
        end
      end else begin
        br_snapshots_8_9 <= _GEN_500;
      end
    end else begin
      br_snapshots_8_9 <= _GEN_500;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_10 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[10]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_10 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_10 <= remap_table_1_10;
        end
      end else begin
        br_snapshots_8_10 <= _GEN_512;
      end
    end else begin
      br_snapshots_8_10 <= _GEN_512;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_11 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[11]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_11 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_11 <= remap_table_1_11;
        end
      end else begin
        br_snapshots_8_11 <= _GEN_524;
      end
    end else begin
      br_snapshots_8_11 <= _GEN_524;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_12 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[12]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_12 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_12 <= remap_table_1_12;
        end
      end else begin
        br_snapshots_8_12 <= _GEN_536;
      end
    end else begin
      br_snapshots_8_12 <= _GEN_536;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_13 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[13]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_13 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_13 <= remap_table_1_13;
        end
      end else begin
        br_snapshots_8_13 <= _GEN_548;
      end
    end else begin
      br_snapshots_8_13 <= _GEN_548;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_14 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[14]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_14 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_14 <= remap_table_1_14;
        end
      end else begin
        br_snapshots_8_14 <= _GEN_560;
      end
    end else begin
      br_snapshots_8_14 <= _GEN_560;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_15 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[15]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_15 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_15 <= remap_table_1_15;
        end
      end else begin
        br_snapshots_8_15 <= _GEN_572;
      end
    end else begin
      br_snapshots_8_15 <= _GEN_572;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_16 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[16]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_16 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_16 <= remap_table_1_16;
        end
      end else begin
        br_snapshots_8_16 <= _GEN_584;
      end
    end else begin
      br_snapshots_8_16 <= _GEN_584;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_17 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[17]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_17 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_17 <= remap_table_1_17;
        end
      end else begin
        br_snapshots_8_17 <= _GEN_596;
      end
    end else begin
      br_snapshots_8_17 <= _GEN_596;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_18 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[18]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_18 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_18 <= remap_table_1_18;
        end
      end else begin
        br_snapshots_8_18 <= _GEN_608;
      end
    end else begin
      br_snapshots_8_18 <= _GEN_608;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_19 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[19]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_19 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_19 <= remap_table_1_19;
        end
      end else begin
        br_snapshots_8_19 <= _GEN_620;
      end
    end else begin
      br_snapshots_8_19 <= _GEN_620;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_20 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[20]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_20 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_20 <= remap_table_1_20;
        end
      end else begin
        br_snapshots_8_20 <= _GEN_632;
      end
    end else begin
      br_snapshots_8_20 <= _GEN_632;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_21 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[21]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_21 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_21 <= remap_table_1_21;
        end
      end else begin
        br_snapshots_8_21 <= _GEN_644;
      end
    end else begin
      br_snapshots_8_21 <= _GEN_644;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_22 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[22]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_22 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_22 <= remap_table_1_22;
        end
      end else begin
        br_snapshots_8_22 <= _GEN_656;
      end
    end else begin
      br_snapshots_8_22 <= _GEN_656;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_23 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[23]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_23 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_23 <= remap_table_1_23;
        end
      end else begin
        br_snapshots_8_23 <= _GEN_668;
      end
    end else begin
      br_snapshots_8_23 <= _GEN_668;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_24 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[24]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_24 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_24 <= remap_table_1_24;
        end
      end else begin
        br_snapshots_8_24 <= _GEN_680;
      end
    end else begin
      br_snapshots_8_24 <= _GEN_680;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_25 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[25]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_25 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_25 <= remap_table_1_25;
        end
      end else begin
        br_snapshots_8_25 <= _GEN_692;
      end
    end else begin
      br_snapshots_8_25 <= _GEN_692;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_26 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[26]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_26 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_26 <= remap_table_1_26;
        end
      end else begin
        br_snapshots_8_26 <= _GEN_704;
      end
    end else begin
      br_snapshots_8_26 <= _GEN_704;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_27 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[27]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_27 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_27 <= remap_table_1_27;
        end
      end else begin
        br_snapshots_8_27 <= _GEN_716;
      end
    end else begin
      br_snapshots_8_27 <= _GEN_716;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_28 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[28]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_28 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_28 <= remap_table_1_28;
        end
      end else begin
        br_snapshots_8_28 <= _GEN_728;
      end
    end else begin
      br_snapshots_8_28 <= _GEN_728;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_29 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[29]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_29 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_29 <= remap_table_1_29;
        end
      end else begin
        br_snapshots_8_29 <= _GEN_740;
      end
    end else begin
      br_snapshots_8_29 <= _GEN_740;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_30 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[30]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_30 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_30 <= remap_table_1_30;
        end
      end else begin
        br_snapshots_8_30 <= _GEN_752;
      end
    end else begin
      br_snapshots_8_30 <= _GEN_752;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_8_31 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h8 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[31]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_8_31 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_8_31 <= remap_table_1_31;
        end
      end else begin
        br_snapshots_8_31 <= _GEN_764;
      end
    end else begin
      br_snapshots_8_31 <= _GEN_764;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_1 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[1]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_1 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_1 <= remap_table_1_1;
        end
      end else begin
        br_snapshots_9_1 <= _GEN_405;
      end
    end else begin
      br_snapshots_9_1 <= _GEN_405;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_2 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[2]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_2 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_2 <= remap_table_1_2;
        end
      end else begin
        br_snapshots_9_2 <= _GEN_417;
      end
    end else begin
      br_snapshots_9_2 <= _GEN_417;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_3 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[3]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_3 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_3 <= remap_table_1_3;
        end
      end else begin
        br_snapshots_9_3 <= _GEN_429;
      end
    end else begin
      br_snapshots_9_3 <= _GEN_429;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_4 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[4]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_4 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_4 <= remap_table_1_4;
        end
      end else begin
        br_snapshots_9_4 <= _GEN_441;
      end
    end else begin
      br_snapshots_9_4 <= _GEN_441;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_5 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[5]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_5 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_5 <= remap_table_1_5;
        end
      end else begin
        br_snapshots_9_5 <= _GEN_453;
      end
    end else begin
      br_snapshots_9_5 <= _GEN_453;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_6 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[6]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_6 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_6 <= remap_table_1_6;
        end
      end else begin
        br_snapshots_9_6 <= _GEN_465;
      end
    end else begin
      br_snapshots_9_6 <= _GEN_465;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_7 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[7]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_7 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_7 <= remap_table_1_7;
        end
      end else begin
        br_snapshots_9_7 <= _GEN_477;
      end
    end else begin
      br_snapshots_9_7 <= _GEN_477;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_8 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[8]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_8 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_8 <= remap_table_1_8;
        end
      end else begin
        br_snapshots_9_8 <= _GEN_489;
      end
    end else begin
      br_snapshots_9_8 <= _GEN_489;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_9 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[9]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_9 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_9 <= remap_table_1_9;
        end
      end else begin
        br_snapshots_9_9 <= _GEN_501;
      end
    end else begin
      br_snapshots_9_9 <= _GEN_501;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_10 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[10]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_10 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_10 <= remap_table_1_10;
        end
      end else begin
        br_snapshots_9_10 <= _GEN_513;
      end
    end else begin
      br_snapshots_9_10 <= _GEN_513;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_11 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[11]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_11 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_11 <= remap_table_1_11;
        end
      end else begin
        br_snapshots_9_11 <= _GEN_525;
      end
    end else begin
      br_snapshots_9_11 <= _GEN_525;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_12 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[12]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_12 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_12 <= remap_table_1_12;
        end
      end else begin
        br_snapshots_9_12 <= _GEN_537;
      end
    end else begin
      br_snapshots_9_12 <= _GEN_537;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_13 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[13]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_13 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_13 <= remap_table_1_13;
        end
      end else begin
        br_snapshots_9_13 <= _GEN_549;
      end
    end else begin
      br_snapshots_9_13 <= _GEN_549;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_14 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[14]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_14 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_14 <= remap_table_1_14;
        end
      end else begin
        br_snapshots_9_14 <= _GEN_561;
      end
    end else begin
      br_snapshots_9_14 <= _GEN_561;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_15 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[15]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_15 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_15 <= remap_table_1_15;
        end
      end else begin
        br_snapshots_9_15 <= _GEN_573;
      end
    end else begin
      br_snapshots_9_15 <= _GEN_573;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_16 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[16]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_16 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_16 <= remap_table_1_16;
        end
      end else begin
        br_snapshots_9_16 <= _GEN_585;
      end
    end else begin
      br_snapshots_9_16 <= _GEN_585;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_17 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[17]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_17 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_17 <= remap_table_1_17;
        end
      end else begin
        br_snapshots_9_17 <= _GEN_597;
      end
    end else begin
      br_snapshots_9_17 <= _GEN_597;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_18 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[18]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_18 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_18 <= remap_table_1_18;
        end
      end else begin
        br_snapshots_9_18 <= _GEN_609;
      end
    end else begin
      br_snapshots_9_18 <= _GEN_609;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_19 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[19]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_19 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_19 <= remap_table_1_19;
        end
      end else begin
        br_snapshots_9_19 <= _GEN_621;
      end
    end else begin
      br_snapshots_9_19 <= _GEN_621;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_20 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[20]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_20 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_20 <= remap_table_1_20;
        end
      end else begin
        br_snapshots_9_20 <= _GEN_633;
      end
    end else begin
      br_snapshots_9_20 <= _GEN_633;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_21 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[21]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_21 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_21 <= remap_table_1_21;
        end
      end else begin
        br_snapshots_9_21 <= _GEN_645;
      end
    end else begin
      br_snapshots_9_21 <= _GEN_645;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_22 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[22]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_22 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_22 <= remap_table_1_22;
        end
      end else begin
        br_snapshots_9_22 <= _GEN_657;
      end
    end else begin
      br_snapshots_9_22 <= _GEN_657;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_23 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[23]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_23 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_23 <= remap_table_1_23;
        end
      end else begin
        br_snapshots_9_23 <= _GEN_669;
      end
    end else begin
      br_snapshots_9_23 <= _GEN_669;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_24 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[24]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_24 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_24 <= remap_table_1_24;
        end
      end else begin
        br_snapshots_9_24 <= _GEN_681;
      end
    end else begin
      br_snapshots_9_24 <= _GEN_681;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_25 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[25]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_25 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_25 <= remap_table_1_25;
        end
      end else begin
        br_snapshots_9_25 <= _GEN_693;
      end
    end else begin
      br_snapshots_9_25 <= _GEN_693;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_26 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[26]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_26 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_26 <= remap_table_1_26;
        end
      end else begin
        br_snapshots_9_26 <= _GEN_705;
      end
    end else begin
      br_snapshots_9_26 <= _GEN_705;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_27 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[27]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_27 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_27 <= remap_table_1_27;
        end
      end else begin
        br_snapshots_9_27 <= _GEN_717;
      end
    end else begin
      br_snapshots_9_27 <= _GEN_717;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_28 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[28]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_28 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_28 <= remap_table_1_28;
        end
      end else begin
        br_snapshots_9_28 <= _GEN_729;
      end
    end else begin
      br_snapshots_9_28 <= _GEN_729;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_29 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[29]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_29 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_29 <= remap_table_1_29;
        end
      end else begin
        br_snapshots_9_29 <= _GEN_741;
      end
    end else begin
      br_snapshots_9_29 <= _GEN_741;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_30 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[30]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_30 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_30 <= remap_table_1_30;
        end
      end else begin
        br_snapshots_9_30 <= _GEN_753;
      end
    end else begin
      br_snapshots_9_30 <= _GEN_753;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_9_31 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'h9 == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[31]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_9_31 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_9_31 <= remap_table_1_31;
        end
      end else begin
        br_snapshots_9_31 <= _GEN_765;
      end
    end else begin
      br_snapshots_9_31 <= _GEN_765;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_1 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[1]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_1 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_1 <= remap_table_1_1;
        end
      end else begin
        br_snapshots_10_1 <= _GEN_406;
      end
    end else begin
      br_snapshots_10_1 <= _GEN_406;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_2 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[2]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_2 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_2 <= remap_table_1_2;
        end
      end else begin
        br_snapshots_10_2 <= _GEN_418;
      end
    end else begin
      br_snapshots_10_2 <= _GEN_418;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_3 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[3]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_3 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_3 <= remap_table_1_3;
        end
      end else begin
        br_snapshots_10_3 <= _GEN_430;
      end
    end else begin
      br_snapshots_10_3 <= _GEN_430;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_4 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[4]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_4 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_4 <= remap_table_1_4;
        end
      end else begin
        br_snapshots_10_4 <= _GEN_442;
      end
    end else begin
      br_snapshots_10_4 <= _GEN_442;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_5 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[5]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_5 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_5 <= remap_table_1_5;
        end
      end else begin
        br_snapshots_10_5 <= _GEN_454;
      end
    end else begin
      br_snapshots_10_5 <= _GEN_454;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_6 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[6]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_6 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_6 <= remap_table_1_6;
        end
      end else begin
        br_snapshots_10_6 <= _GEN_466;
      end
    end else begin
      br_snapshots_10_6 <= _GEN_466;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_7 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[7]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_7 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_7 <= remap_table_1_7;
        end
      end else begin
        br_snapshots_10_7 <= _GEN_478;
      end
    end else begin
      br_snapshots_10_7 <= _GEN_478;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_8 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[8]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_8 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_8 <= remap_table_1_8;
        end
      end else begin
        br_snapshots_10_8 <= _GEN_490;
      end
    end else begin
      br_snapshots_10_8 <= _GEN_490;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_9 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[9]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_9 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_9 <= remap_table_1_9;
        end
      end else begin
        br_snapshots_10_9 <= _GEN_502;
      end
    end else begin
      br_snapshots_10_9 <= _GEN_502;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_10 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[10]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_10 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_10 <= remap_table_1_10;
        end
      end else begin
        br_snapshots_10_10 <= _GEN_514;
      end
    end else begin
      br_snapshots_10_10 <= _GEN_514;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_11 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[11]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_11 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_11 <= remap_table_1_11;
        end
      end else begin
        br_snapshots_10_11 <= _GEN_526;
      end
    end else begin
      br_snapshots_10_11 <= _GEN_526;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_12 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[12]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_12 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_12 <= remap_table_1_12;
        end
      end else begin
        br_snapshots_10_12 <= _GEN_538;
      end
    end else begin
      br_snapshots_10_12 <= _GEN_538;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_13 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[13]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_13 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_13 <= remap_table_1_13;
        end
      end else begin
        br_snapshots_10_13 <= _GEN_550;
      end
    end else begin
      br_snapshots_10_13 <= _GEN_550;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_14 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[14]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_14 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_14 <= remap_table_1_14;
        end
      end else begin
        br_snapshots_10_14 <= _GEN_562;
      end
    end else begin
      br_snapshots_10_14 <= _GEN_562;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_15 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[15]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_15 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_15 <= remap_table_1_15;
        end
      end else begin
        br_snapshots_10_15 <= _GEN_574;
      end
    end else begin
      br_snapshots_10_15 <= _GEN_574;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_16 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[16]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_16 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_16 <= remap_table_1_16;
        end
      end else begin
        br_snapshots_10_16 <= _GEN_586;
      end
    end else begin
      br_snapshots_10_16 <= _GEN_586;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_17 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[17]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_17 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_17 <= remap_table_1_17;
        end
      end else begin
        br_snapshots_10_17 <= _GEN_598;
      end
    end else begin
      br_snapshots_10_17 <= _GEN_598;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_18 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[18]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_18 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_18 <= remap_table_1_18;
        end
      end else begin
        br_snapshots_10_18 <= _GEN_610;
      end
    end else begin
      br_snapshots_10_18 <= _GEN_610;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_19 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[19]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_19 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_19 <= remap_table_1_19;
        end
      end else begin
        br_snapshots_10_19 <= _GEN_622;
      end
    end else begin
      br_snapshots_10_19 <= _GEN_622;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_20 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[20]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_20 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_20 <= remap_table_1_20;
        end
      end else begin
        br_snapshots_10_20 <= _GEN_634;
      end
    end else begin
      br_snapshots_10_20 <= _GEN_634;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_21 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[21]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_21 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_21 <= remap_table_1_21;
        end
      end else begin
        br_snapshots_10_21 <= _GEN_646;
      end
    end else begin
      br_snapshots_10_21 <= _GEN_646;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_22 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[22]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_22 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_22 <= remap_table_1_22;
        end
      end else begin
        br_snapshots_10_22 <= _GEN_658;
      end
    end else begin
      br_snapshots_10_22 <= _GEN_658;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_23 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[23]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_23 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_23 <= remap_table_1_23;
        end
      end else begin
        br_snapshots_10_23 <= _GEN_670;
      end
    end else begin
      br_snapshots_10_23 <= _GEN_670;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_24 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[24]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_24 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_24 <= remap_table_1_24;
        end
      end else begin
        br_snapshots_10_24 <= _GEN_682;
      end
    end else begin
      br_snapshots_10_24 <= _GEN_682;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_25 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[25]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_25 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_25 <= remap_table_1_25;
        end
      end else begin
        br_snapshots_10_25 <= _GEN_694;
      end
    end else begin
      br_snapshots_10_25 <= _GEN_694;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_26 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[26]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_26 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_26 <= remap_table_1_26;
        end
      end else begin
        br_snapshots_10_26 <= _GEN_706;
      end
    end else begin
      br_snapshots_10_26 <= _GEN_706;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_27 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[27]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_27 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_27 <= remap_table_1_27;
        end
      end else begin
        br_snapshots_10_27 <= _GEN_718;
      end
    end else begin
      br_snapshots_10_27 <= _GEN_718;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_28 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[28]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_28 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_28 <= remap_table_1_28;
        end
      end else begin
        br_snapshots_10_28 <= _GEN_730;
      end
    end else begin
      br_snapshots_10_28 <= _GEN_730;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_29 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[29]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_29 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_29 <= remap_table_1_29;
        end
      end else begin
        br_snapshots_10_29 <= _GEN_742;
      end
    end else begin
      br_snapshots_10_29 <= _GEN_742;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_30 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[30]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_30 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_30 <= remap_table_1_30;
        end
      end else begin
        br_snapshots_10_30 <= _GEN_754;
      end
    end else begin
      br_snapshots_10_30 <= _GEN_754;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_10_31 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'ha == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[31]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_10_31 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_10_31 <= remap_table_1_31;
        end
      end else begin
        br_snapshots_10_31 <= _GEN_766;
      end
    end else begin
      br_snapshots_10_31 <= _GEN_766;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_1 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[1]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_1 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_1 <= remap_table_1_1;
        end
      end else begin
        br_snapshots_11_1 <= _GEN_407;
      end
    end else begin
      br_snapshots_11_1 <= _GEN_407;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_2 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[2]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_2 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_2 <= remap_table_1_2;
        end
      end else begin
        br_snapshots_11_2 <= _GEN_419;
      end
    end else begin
      br_snapshots_11_2 <= _GEN_419;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_3 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[3]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_3 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_3 <= remap_table_1_3;
        end
      end else begin
        br_snapshots_11_3 <= _GEN_431;
      end
    end else begin
      br_snapshots_11_3 <= _GEN_431;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_4 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[4]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_4 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_4 <= remap_table_1_4;
        end
      end else begin
        br_snapshots_11_4 <= _GEN_443;
      end
    end else begin
      br_snapshots_11_4 <= _GEN_443;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_5 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[5]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_5 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_5 <= remap_table_1_5;
        end
      end else begin
        br_snapshots_11_5 <= _GEN_455;
      end
    end else begin
      br_snapshots_11_5 <= _GEN_455;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_6 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[6]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_6 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_6 <= remap_table_1_6;
        end
      end else begin
        br_snapshots_11_6 <= _GEN_467;
      end
    end else begin
      br_snapshots_11_6 <= _GEN_467;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_7 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[7]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_7 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_7 <= remap_table_1_7;
        end
      end else begin
        br_snapshots_11_7 <= _GEN_479;
      end
    end else begin
      br_snapshots_11_7 <= _GEN_479;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_8 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[8]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_8 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_8 <= remap_table_1_8;
        end
      end else begin
        br_snapshots_11_8 <= _GEN_491;
      end
    end else begin
      br_snapshots_11_8 <= _GEN_491;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_9 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[9]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_9 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_9 <= remap_table_1_9;
        end
      end else begin
        br_snapshots_11_9 <= _GEN_503;
      end
    end else begin
      br_snapshots_11_9 <= _GEN_503;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_10 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[10]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_10 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_10 <= remap_table_1_10;
        end
      end else begin
        br_snapshots_11_10 <= _GEN_515;
      end
    end else begin
      br_snapshots_11_10 <= _GEN_515;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_11 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[11]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_11 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_11 <= remap_table_1_11;
        end
      end else begin
        br_snapshots_11_11 <= _GEN_527;
      end
    end else begin
      br_snapshots_11_11 <= _GEN_527;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_12 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[12]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_12 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_12 <= remap_table_1_12;
        end
      end else begin
        br_snapshots_11_12 <= _GEN_539;
      end
    end else begin
      br_snapshots_11_12 <= _GEN_539;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_13 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[13]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_13 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_13 <= remap_table_1_13;
        end
      end else begin
        br_snapshots_11_13 <= _GEN_551;
      end
    end else begin
      br_snapshots_11_13 <= _GEN_551;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_14 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[14]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_14 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_14 <= remap_table_1_14;
        end
      end else begin
        br_snapshots_11_14 <= _GEN_563;
      end
    end else begin
      br_snapshots_11_14 <= _GEN_563;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_15 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[15]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_15 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_15 <= remap_table_1_15;
        end
      end else begin
        br_snapshots_11_15 <= _GEN_575;
      end
    end else begin
      br_snapshots_11_15 <= _GEN_575;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_16 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[16]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_16 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_16 <= remap_table_1_16;
        end
      end else begin
        br_snapshots_11_16 <= _GEN_587;
      end
    end else begin
      br_snapshots_11_16 <= _GEN_587;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_17 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[17]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_17 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_17 <= remap_table_1_17;
        end
      end else begin
        br_snapshots_11_17 <= _GEN_599;
      end
    end else begin
      br_snapshots_11_17 <= _GEN_599;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_18 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[18]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_18 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_18 <= remap_table_1_18;
        end
      end else begin
        br_snapshots_11_18 <= _GEN_611;
      end
    end else begin
      br_snapshots_11_18 <= _GEN_611;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_19 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[19]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_19 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_19 <= remap_table_1_19;
        end
      end else begin
        br_snapshots_11_19 <= _GEN_623;
      end
    end else begin
      br_snapshots_11_19 <= _GEN_623;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_20 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[20]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_20 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_20 <= remap_table_1_20;
        end
      end else begin
        br_snapshots_11_20 <= _GEN_635;
      end
    end else begin
      br_snapshots_11_20 <= _GEN_635;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_21 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[21]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_21 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_21 <= remap_table_1_21;
        end
      end else begin
        br_snapshots_11_21 <= _GEN_647;
      end
    end else begin
      br_snapshots_11_21 <= _GEN_647;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_22 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[22]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_22 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_22 <= remap_table_1_22;
        end
      end else begin
        br_snapshots_11_22 <= _GEN_659;
      end
    end else begin
      br_snapshots_11_22 <= _GEN_659;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_23 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[23]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_23 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_23 <= remap_table_1_23;
        end
      end else begin
        br_snapshots_11_23 <= _GEN_671;
      end
    end else begin
      br_snapshots_11_23 <= _GEN_671;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_24 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[24]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_24 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_24 <= remap_table_1_24;
        end
      end else begin
        br_snapshots_11_24 <= _GEN_683;
      end
    end else begin
      br_snapshots_11_24 <= _GEN_683;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_25 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[25]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_25 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_25 <= remap_table_1_25;
        end
      end else begin
        br_snapshots_11_25 <= _GEN_695;
      end
    end else begin
      br_snapshots_11_25 <= _GEN_695;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_26 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[26]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_26 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_26 <= remap_table_1_26;
        end
      end else begin
        br_snapshots_11_26 <= _GEN_707;
      end
    end else begin
      br_snapshots_11_26 <= _GEN_707;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_27 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[27]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_27 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_27 <= remap_table_1_27;
        end
      end else begin
        br_snapshots_11_27 <= _GEN_719;
      end
    end else begin
      br_snapshots_11_27 <= _GEN_719;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_28 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[28]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_28 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_28 <= remap_table_1_28;
        end
      end else begin
        br_snapshots_11_28 <= _GEN_731;
      end
    end else begin
      br_snapshots_11_28 <= _GEN_731;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_29 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[29]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_29 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_29 <= remap_table_1_29;
        end
      end else begin
        br_snapshots_11_29 <= _GEN_743;
      end
    end else begin
      br_snapshots_11_29 <= _GEN_743;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_30 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[30]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_30 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_30 <= remap_table_1_30;
        end
      end else begin
        br_snapshots_11_30 <= _GEN_755;
      end
    end else begin
      br_snapshots_11_30 <= _GEN_755;
    end
    if (io_flush) begin // @[rename-maptable.scala 137:19]
      br_snapshots_11_31 <= 6'h0; // @[rename-maptable.scala 143:28]
    end else if (io_ren_br_tags_1_valid) begin // @[rename-maptable.scala 132:36]
      if (4'hb == io_ren_br_tags_1_bits) begin // @[rename-maptable.scala 133:44]
        if (remap_ldsts_oh_1[31]) begin // @[rename-maptable.scala 122:70]
          br_snapshots_11_31 <= io_remap_reqs_1_pdst;
        end else begin
          br_snapshots_11_31 <= remap_table_1_31;
        end
      end else begin
        br_snapshots_11_31 <= _GEN_767;
      end
    end else begin
      br_snapshots_11_31 <= _GEN_767;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~io_remap_reqs_0_valid | ~(_T_612 | map_table_31 == io_remap_reqs_0_pdst) | io_remap_reqs_0_pdst == 6'h0
           & io_rollback | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [maptable] Trying to write a duplicate mapping.\n    at rename-maptable.scala:176 assert (!r || !map_table.contains(p) || p === 0.U && io.rollback, \"[maptable] Trying to write a duplicate mapping.\")}\n"
            ); // @[rename-maptable.scala 176:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~io_remap_reqs_0_valid | ~(_T_612 | map_table_31 == io_remap_reqs_0_pdst) | io_remap_reqs_0_pdst == 6'h0
           & io_rollback | reset)) begin
          $fatal; // @[rename-maptable.scala 176:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~io_remap_reqs_1_valid | ~(_T_685 | map_table_31 == io_remap_reqs_1_pdst) | io_remap_reqs_1_pdst == 6'h0
           & io_rollback | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [maptable] Trying to write a duplicate mapping.\n    at rename-maptable.scala:176 assert (!r || !map_table.contains(p) || p === 0.U && io.rollback, \"[maptable] Trying to write a duplicate mapping.\")}\n"
            ); // @[rename-maptable.scala 176:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~io_remap_reqs_1_valid | ~(_T_685 | map_table_31 == io_remap_reqs_1_pdst) | io_remap_reqs_1_pdst == 6'h0
           & io_rollback | reset)) begin
          $fatal; // @[rename-maptable.scala 176:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  map_table_0 = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  map_table_1 = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  map_table_2 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  map_table_3 = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  map_table_4 = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  map_table_5 = _RAND_5[5:0];
  _RAND_6 = {1{`RANDOM}};
  map_table_6 = _RAND_6[5:0];
  _RAND_7 = {1{`RANDOM}};
  map_table_7 = _RAND_7[5:0];
  _RAND_8 = {1{`RANDOM}};
  map_table_8 = _RAND_8[5:0];
  _RAND_9 = {1{`RANDOM}};
  map_table_9 = _RAND_9[5:0];
  _RAND_10 = {1{`RANDOM}};
  map_table_10 = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  map_table_11 = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  map_table_12 = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  map_table_13 = _RAND_13[5:0];
  _RAND_14 = {1{`RANDOM}};
  map_table_14 = _RAND_14[5:0];
  _RAND_15 = {1{`RANDOM}};
  map_table_15 = _RAND_15[5:0];
  _RAND_16 = {1{`RANDOM}};
  map_table_16 = _RAND_16[5:0];
  _RAND_17 = {1{`RANDOM}};
  map_table_17 = _RAND_17[5:0];
  _RAND_18 = {1{`RANDOM}};
  map_table_18 = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
  map_table_19 = _RAND_19[5:0];
  _RAND_20 = {1{`RANDOM}};
  map_table_20 = _RAND_20[5:0];
  _RAND_21 = {1{`RANDOM}};
  map_table_21 = _RAND_21[5:0];
  _RAND_22 = {1{`RANDOM}};
  map_table_22 = _RAND_22[5:0];
  _RAND_23 = {1{`RANDOM}};
  map_table_23 = _RAND_23[5:0];
  _RAND_24 = {1{`RANDOM}};
  map_table_24 = _RAND_24[5:0];
  _RAND_25 = {1{`RANDOM}};
  map_table_25 = _RAND_25[5:0];
  _RAND_26 = {1{`RANDOM}};
  map_table_26 = _RAND_26[5:0];
  _RAND_27 = {1{`RANDOM}};
  map_table_27 = _RAND_27[5:0];
  _RAND_28 = {1{`RANDOM}};
  map_table_28 = _RAND_28[5:0];
  _RAND_29 = {1{`RANDOM}};
  map_table_29 = _RAND_29[5:0];
  _RAND_30 = {1{`RANDOM}};
  map_table_30 = _RAND_30[5:0];
  _RAND_31 = {1{`RANDOM}};
  map_table_31 = _RAND_31[5:0];
  _RAND_32 = {1{`RANDOM}};
  commit_map_table_0 = _RAND_32[5:0];
  _RAND_33 = {1{`RANDOM}};
  commit_map_table_1 = _RAND_33[5:0];
  _RAND_34 = {1{`RANDOM}};
  commit_map_table_2 = _RAND_34[5:0];
  _RAND_35 = {1{`RANDOM}};
  commit_map_table_3 = _RAND_35[5:0];
  _RAND_36 = {1{`RANDOM}};
  commit_map_table_4 = _RAND_36[5:0];
  _RAND_37 = {1{`RANDOM}};
  commit_map_table_5 = _RAND_37[5:0];
  _RAND_38 = {1{`RANDOM}};
  commit_map_table_6 = _RAND_38[5:0];
  _RAND_39 = {1{`RANDOM}};
  commit_map_table_7 = _RAND_39[5:0];
  _RAND_40 = {1{`RANDOM}};
  commit_map_table_8 = _RAND_40[5:0];
  _RAND_41 = {1{`RANDOM}};
  commit_map_table_9 = _RAND_41[5:0];
  _RAND_42 = {1{`RANDOM}};
  commit_map_table_10 = _RAND_42[5:0];
  _RAND_43 = {1{`RANDOM}};
  commit_map_table_11 = _RAND_43[5:0];
  _RAND_44 = {1{`RANDOM}};
  commit_map_table_12 = _RAND_44[5:0];
  _RAND_45 = {1{`RANDOM}};
  commit_map_table_13 = _RAND_45[5:0];
  _RAND_46 = {1{`RANDOM}};
  commit_map_table_14 = _RAND_46[5:0];
  _RAND_47 = {1{`RANDOM}};
  commit_map_table_15 = _RAND_47[5:0];
  _RAND_48 = {1{`RANDOM}};
  commit_map_table_16 = _RAND_48[5:0];
  _RAND_49 = {1{`RANDOM}};
  commit_map_table_17 = _RAND_49[5:0];
  _RAND_50 = {1{`RANDOM}};
  commit_map_table_18 = _RAND_50[5:0];
  _RAND_51 = {1{`RANDOM}};
  commit_map_table_19 = _RAND_51[5:0];
  _RAND_52 = {1{`RANDOM}};
  commit_map_table_20 = _RAND_52[5:0];
  _RAND_53 = {1{`RANDOM}};
  commit_map_table_21 = _RAND_53[5:0];
  _RAND_54 = {1{`RANDOM}};
  commit_map_table_22 = _RAND_54[5:0];
  _RAND_55 = {1{`RANDOM}};
  commit_map_table_23 = _RAND_55[5:0];
  _RAND_56 = {1{`RANDOM}};
  commit_map_table_24 = _RAND_56[5:0];
  _RAND_57 = {1{`RANDOM}};
  commit_map_table_25 = _RAND_57[5:0];
  _RAND_58 = {1{`RANDOM}};
  commit_map_table_26 = _RAND_58[5:0];
  _RAND_59 = {1{`RANDOM}};
  commit_map_table_27 = _RAND_59[5:0];
  _RAND_60 = {1{`RANDOM}};
  commit_map_table_28 = _RAND_60[5:0];
  _RAND_61 = {1{`RANDOM}};
  commit_map_table_29 = _RAND_61[5:0];
  _RAND_62 = {1{`RANDOM}};
  commit_map_table_30 = _RAND_62[5:0];
  _RAND_63 = {1{`RANDOM}};
  commit_map_table_31 = _RAND_63[5:0];
  _RAND_64 = {1{`RANDOM}};
  br_snapshots_0_1 = _RAND_64[5:0];
  _RAND_65 = {1{`RANDOM}};
  br_snapshots_0_2 = _RAND_65[5:0];
  _RAND_66 = {1{`RANDOM}};
  br_snapshots_0_3 = _RAND_66[5:0];
  _RAND_67 = {1{`RANDOM}};
  br_snapshots_0_4 = _RAND_67[5:0];
  _RAND_68 = {1{`RANDOM}};
  br_snapshots_0_5 = _RAND_68[5:0];
  _RAND_69 = {1{`RANDOM}};
  br_snapshots_0_6 = _RAND_69[5:0];
  _RAND_70 = {1{`RANDOM}};
  br_snapshots_0_7 = _RAND_70[5:0];
  _RAND_71 = {1{`RANDOM}};
  br_snapshots_0_8 = _RAND_71[5:0];
  _RAND_72 = {1{`RANDOM}};
  br_snapshots_0_9 = _RAND_72[5:0];
  _RAND_73 = {1{`RANDOM}};
  br_snapshots_0_10 = _RAND_73[5:0];
  _RAND_74 = {1{`RANDOM}};
  br_snapshots_0_11 = _RAND_74[5:0];
  _RAND_75 = {1{`RANDOM}};
  br_snapshots_0_12 = _RAND_75[5:0];
  _RAND_76 = {1{`RANDOM}};
  br_snapshots_0_13 = _RAND_76[5:0];
  _RAND_77 = {1{`RANDOM}};
  br_snapshots_0_14 = _RAND_77[5:0];
  _RAND_78 = {1{`RANDOM}};
  br_snapshots_0_15 = _RAND_78[5:0];
  _RAND_79 = {1{`RANDOM}};
  br_snapshots_0_16 = _RAND_79[5:0];
  _RAND_80 = {1{`RANDOM}};
  br_snapshots_0_17 = _RAND_80[5:0];
  _RAND_81 = {1{`RANDOM}};
  br_snapshots_0_18 = _RAND_81[5:0];
  _RAND_82 = {1{`RANDOM}};
  br_snapshots_0_19 = _RAND_82[5:0];
  _RAND_83 = {1{`RANDOM}};
  br_snapshots_0_20 = _RAND_83[5:0];
  _RAND_84 = {1{`RANDOM}};
  br_snapshots_0_21 = _RAND_84[5:0];
  _RAND_85 = {1{`RANDOM}};
  br_snapshots_0_22 = _RAND_85[5:0];
  _RAND_86 = {1{`RANDOM}};
  br_snapshots_0_23 = _RAND_86[5:0];
  _RAND_87 = {1{`RANDOM}};
  br_snapshots_0_24 = _RAND_87[5:0];
  _RAND_88 = {1{`RANDOM}};
  br_snapshots_0_25 = _RAND_88[5:0];
  _RAND_89 = {1{`RANDOM}};
  br_snapshots_0_26 = _RAND_89[5:0];
  _RAND_90 = {1{`RANDOM}};
  br_snapshots_0_27 = _RAND_90[5:0];
  _RAND_91 = {1{`RANDOM}};
  br_snapshots_0_28 = _RAND_91[5:0];
  _RAND_92 = {1{`RANDOM}};
  br_snapshots_0_29 = _RAND_92[5:0];
  _RAND_93 = {1{`RANDOM}};
  br_snapshots_0_30 = _RAND_93[5:0];
  _RAND_94 = {1{`RANDOM}};
  br_snapshots_0_31 = _RAND_94[5:0];
  _RAND_95 = {1{`RANDOM}};
  br_snapshots_1_1 = _RAND_95[5:0];
  _RAND_96 = {1{`RANDOM}};
  br_snapshots_1_2 = _RAND_96[5:0];
  _RAND_97 = {1{`RANDOM}};
  br_snapshots_1_3 = _RAND_97[5:0];
  _RAND_98 = {1{`RANDOM}};
  br_snapshots_1_4 = _RAND_98[5:0];
  _RAND_99 = {1{`RANDOM}};
  br_snapshots_1_5 = _RAND_99[5:0];
  _RAND_100 = {1{`RANDOM}};
  br_snapshots_1_6 = _RAND_100[5:0];
  _RAND_101 = {1{`RANDOM}};
  br_snapshots_1_7 = _RAND_101[5:0];
  _RAND_102 = {1{`RANDOM}};
  br_snapshots_1_8 = _RAND_102[5:0];
  _RAND_103 = {1{`RANDOM}};
  br_snapshots_1_9 = _RAND_103[5:0];
  _RAND_104 = {1{`RANDOM}};
  br_snapshots_1_10 = _RAND_104[5:0];
  _RAND_105 = {1{`RANDOM}};
  br_snapshots_1_11 = _RAND_105[5:0];
  _RAND_106 = {1{`RANDOM}};
  br_snapshots_1_12 = _RAND_106[5:0];
  _RAND_107 = {1{`RANDOM}};
  br_snapshots_1_13 = _RAND_107[5:0];
  _RAND_108 = {1{`RANDOM}};
  br_snapshots_1_14 = _RAND_108[5:0];
  _RAND_109 = {1{`RANDOM}};
  br_snapshots_1_15 = _RAND_109[5:0];
  _RAND_110 = {1{`RANDOM}};
  br_snapshots_1_16 = _RAND_110[5:0];
  _RAND_111 = {1{`RANDOM}};
  br_snapshots_1_17 = _RAND_111[5:0];
  _RAND_112 = {1{`RANDOM}};
  br_snapshots_1_18 = _RAND_112[5:0];
  _RAND_113 = {1{`RANDOM}};
  br_snapshots_1_19 = _RAND_113[5:0];
  _RAND_114 = {1{`RANDOM}};
  br_snapshots_1_20 = _RAND_114[5:0];
  _RAND_115 = {1{`RANDOM}};
  br_snapshots_1_21 = _RAND_115[5:0];
  _RAND_116 = {1{`RANDOM}};
  br_snapshots_1_22 = _RAND_116[5:0];
  _RAND_117 = {1{`RANDOM}};
  br_snapshots_1_23 = _RAND_117[5:0];
  _RAND_118 = {1{`RANDOM}};
  br_snapshots_1_24 = _RAND_118[5:0];
  _RAND_119 = {1{`RANDOM}};
  br_snapshots_1_25 = _RAND_119[5:0];
  _RAND_120 = {1{`RANDOM}};
  br_snapshots_1_26 = _RAND_120[5:0];
  _RAND_121 = {1{`RANDOM}};
  br_snapshots_1_27 = _RAND_121[5:0];
  _RAND_122 = {1{`RANDOM}};
  br_snapshots_1_28 = _RAND_122[5:0];
  _RAND_123 = {1{`RANDOM}};
  br_snapshots_1_29 = _RAND_123[5:0];
  _RAND_124 = {1{`RANDOM}};
  br_snapshots_1_30 = _RAND_124[5:0];
  _RAND_125 = {1{`RANDOM}};
  br_snapshots_1_31 = _RAND_125[5:0];
  _RAND_126 = {1{`RANDOM}};
  br_snapshots_2_1 = _RAND_126[5:0];
  _RAND_127 = {1{`RANDOM}};
  br_snapshots_2_2 = _RAND_127[5:0];
  _RAND_128 = {1{`RANDOM}};
  br_snapshots_2_3 = _RAND_128[5:0];
  _RAND_129 = {1{`RANDOM}};
  br_snapshots_2_4 = _RAND_129[5:0];
  _RAND_130 = {1{`RANDOM}};
  br_snapshots_2_5 = _RAND_130[5:0];
  _RAND_131 = {1{`RANDOM}};
  br_snapshots_2_6 = _RAND_131[5:0];
  _RAND_132 = {1{`RANDOM}};
  br_snapshots_2_7 = _RAND_132[5:0];
  _RAND_133 = {1{`RANDOM}};
  br_snapshots_2_8 = _RAND_133[5:0];
  _RAND_134 = {1{`RANDOM}};
  br_snapshots_2_9 = _RAND_134[5:0];
  _RAND_135 = {1{`RANDOM}};
  br_snapshots_2_10 = _RAND_135[5:0];
  _RAND_136 = {1{`RANDOM}};
  br_snapshots_2_11 = _RAND_136[5:0];
  _RAND_137 = {1{`RANDOM}};
  br_snapshots_2_12 = _RAND_137[5:0];
  _RAND_138 = {1{`RANDOM}};
  br_snapshots_2_13 = _RAND_138[5:0];
  _RAND_139 = {1{`RANDOM}};
  br_snapshots_2_14 = _RAND_139[5:0];
  _RAND_140 = {1{`RANDOM}};
  br_snapshots_2_15 = _RAND_140[5:0];
  _RAND_141 = {1{`RANDOM}};
  br_snapshots_2_16 = _RAND_141[5:0];
  _RAND_142 = {1{`RANDOM}};
  br_snapshots_2_17 = _RAND_142[5:0];
  _RAND_143 = {1{`RANDOM}};
  br_snapshots_2_18 = _RAND_143[5:0];
  _RAND_144 = {1{`RANDOM}};
  br_snapshots_2_19 = _RAND_144[5:0];
  _RAND_145 = {1{`RANDOM}};
  br_snapshots_2_20 = _RAND_145[5:0];
  _RAND_146 = {1{`RANDOM}};
  br_snapshots_2_21 = _RAND_146[5:0];
  _RAND_147 = {1{`RANDOM}};
  br_snapshots_2_22 = _RAND_147[5:0];
  _RAND_148 = {1{`RANDOM}};
  br_snapshots_2_23 = _RAND_148[5:0];
  _RAND_149 = {1{`RANDOM}};
  br_snapshots_2_24 = _RAND_149[5:0];
  _RAND_150 = {1{`RANDOM}};
  br_snapshots_2_25 = _RAND_150[5:0];
  _RAND_151 = {1{`RANDOM}};
  br_snapshots_2_26 = _RAND_151[5:0];
  _RAND_152 = {1{`RANDOM}};
  br_snapshots_2_27 = _RAND_152[5:0];
  _RAND_153 = {1{`RANDOM}};
  br_snapshots_2_28 = _RAND_153[5:0];
  _RAND_154 = {1{`RANDOM}};
  br_snapshots_2_29 = _RAND_154[5:0];
  _RAND_155 = {1{`RANDOM}};
  br_snapshots_2_30 = _RAND_155[5:0];
  _RAND_156 = {1{`RANDOM}};
  br_snapshots_2_31 = _RAND_156[5:0];
  _RAND_157 = {1{`RANDOM}};
  br_snapshots_3_1 = _RAND_157[5:0];
  _RAND_158 = {1{`RANDOM}};
  br_snapshots_3_2 = _RAND_158[5:0];
  _RAND_159 = {1{`RANDOM}};
  br_snapshots_3_3 = _RAND_159[5:0];
  _RAND_160 = {1{`RANDOM}};
  br_snapshots_3_4 = _RAND_160[5:0];
  _RAND_161 = {1{`RANDOM}};
  br_snapshots_3_5 = _RAND_161[5:0];
  _RAND_162 = {1{`RANDOM}};
  br_snapshots_3_6 = _RAND_162[5:0];
  _RAND_163 = {1{`RANDOM}};
  br_snapshots_3_7 = _RAND_163[5:0];
  _RAND_164 = {1{`RANDOM}};
  br_snapshots_3_8 = _RAND_164[5:0];
  _RAND_165 = {1{`RANDOM}};
  br_snapshots_3_9 = _RAND_165[5:0];
  _RAND_166 = {1{`RANDOM}};
  br_snapshots_3_10 = _RAND_166[5:0];
  _RAND_167 = {1{`RANDOM}};
  br_snapshots_3_11 = _RAND_167[5:0];
  _RAND_168 = {1{`RANDOM}};
  br_snapshots_3_12 = _RAND_168[5:0];
  _RAND_169 = {1{`RANDOM}};
  br_snapshots_3_13 = _RAND_169[5:0];
  _RAND_170 = {1{`RANDOM}};
  br_snapshots_3_14 = _RAND_170[5:0];
  _RAND_171 = {1{`RANDOM}};
  br_snapshots_3_15 = _RAND_171[5:0];
  _RAND_172 = {1{`RANDOM}};
  br_snapshots_3_16 = _RAND_172[5:0];
  _RAND_173 = {1{`RANDOM}};
  br_snapshots_3_17 = _RAND_173[5:0];
  _RAND_174 = {1{`RANDOM}};
  br_snapshots_3_18 = _RAND_174[5:0];
  _RAND_175 = {1{`RANDOM}};
  br_snapshots_3_19 = _RAND_175[5:0];
  _RAND_176 = {1{`RANDOM}};
  br_snapshots_3_20 = _RAND_176[5:0];
  _RAND_177 = {1{`RANDOM}};
  br_snapshots_3_21 = _RAND_177[5:0];
  _RAND_178 = {1{`RANDOM}};
  br_snapshots_3_22 = _RAND_178[5:0];
  _RAND_179 = {1{`RANDOM}};
  br_snapshots_3_23 = _RAND_179[5:0];
  _RAND_180 = {1{`RANDOM}};
  br_snapshots_3_24 = _RAND_180[5:0];
  _RAND_181 = {1{`RANDOM}};
  br_snapshots_3_25 = _RAND_181[5:0];
  _RAND_182 = {1{`RANDOM}};
  br_snapshots_3_26 = _RAND_182[5:0];
  _RAND_183 = {1{`RANDOM}};
  br_snapshots_3_27 = _RAND_183[5:0];
  _RAND_184 = {1{`RANDOM}};
  br_snapshots_3_28 = _RAND_184[5:0];
  _RAND_185 = {1{`RANDOM}};
  br_snapshots_3_29 = _RAND_185[5:0];
  _RAND_186 = {1{`RANDOM}};
  br_snapshots_3_30 = _RAND_186[5:0];
  _RAND_187 = {1{`RANDOM}};
  br_snapshots_3_31 = _RAND_187[5:0];
  _RAND_188 = {1{`RANDOM}};
  br_snapshots_4_1 = _RAND_188[5:0];
  _RAND_189 = {1{`RANDOM}};
  br_snapshots_4_2 = _RAND_189[5:0];
  _RAND_190 = {1{`RANDOM}};
  br_snapshots_4_3 = _RAND_190[5:0];
  _RAND_191 = {1{`RANDOM}};
  br_snapshots_4_4 = _RAND_191[5:0];
  _RAND_192 = {1{`RANDOM}};
  br_snapshots_4_5 = _RAND_192[5:0];
  _RAND_193 = {1{`RANDOM}};
  br_snapshots_4_6 = _RAND_193[5:0];
  _RAND_194 = {1{`RANDOM}};
  br_snapshots_4_7 = _RAND_194[5:0];
  _RAND_195 = {1{`RANDOM}};
  br_snapshots_4_8 = _RAND_195[5:0];
  _RAND_196 = {1{`RANDOM}};
  br_snapshots_4_9 = _RAND_196[5:0];
  _RAND_197 = {1{`RANDOM}};
  br_snapshots_4_10 = _RAND_197[5:0];
  _RAND_198 = {1{`RANDOM}};
  br_snapshots_4_11 = _RAND_198[5:0];
  _RAND_199 = {1{`RANDOM}};
  br_snapshots_4_12 = _RAND_199[5:0];
  _RAND_200 = {1{`RANDOM}};
  br_snapshots_4_13 = _RAND_200[5:0];
  _RAND_201 = {1{`RANDOM}};
  br_snapshots_4_14 = _RAND_201[5:0];
  _RAND_202 = {1{`RANDOM}};
  br_snapshots_4_15 = _RAND_202[5:0];
  _RAND_203 = {1{`RANDOM}};
  br_snapshots_4_16 = _RAND_203[5:0];
  _RAND_204 = {1{`RANDOM}};
  br_snapshots_4_17 = _RAND_204[5:0];
  _RAND_205 = {1{`RANDOM}};
  br_snapshots_4_18 = _RAND_205[5:0];
  _RAND_206 = {1{`RANDOM}};
  br_snapshots_4_19 = _RAND_206[5:0];
  _RAND_207 = {1{`RANDOM}};
  br_snapshots_4_20 = _RAND_207[5:0];
  _RAND_208 = {1{`RANDOM}};
  br_snapshots_4_21 = _RAND_208[5:0];
  _RAND_209 = {1{`RANDOM}};
  br_snapshots_4_22 = _RAND_209[5:0];
  _RAND_210 = {1{`RANDOM}};
  br_snapshots_4_23 = _RAND_210[5:0];
  _RAND_211 = {1{`RANDOM}};
  br_snapshots_4_24 = _RAND_211[5:0];
  _RAND_212 = {1{`RANDOM}};
  br_snapshots_4_25 = _RAND_212[5:0];
  _RAND_213 = {1{`RANDOM}};
  br_snapshots_4_26 = _RAND_213[5:0];
  _RAND_214 = {1{`RANDOM}};
  br_snapshots_4_27 = _RAND_214[5:0];
  _RAND_215 = {1{`RANDOM}};
  br_snapshots_4_28 = _RAND_215[5:0];
  _RAND_216 = {1{`RANDOM}};
  br_snapshots_4_29 = _RAND_216[5:0];
  _RAND_217 = {1{`RANDOM}};
  br_snapshots_4_30 = _RAND_217[5:0];
  _RAND_218 = {1{`RANDOM}};
  br_snapshots_4_31 = _RAND_218[5:0];
  _RAND_219 = {1{`RANDOM}};
  br_snapshots_5_1 = _RAND_219[5:0];
  _RAND_220 = {1{`RANDOM}};
  br_snapshots_5_2 = _RAND_220[5:0];
  _RAND_221 = {1{`RANDOM}};
  br_snapshots_5_3 = _RAND_221[5:0];
  _RAND_222 = {1{`RANDOM}};
  br_snapshots_5_4 = _RAND_222[5:0];
  _RAND_223 = {1{`RANDOM}};
  br_snapshots_5_5 = _RAND_223[5:0];
  _RAND_224 = {1{`RANDOM}};
  br_snapshots_5_6 = _RAND_224[5:0];
  _RAND_225 = {1{`RANDOM}};
  br_snapshots_5_7 = _RAND_225[5:0];
  _RAND_226 = {1{`RANDOM}};
  br_snapshots_5_8 = _RAND_226[5:0];
  _RAND_227 = {1{`RANDOM}};
  br_snapshots_5_9 = _RAND_227[5:0];
  _RAND_228 = {1{`RANDOM}};
  br_snapshots_5_10 = _RAND_228[5:0];
  _RAND_229 = {1{`RANDOM}};
  br_snapshots_5_11 = _RAND_229[5:0];
  _RAND_230 = {1{`RANDOM}};
  br_snapshots_5_12 = _RAND_230[5:0];
  _RAND_231 = {1{`RANDOM}};
  br_snapshots_5_13 = _RAND_231[5:0];
  _RAND_232 = {1{`RANDOM}};
  br_snapshots_5_14 = _RAND_232[5:0];
  _RAND_233 = {1{`RANDOM}};
  br_snapshots_5_15 = _RAND_233[5:0];
  _RAND_234 = {1{`RANDOM}};
  br_snapshots_5_16 = _RAND_234[5:0];
  _RAND_235 = {1{`RANDOM}};
  br_snapshots_5_17 = _RAND_235[5:0];
  _RAND_236 = {1{`RANDOM}};
  br_snapshots_5_18 = _RAND_236[5:0];
  _RAND_237 = {1{`RANDOM}};
  br_snapshots_5_19 = _RAND_237[5:0];
  _RAND_238 = {1{`RANDOM}};
  br_snapshots_5_20 = _RAND_238[5:0];
  _RAND_239 = {1{`RANDOM}};
  br_snapshots_5_21 = _RAND_239[5:0];
  _RAND_240 = {1{`RANDOM}};
  br_snapshots_5_22 = _RAND_240[5:0];
  _RAND_241 = {1{`RANDOM}};
  br_snapshots_5_23 = _RAND_241[5:0];
  _RAND_242 = {1{`RANDOM}};
  br_snapshots_5_24 = _RAND_242[5:0];
  _RAND_243 = {1{`RANDOM}};
  br_snapshots_5_25 = _RAND_243[5:0];
  _RAND_244 = {1{`RANDOM}};
  br_snapshots_5_26 = _RAND_244[5:0];
  _RAND_245 = {1{`RANDOM}};
  br_snapshots_5_27 = _RAND_245[5:0];
  _RAND_246 = {1{`RANDOM}};
  br_snapshots_5_28 = _RAND_246[5:0];
  _RAND_247 = {1{`RANDOM}};
  br_snapshots_5_29 = _RAND_247[5:0];
  _RAND_248 = {1{`RANDOM}};
  br_snapshots_5_30 = _RAND_248[5:0];
  _RAND_249 = {1{`RANDOM}};
  br_snapshots_5_31 = _RAND_249[5:0];
  _RAND_250 = {1{`RANDOM}};
  br_snapshots_6_1 = _RAND_250[5:0];
  _RAND_251 = {1{`RANDOM}};
  br_snapshots_6_2 = _RAND_251[5:0];
  _RAND_252 = {1{`RANDOM}};
  br_snapshots_6_3 = _RAND_252[5:0];
  _RAND_253 = {1{`RANDOM}};
  br_snapshots_6_4 = _RAND_253[5:0];
  _RAND_254 = {1{`RANDOM}};
  br_snapshots_6_5 = _RAND_254[5:0];
  _RAND_255 = {1{`RANDOM}};
  br_snapshots_6_6 = _RAND_255[5:0];
  _RAND_256 = {1{`RANDOM}};
  br_snapshots_6_7 = _RAND_256[5:0];
  _RAND_257 = {1{`RANDOM}};
  br_snapshots_6_8 = _RAND_257[5:0];
  _RAND_258 = {1{`RANDOM}};
  br_snapshots_6_9 = _RAND_258[5:0];
  _RAND_259 = {1{`RANDOM}};
  br_snapshots_6_10 = _RAND_259[5:0];
  _RAND_260 = {1{`RANDOM}};
  br_snapshots_6_11 = _RAND_260[5:0];
  _RAND_261 = {1{`RANDOM}};
  br_snapshots_6_12 = _RAND_261[5:0];
  _RAND_262 = {1{`RANDOM}};
  br_snapshots_6_13 = _RAND_262[5:0];
  _RAND_263 = {1{`RANDOM}};
  br_snapshots_6_14 = _RAND_263[5:0];
  _RAND_264 = {1{`RANDOM}};
  br_snapshots_6_15 = _RAND_264[5:0];
  _RAND_265 = {1{`RANDOM}};
  br_snapshots_6_16 = _RAND_265[5:0];
  _RAND_266 = {1{`RANDOM}};
  br_snapshots_6_17 = _RAND_266[5:0];
  _RAND_267 = {1{`RANDOM}};
  br_snapshots_6_18 = _RAND_267[5:0];
  _RAND_268 = {1{`RANDOM}};
  br_snapshots_6_19 = _RAND_268[5:0];
  _RAND_269 = {1{`RANDOM}};
  br_snapshots_6_20 = _RAND_269[5:0];
  _RAND_270 = {1{`RANDOM}};
  br_snapshots_6_21 = _RAND_270[5:0];
  _RAND_271 = {1{`RANDOM}};
  br_snapshots_6_22 = _RAND_271[5:0];
  _RAND_272 = {1{`RANDOM}};
  br_snapshots_6_23 = _RAND_272[5:0];
  _RAND_273 = {1{`RANDOM}};
  br_snapshots_6_24 = _RAND_273[5:0];
  _RAND_274 = {1{`RANDOM}};
  br_snapshots_6_25 = _RAND_274[5:0];
  _RAND_275 = {1{`RANDOM}};
  br_snapshots_6_26 = _RAND_275[5:0];
  _RAND_276 = {1{`RANDOM}};
  br_snapshots_6_27 = _RAND_276[5:0];
  _RAND_277 = {1{`RANDOM}};
  br_snapshots_6_28 = _RAND_277[5:0];
  _RAND_278 = {1{`RANDOM}};
  br_snapshots_6_29 = _RAND_278[5:0];
  _RAND_279 = {1{`RANDOM}};
  br_snapshots_6_30 = _RAND_279[5:0];
  _RAND_280 = {1{`RANDOM}};
  br_snapshots_6_31 = _RAND_280[5:0];
  _RAND_281 = {1{`RANDOM}};
  br_snapshots_7_1 = _RAND_281[5:0];
  _RAND_282 = {1{`RANDOM}};
  br_snapshots_7_2 = _RAND_282[5:0];
  _RAND_283 = {1{`RANDOM}};
  br_snapshots_7_3 = _RAND_283[5:0];
  _RAND_284 = {1{`RANDOM}};
  br_snapshots_7_4 = _RAND_284[5:0];
  _RAND_285 = {1{`RANDOM}};
  br_snapshots_7_5 = _RAND_285[5:0];
  _RAND_286 = {1{`RANDOM}};
  br_snapshots_7_6 = _RAND_286[5:0];
  _RAND_287 = {1{`RANDOM}};
  br_snapshots_7_7 = _RAND_287[5:0];
  _RAND_288 = {1{`RANDOM}};
  br_snapshots_7_8 = _RAND_288[5:0];
  _RAND_289 = {1{`RANDOM}};
  br_snapshots_7_9 = _RAND_289[5:0];
  _RAND_290 = {1{`RANDOM}};
  br_snapshots_7_10 = _RAND_290[5:0];
  _RAND_291 = {1{`RANDOM}};
  br_snapshots_7_11 = _RAND_291[5:0];
  _RAND_292 = {1{`RANDOM}};
  br_snapshots_7_12 = _RAND_292[5:0];
  _RAND_293 = {1{`RANDOM}};
  br_snapshots_7_13 = _RAND_293[5:0];
  _RAND_294 = {1{`RANDOM}};
  br_snapshots_7_14 = _RAND_294[5:0];
  _RAND_295 = {1{`RANDOM}};
  br_snapshots_7_15 = _RAND_295[5:0];
  _RAND_296 = {1{`RANDOM}};
  br_snapshots_7_16 = _RAND_296[5:0];
  _RAND_297 = {1{`RANDOM}};
  br_snapshots_7_17 = _RAND_297[5:0];
  _RAND_298 = {1{`RANDOM}};
  br_snapshots_7_18 = _RAND_298[5:0];
  _RAND_299 = {1{`RANDOM}};
  br_snapshots_7_19 = _RAND_299[5:0];
  _RAND_300 = {1{`RANDOM}};
  br_snapshots_7_20 = _RAND_300[5:0];
  _RAND_301 = {1{`RANDOM}};
  br_snapshots_7_21 = _RAND_301[5:0];
  _RAND_302 = {1{`RANDOM}};
  br_snapshots_7_22 = _RAND_302[5:0];
  _RAND_303 = {1{`RANDOM}};
  br_snapshots_7_23 = _RAND_303[5:0];
  _RAND_304 = {1{`RANDOM}};
  br_snapshots_7_24 = _RAND_304[5:0];
  _RAND_305 = {1{`RANDOM}};
  br_snapshots_7_25 = _RAND_305[5:0];
  _RAND_306 = {1{`RANDOM}};
  br_snapshots_7_26 = _RAND_306[5:0];
  _RAND_307 = {1{`RANDOM}};
  br_snapshots_7_27 = _RAND_307[5:0];
  _RAND_308 = {1{`RANDOM}};
  br_snapshots_7_28 = _RAND_308[5:0];
  _RAND_309 = {1{`RANDOM}};
  br_snapshots_7_29 = _RAND_309[5:0];
  _RAND_310 = {1{`RANDOM}};
  br_snapshots_7_30 = _RAND_310[5:0];
  _RAND_311 = {1{`RANDOM}};
  br_snapshots_7_31 = _RAND_311[5:0];
  _RAND_312 = {1{`RANDOM}};
  br_snapshots_8_1 = _RAND_312[5:0];
  _RAND_313 = {1{`RANDOM}};
  br_snapshots_8_2 = _RAND_313[5:0];
  _RAND_314 = {1{`RANDOM}};
  br_snapshots_8_3 = _RAND_314[5:0];
  _RAND_315 = {1{`RANDOM}};
  br_snapshots_8_4 = _RAND_315[5:0];
  _RAND_316 = {1{`RANDOM}};
  br_snapshots_8_5 = _RAND_316[5:0];
  _RAND_317 = {1{`RANDOM}};
  br_snapshots_8_6 = _RAND_317[5:0];
  _RAND_318 = {1{`RANDOM}};
  br_snapshots_8_7 = _RAND_318[5:0];
  _RAND_319 = {1{`RANDOM}};
  br_snapshots_8_8 = _RAND_319[5:0];
  _RAND_320 = {1{`RANDOM}};
  br_snapshots_8_9 = _RAND_320[5:0];
  _RAND_321 = {1{`RANDOM}};
  br_snapshots_8_10 = _RAND_321[5:0];
  _RAND_322 = {1{`RANDOM}};
  br_snapshots_8_11 = _RAND_322[5:0];
  _RAND_323 = {1{`RANDOM}};
  br_snapshots_8_12 = _RAND_323[5:0];
  _RAND_324 = {1{`RANDOM}};
  br_snapshots_8_13 = _RAND_324[5:0];
  _RAND_325 = {1{`RANDOM}};
  br_snapshots_8_14 = _RAND_325[5:0];
  _RAND_326 = {1{`RANDOM}};
  br_snapshots_8_15 = _RAND_326[5:0];
  _RAND_327 = {1{`RANDOM}};
  br_snapshots_8_16 = _RAND_327[5:0];
  _RAND_328 = {1{`RANDOM}};
  br_snapshots_8_17 = _RAND_328[5:0];
  _RAND_329 = {1{`RANDOM}};
  br_snapshots_8_18 = _RAND_329[5:0];
  _RAND_330 = {1{`RANDOM}};
  br_snapshots_8_19 = _RAND_330[5:0];
  _RAND_331 = {1{`RANDOM}};
  br_snapshots_8_20 = _RAND_331[5:0];
  _RAND_332 = {1{`RANDOM}};
  br_snapshots_8_21 = _RAND_332[5:0];
  _RAND_333 = {1{`RANDOM}};
  br_snapshots_8_22 = _RAND_333[5:0];
  _RAND_334 = {1{`RANDOM}};
  br_snapshots_8_23 = _RAND_334[5:0];
  _RAND_335 = {1{`RANDOM}};
  br_snapshots_8_24 = _RAND_335[5:0];
  _RAND_336 = {1{`RANDOM}};
  br_snapshots_8_25 = _RAND_336[5:0];
  _RAND_337 = {1{`RANDOM}};
  br_snapshots_8_26 = _RAND_337[5:0];
  _RAND_338 = {1{`RANDOM}};
  br_snapshots_8_27 = _RAND_338[5:0];
  _RAND_339 = {1{`RANDOM}};
  br_snapshots_8_28 = _RAND_339[5:0];
  _RAND_340 = {1{`RANDOM}};
  br_snapshots_8_29 = _RAND_340[5:0];
  _RAND_341 = {1{`RANDOM}};
  br_snapshots_8_30 = _RAND_341[5:0];
  _RAND_342 = {1{`RANDOM}};
  br_snapshots_8_31 = _RAND_342[5:0];
  _RAND_343 = {1{`RANDOM}};
  br_snapshots_9_1 = _RAND_343[5:0];
  _RAND_344 = {1{`RANDOM}};
  br_snapshots_9_2 = _RAND_344[5:0];
  _RAND_345 = {1{`RANDOM}};
  br_snapshots_9_3 = _RAND_345[5:0];
  _RAND_346 = {1{`RANDOM}};
  br_snapshots_9_4 = _RAND_346[5:0];
  _RAND_347 = {1{`RANDOM}};
  br_snapshots_9_5 = _RAND_347[5:0];
  _RAND_348 = {1{`RANDOM}};
  br_snapshots_9_6 = _RAND_348[5:0];
  _RAND_349 = {1{`RANDOM}};
  br_snapshots_9_7 = _RAND_349[5:0];
  _RAND_350 = {1{`RANDOM}};
  br_snapshots_9_8 = _RAND_350[5:0];
  _RAND_351 = {1{`RANDOM}};
  br_snapshots_9_9 = _RAND_351[5:0];
  _RAND_352 = {1{`RANDOM}};
  br_snapshots_9_10 = _RAND_352[5:0];
  _RAND_353 = {1{`RANDOM}};
  br_snapshots_9_11 = _RAND_353[5:0];
  _RAND_354 = {1{`RANDOM}};
  br_snapshots_9_12 = _RAND_354[5:0];
  _RAND_355 = {1{`RANDOM}};
  br_snapshots_9_13 = _RAND_355[5:0];
  _RAND_356 = {1{`RANDOM}};
  br_snapshots_9_14 = _RAND_356[5:0];
  _RAND_357 = {1{`RANDOM}};
  br_snapshots_9_15 = _RAND_357[5:0];
  _RAND_358 = {1{`RANDOM}};
  br_snapshots_9_16 = _RAND_358[5:0];
  _RAND_359 = {1{`RANDOM}};
  br_snapshots_9_17 = _RAND_359[5:0];
  _RAND_360 = {1{`RANDOM}};
  br_snapshots_9_18 = _RAND_360[5:0];
  _RAND_361 = {1{`RANDOM}};
  br_snapshots_9_19 = _RAND_361[5:0];
  _RAND_362 = {1{`RANDOM}};
  br_snapshots_9_20 = _RAND_362[5:0];
  _RAND_363 = {1{`RANDOM}};
  br_snapshots_9_21 = _RAND_363[5:0];
  _RAND_364 = {1{`RANDOM}};
  br_snapshots_9_22 = _RAND_364[5:0];
  _RAND_365 = {1{`RANDOM}};
  br_snapshots_9_23 = _RAND_365[5:0];
  _RAND_366 = {1{`RANDOM}};
  br_snapshots_9_24 = _RAND_366[5:0];
  _RAND_367 = {1{`RANDOM}};
  br_snapshots_9_25 = _RAND_367[5:0];
  _RAND_368 = {1{`RANDOM}};
  br_snapshots_9_26 = _RAND_368[5:0];
  _RAND_369 = {1{`RANDOM}};
  br_snapshots_9_27 = _RAND_369[5:0];
  _RAND_370 = {1{`RANDOM}};
  br_snapshots_9_28 = _RAND_370[5:0];
  _RAND_371 = {1{`RANDOM}};
  br_snapshots_9_29 = _RAND_371[5:0];
  _RAND_372 = {1{`RANDOM}};
  br_snapshots_9_30 = _RAND_372[5:0];
  _RAND_373 = {1{`RANDOM}};
  br_snapshots_9_31 = _RAND_373[5:0];
  _RAND_374 = {1{`RANDOM}};
  br_snapshots_10_1 = _RAND_374[5:0];
  _RAND_375 = {1{`RANDOM}};
  br_snapshots_10_2 = _RAND_375[5:0];
  _RAND_376 = {1{`RANDOM}};
  br_snapshots_10_3 = _RAND_376[5:0];
  _RAND_377 = {1{`RANDOM}};
  br_snapshots_10_4 = _RAND_377[5:0];
  _RAND_378 = {1{`RANDOM}};
  br_snapshots_10_5 = _RAND_378[5:0];
  _RAND_379 = {1{`RANDOM}};
  br_snapshots_10_6 = _RAND_379[5:0];
  _RAND_380 = {1{`RANDOM}};
  br_snapshots_10_7 = _RAND_380[5:0];
  _RAND_381 = {1{`RANDOM}};
  br_snapshots_10_8 = _RAND_381[5:0];
  _RAND_382 = {1{`RANDOM}};
  br_snapshots_10_9 = _RAND_382[5:0];
  _RAND_383 = {1{`RANDOM}};
  br_snapshots_10_10 = _RAND_383[5:0];
  _RAND_384 = {1{`RANDOM}};
  br_snapshots_10_11 = _RAND_384[5:0];
  _RAND_385 = {1{`RANDOM}};
  br_snapshots_10_12 = _RAND_385[5:0];
  _RAND_386 = {1{`RANDOM}};
  br_snapshots_10_13 = _RAND_386[5:0];
  _RAND_387 = {1{`RANDOM}};
  br_snapshots_10_14 = _RAND_387[5:0];
  _RAND_388 = {1{`RANDOM}};
  br_snapshots_10_15 = _RAND_388[5:0];
  _RAND_389 = {1{`RANDOM}};
  br_snapshots_10_16 = _RAND_389[5:0];
  _RAND_390 = {1{`RANDOM}};
  br_snapshots_10_17 = _RAND_390[5:0];
  _RAND_391 = {1{`RANDOM}};
  br_snapshots_10_18 = _RAND_391[5:0];
  _RAND_392 = {1{`RANDOM}};
  br_snapshots_10_19 = _RAND_392[5:0];
  _RAND_393 = {1{`RANDOM}};
  br_snapshots_10_20 = _RAND_393[5:0];
  _RAND_394 = {1{`RANDOM}};
  br_snapshots_10_21 = _RAND_394[5:0];
  _RAND_395 = {1{`RANDOM}};
  br_snapshots_10_22 = _RAND_395[5:0];
  _RAND_396 = {1{`RANDOM}};
  br_snapshots_10_23 = _RAND_396[5:0];
  _RAND_397 = {1{`RANDOM}};
  br_snapshots_10_24 = _RAND_397[5:0];
  _RAND_398 = {1{`RANDOM}};
  br_snapshots_10_25 = _RAND_398[5:0];
  _RAND_399 = {1{`RANDOM}};
  br_snapshots_10_26 = _RAND_399[5:0];
  _RAND_400 = {1{`RANDOM}};
  br_snapshots_10_27 = _RAND_400[5:0];
  _RAND_401 = {1{`RANDOM}};
  br_snapshots_10_28 = _RAND_401[5:0];
  _RAND_402 = {1{`RANDOM}};
  br_snapshots_10_29 = _RAND_402[5:0];
  _RAND_403 = {1{`RANDOM}};
  br_snapshots_10_30 = _RAND_403[5:0];
  _RAND_404 = {1{`RANDOM}};
  br_snapshots_10_31 = _RAND_404[5:0];
  _RAND_405 = {1{`RANDOM}};
  br_snapshots_11_1 = _RAND_405[5:0];
  _RAND_406 = {1{`RANDOM}};
  br_snapshots_11_2 = _RAND_406[5:0];
  _RAND_407 = {1{`RANDOM}};
  br_snapshots_11_3 = _RAND_407[5:0];
  _RAND_408 = {1{`RANDOM}};
  br_snapshots_11_4 = _RAND_408[5:0];
  _RAND_409 = {1{`RANDOM}};
  br_snapshots_11_5 = _RAND_409[5:0];
  _RAND_410 = {1{`RANDOM}};
  br_snapshots_11_6 = _RAND_410[5:0];
  _RAND_411 = {1{`RANDOM}};
  br_snapshots_11_7 = _RAND_411[5:0];
  _RAND_412 = {1{`RANDOM}};
  br_snapshots_11_8 = _RAND_412[5:0];
  _RAND_413 = {1{`RANDOM}};
  br_snapshots_11_9 = _RAND_413[5:0];
  _RAND_414 = {1{`RANDOM}};
  br_snapshots_11_10 = _RAND_414[5:0];
  _RAND_415 = {1{`RANDOM}};
  br_snapshots_11_11 = _RAND_415[5:0];
  _RAND_416 = {1{`RANDOM}};
  br_snapshots_11_12 = _RAND_416[5:0];
  _RAND_417 = {1{`RANDOM}};
  br_snapshots_11_13 = _RAND_417[5:0];
  _RAND_418 = {1{`RANDOM}};
  br_snapshots_11_14 = _RAND_418[5:0];
  _RAND_419 = {1{`RANDOM}};
  br_snapshots_11_15 = _RAND_419[5:0];
  _RAND_420 = {1{`RANDOM}};
  br_snapshots_11_16 = _RAND_420[5:0];
  _RAND_421 = {1{`RANDOM}};
  br_snapshots_11_17 = _RAND_421[5:0];
  _RAND_422 = {1{`RANDOM}};
  br_snapshots_11_18 = _RAND_422[5:0];
  _RAND_423 = {1{`RANDOM}};
  br_snapshots_11_19 = _RAND_423[5:0];
  _RAND_424 = {1{`RANDOM}};
  br_snapshots_11_20 = _RAND_424[5:0];
  _RAND_425 = {1{`RANDOM}};
  br_snapshots_11_21 = _RAND_425[5:0];
  _RAND_426 = {1{`RANDOM}};
  br_snapshots_11_22 = _RAND_426[5:0];
  _RAND_427 = {1{`RANDOM}};
  br_snapshots_11_23 = _RAND_427[5:0];
  _RAND_428 = {1{`RANDOM}};
  br_snapshots_11_24 = _RAND_428[5:0];
  _RAND_429 = {1{`RANDOM}};
  br_snapshots_11_25 = _RAND_429[5:0];
  _RAND_430 = {1{`RANDOM}};
  br_snapshots_11_26 = _RAND_430[5:0];
  _RAND_431 = {1{`RANDOM}};
  br_snapshots_11_27 = _RAND_431[5:0];
  _RAND_432 = {1{`RANDOM}};
  br_snapshots_11_28 = _RAND_432[5:0];
  _RAND_433 = {1{`RANDOM}};
  br_snapshots_11_29 = _RAND_433[5:0];
  _RAND_434 = {1{`RANDOM}};
  br_snapshots_11_30 = _RAND_434[5:0];
  _RAND_435 = {1{`RANDOM}};
  br_snapshots_11_31 = _RAND_435[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
