module IssueUnitCollapsing_1(
  input         clock,
  input         reset,
  output        io_dis_uops_0_ready,
  input         io_dis_uops_0_valid,
  input  [6:0]  io_dis_uops_0_bits_uopc,
  input  [31:0] io_dis_uops_0_bits_inst,
  input  [31:0] io_dis_uops_0_bits_debug_inst,
  input         io_dis_uops_0_bits_is_rvc,
  input  [39:0] io_dis_uops_0_bits_debug_pc,
  input  [2:0]  io_dis_uops_0_bits_iq_type,
  input  [9:0]  io_dis_uops_0_bits_fu_code,
  input  [3:0]  io_dis_uops_0_bits_ctrl_br_type,
  input  [1:0]  io_dis_uops_0_bits_ctrl_op1_sel,
  input  [2:0]  io_dis_uops_0_bits_ctrl_op2_sel,
  input  [2:0]  io_dis_uops_0_bits_ctrl_imm_sel,
  input  [3:0]  io_dis_uops_0_bits_ctrl_op_fcn,
  input         io_dis_uops_0_bits_ctrl_fcn_dw,
  input  [2:0]  io_dis_uops_0_bits_ctrl_csr_cmd,
  input         io_dis_uops_0_bits_ctrl_is_load,
  input         io_dis_uops_0_bits_ctrl_is_sta,
  input         io_dis_uops_0_bits_ctrl_is_std,
  input  [1:0]  io_dis_uops_0_bits_iw_state,
  input         io_dis_uops_0_bits_iw_p1_poisoned,
  input         io_dis_uops_0_bits_iw_p2_poisoned,
  input         io_dis_uops_0_bits_is_br,
  input         io_dis_uops_0_bits_is_jalr,
  input         io_dis_uops_0_bits_is_jal,
  input         io_dis_uops_0_bits_is_sfb,
  input  [11:0] io_dis_uops_0_bits_br_mask,
  input  [3:0]  io_dis_uops_0_bits_br_tag,
  input  [4:0]  io_dis_uops_0_bits_ftq_idx,
  input         io_dis_uops_0_bits_edge_inst,
  input  [5:0]  io_dis_uops_0_bits_pc_lob,
  input         io_dis_uops_0_bits_taken,
  input  [19:0] io_dis_uops_0_bits_imm_packed,
  input  [11:0] io_dis_uops_0_bits_csr_addr,
  input  [5:0]  io_dis_uops_0_bits_rob_idx,
  input  [3:0]  io_dis_uops_0_bits_ldq_idx,
  input  [3:0]  io_dis_uops_0_bits_stq_idx,
  input  [1:0]  io_dis_uops_0_bits_rxq_idx,
  input  [5:0]  io_dis_uops_0_bits_pdst,
  input  [5:0]  io_dis_uops_0_bits_prs1,
  input  [5:0]  io_dis_uops_0_bits_prs2,
  input  [5:0]  io_dis_uops_0_bits_prs3,
  input  [4:0]  io_dis_uops_0_bits_ppred,
  input         io_dis_uops_0_bits_prs1_busy,
  input         io_dis_uops_0_bits_prs2_busy,
  input         io_dis_uops_0_bits_prs3_busy,
  input         io_dis_uops_0_bits_ppred_busy,
  input  [5:0]  io_dis_uops_0_bits_stale_pdst,
  input         io_dis_uops_0_bits_exception,
  input  [63:0] io_dis_uops_0_bits_exc_cause,
  input         io_dis_uops_0_bits_bypassable,
  input  [4:0]  io_dis_uops_0_bits_mem_cmd,
  input  [1:0]  io_dis_uops_0_bits_mem_size,
  input         io_dis_uops_0_bits_mem_signed,
  input         io_dis_uops_0_bits_is_fence,
  input         io_dis_uops_0_bits_is_fencei,
  input         io_dis_uops_0_bits_is_amo,
  input         io_dis_uops_0_bits_uses_ldq,
  input         io_dis_uops_0_bits_uses_stq,
  input         io_dis_uops_0_bits_is_sys_pc2epc,
  input         io_dis_uops_0_bits_is_unique,
  input         io_dis_uops_0_bits_flush_on_commit,
  input         io_dis_uops_0_bits_ldst_is_rs1,
  input  [5:0]  io_dis_uops_0_bits_ldst,
  input  [5:0]  io_dis_uops_0_bits_lrs1,
  input  [5:0]  io_dis_uops_0_bits_lrs2,
  input  [5:0]  io_dis_uops_0_bits_lrs3,
  input         io_dis_uops_0_bits_ldst_val,
  input  [1:0]  io_dis_uops_0_bits_dst_rtype,
  input  [1:0]  io_dis_uops_0_bits_lrs1_rtype,
  input  [1:0]  io_dis_uops_0_bits_lrs2_rtype,
  input         io_dis_uops_0_bits_frs3_en,
  input         io_dis_uops_0_bits_fp_val,
  input         io_dis_uops_0_bits_fp_single,
  input         io_dis_uops_0_bits_xcpt_pf_if,
  input         io_dis_uops_0_bits_xcpt_ae_if,
  input         io_dis_uops_0_bits_xcpt_ma_if,
  input         io_dis_uops_0_bits_bp_debug_if,
  input         io_dis_uops_0_bits_bp_xcpt_if,
  input  [1:0]  io_dis_uops_0_bits_debug_fsrc,
  input  [1:0]  io_dis_uops_0_bits_debug_tsrc,
  output        io_dis_uops_1_ready,
  input         io_dis_uops_1_valid,
  input  [6:0]  io_dis_uops_1_bits_uopc,
  input  [31:0] io_dis_uops_1_bits_inst,
  input  [31:0] io_dis_uops_1_bits_debug_inst,
  input         io_dis_uops_1_bits_is_rvc,
  input  [39:0] io_dis_uops_1_bits_debug_pc,
  input  [2:0]  io_dis_uops_1_bits_iq_type,
  input  [9:0]  io_dis_uops_1_bits_fu_code,
  input  [3:0]  io_dis_uops_1_bits_ctrl_br_type,
  input  [1:0]  io_dis_uops_1_bits_ctrl_op1_sel,
  input  [2:0]  io_dis_uops_1_bits_ctrl_op2_sel,
  input  [2:0]  io_dis_uops_1_bits_ctrl_imm_sel,
  input  [3:0]  io_dis_uops_1_bits_ctrl_op_fcn,
  input         io_dis_uops_1_bits_ctrl_fcn_dw,
  input  [2:0]  io_dis_uops_1_bits_ctrl_csr_cmd,
  input         io_dis_uops_1_bits_ctrl_is_load,
  input         io_dis_uops_1_bits_ctrl_is_sta,
  input         io_dis_uops_1_bits_ctrl_is_std,
  input  [1:0]  io_dis_uops_1_bits_iw_state,
  input         io_dis_uops_1_bits_iw_p1_poisoned,
  input         io_dis_uops_1_bits_iw_p2_poisoned,
  input         io_dis_uops_1_bits_is_br,
  input         io_dis_uops_1_bits_is_jalr,
  input         io_dis_uops_1_bits_is_jal,
  input         io_dis_uops_1_bits_is_sfb,
  input  [11:0] io_dis_uops_1_bits_br_mask,
  input  [3:0]  io_dis_uops_1_bits_br_tag,
  input  [4:0]  io_dis_uops_1_bits_ftq_idx,
  input         io_dis_uops_1_bits_edge_inst,
  input  [5:0]  io_dis_uops_1_bits_pc_lob,
  input         io_dis_uops_1_bits_taken,
  input  [19:0] io_dis_uops_1_bits_imm_packed,
  input  [11:0] io_dis_uops_1_bits_csr_addr,
  input  [5:0]  io_dis_uops_1_bits_rob_idx,
  input  [3:0]  io_dis_uops_1_bits_ldq_idx,
  input  [3:0]  io_dis_uops_1_bits_stq_idx,
  input  [1:0]  io_dis_uops_1_bits_rxq_idx,
  input  [5:0]  io_dis_uops_1_bits_pdst,
  input  [5:0]  io_dis_uops_1_bits_prs1,
  input  [5:0]  io_dis_uops_1_bits_prs2,
  input  [5:0]  io_dis_uops_1_bits_prs3,
  input  [4:0]  io_dis_uops_1_bits_ppred,
  input         io_dis_uops_1_bits_prs1_busy,
  input         io_dis_uops_1_bits_prs2_busy,
  input         io_dis_uops_1_bits_prs3_busy,
  input         io_dis_uops_1_bits_ppred_busy,
  input  [5:0]  io_dis_uops_1_bits_stale_pdst,
  input         io_dis_uops_1_bits_exception,
  input  [63:0] io_dis_uops_1_bits_exc_cause,
  input         io_dis_uops_1_bits_bypassable,
  input  [4:0]  io_dis_uops_1_bits_mem_cmd,
  input  [1:0]  io_dis_uops_1_bits_mem_size,
  input         io_dis_uops_1_bits_mem_signed,
  input         io_dis_uops_1_bits_is_fence,
  input         io_dis_uops_1_bits_is_fencei,
  input         io_dis_uops_1_bits_is_amo,
  input         io_dis_uops_1_bits_uses_ldq,
  input         io_dis_uops_1_bits_uses_stq,
  input         io_dis_uops_1_bits_is_sys_pc2epc,
  input         io_dis_uops_1_bits_is_unique,
  input         io_dis_uops_1_bits_flush_on_commit,
  input         io_dis_uops_1_bits_ldst_is_rs1,
  input  [5:0]  io_dis_uops_1_bits_ldst,
  input  [5:0]  io_dis_uops_1_bits_lrs1,
  input  [5:0]  io_dis_uops_1_bits_lrs2,
  input  [5:0]  io_dis_uops_1_bits_lrs3,
  input         io_dis_uops_1_bits_ldst_val,
  input  [1:0]  io_dis_uops_1_bits_dst_rtype,
  input  [1:0]  io_dis_uops_1_bits_lrs1_rtype,
  input  [1:0]  io_dis_uops_1_bits_lrs2_rtype,
  input         io_dis_uops_1_bits_frs3_en,
  input         io_dis_uops_1_bits_fp_val,
  input         io_dis_uops_1_bits_fp_single,
  input         io_dis_uops_1_bits_xcpt_pf_if,
  input         io_dis_uops_1_bits_xcpt_ae_if,
  input         io_dis_uops_1_bits_xcpt_ma_if,
  input         io_dis_uops_1_bits_bp_debug_if,
  input         io_dis_uops_1_bits_bp_xcpt_if,
  input  [1:0]  io_dis_uops_1_bits_debug_fsrc,
  input  [1:0]  io_dis_uops_1_bits_debug_tsrc,
  output        io_iss_valids_0,
  output [6:0]  io_iss_uops_0_uopc,
  output [31:0] io_iss_uops_0_inst,
  output [31:0] io_iss_uops_0_debug_inst,
  output        io_iss_uops_0_is_rvc,
  output [39:0] io_iss_uops_0_debug_pc,
  output [2:0]  io_iss_uops_0_iq_type,
  output [9:0]  io_iss_uops_0_fu_code,
  output [3:0]  io_iss_uops_0_ctrl_br_type,
  output [1:0]  io_iss_uops_0_ctrl_op1_sel,
  output [2:0]  io_iss_uops_0_ctrl_op2_sel,
  output [2:0]  io_iss_uops_0_ctrl_imm_sel,
  output [3:0]  io_iss_uops_0_ctrl_op_fcn,
  output        io_iss_uops_0_ctrl_fcn_dw,
  output [2:0]  io_iss_uops_0_ctrl_csr_cmd,
  output        io_iss_uops_0_ctrl_is_load,
  output        io_iss_uops_0_ctrl_is_sta,
  output        io_iss_uops_0_ctrl_is_std,
  output [1:0]  io_iss_uops_0_iw_state,
  output        io_iss_uops_0_iw_p1_poisoned,
  output        io_iss_uops_0_iw_p2_poisoned,
  output        io_iss_uops_0_is_br,
  output        io_iss_uops_0_is_jalr,
  output        io_iss_uops_0_is_jal,
  output        io_iss_uops_0_is_sfb,
  output [11:0] io_iss_uops_0_br_mask,
  output [3:0]  io_iss_uops_0_br_tag,
  output [4:0]  io_iss_uops_0_ftq_idx,
  output        io_iss_uops_0_edge_inst,
  output [5:0]  io_iss_uops_0_pc_lob,
  output        io_iss_uops_0_taken,
  output [19:0] io_iss_uops_0_imm_packed,
  output [11:0] io_iss_uops_0_csr_addr,
  output [5:0]  io_iss_uops_0_rob_idx,
  output [3:0]  io_iss_uops_0_ldq_idx,
  output [3:0]  io_iss_uops_0_stq_idx,
  output [1:0]  io_iss_uops_0_rxq_idx,
  output [5:0]  io_iss_uops_0_pdst,
  output [5:0]  io_iss_uops_0_prs1,
  output [5:0]  io_iss_uops_0_prs2,
  output [5:0]  io_iss_uops_0_prs3,
  output [4:0]  io_iss_uops_0_ppred,
  output        io_iss_uops_0_prs1_busy,
  output        io_iss_uops_0_prs2_busy,
  output        io_iss_uops_0_prs3_busy,
  output        io_iss_uops_0_ppred_busy,
  output [5:0]  io_iss_uops_0_stale_pdst,
  output        io_iss_uops_0_exception,
  output [63:0] io_iss_uops_0_exc_cause,
  output        io_iss_uops_0_bypassable,
  output [4:0]  io_iss_uops_0_mem_cmd,
  output [1:0]  io_iss_uops_0_mem_size,
  output        io_iss_uops_0_mem_signed,
  output        io_iss_uops_0_is_fence,
  output        io_iss_uops_0_is_fencei,
  output        io_iss_uops_0_is_amo,
  output        io_iss_uops_0_uses_ldq,
  output        io_iss_uops_0_uses_stq,
  output        io_iss_uops_0_is_sys_pc2epc,
  output        io_iss_uops_0_is_unique,
  output        io_iss_uops_0_flush_on_commit,
  output        io_iss_uops_0_ldst_is_rs1,
  output [5:0]  io_iss_uops_0_ldst,
  output [5:0]  io_iss_uops_0_lrs1,
  output [5:0]  io_iss_uops_0_lrs2,
  output [5:0]  io_iss_uops_0_lrs3,
  output        io_iss_uops_0_ldst_val,
  output [1:0]  io_iss_uops_0_dst_rtype,
  output [1:0]  io_iss_uops_0_lrs1_rtype,
  output [1:0]  io_iss_uops_0_lrs2_rtype,
  output        io_iss_uops_0_frs3_en,
  output        io_iss_uops_0_fp_val,
  output        io_iss_uops_0_fp_single,
  output        io_iss_uops_0_xcpt_pf_if,
  output        io_iss_uops_0_xcpt_ae_if,
  output        io_iss_uops_0_xcpt_ma_if,
  output        io_iss_uops_0_bp_debug_if,
  output        io_iss_uops_0_bp_xcpt_if,
  output [1:0]  io_iss_uops_0_debug_fsrc,
  output [1:0]  io_iss_uops_0_debug_tsrc,
  input         io_wakeup_ports_0_valid,
  input  [5:0]  io_wakeup_ports_0_bits_pdst,
  input         io_wakeup_ports_0_bits_poisoned,
  input         io_wakeup_ports_1_valid,
  input  [5:0]  io_wakeup_ports_1_bits_pdst,
  input         io_wakeup_ports_1_bits_poisoned,
  input         io_wakeup_ports_2_valid,
  input  [5:0]  io_wakeup_ports_2_bits_pdst,
  input         io_wakeup_ports_2_bits_poisoned,
  input         io_wakeup_ports_3_valid,
  input  [5:0]  io_wakeup_ports_3_bits_pdst,
  input         io_wakeup_ports_3_bits_poisoned,
  input         io_wakeup_ports_4_valid,
  input  [5:0]  io_wakeup_ports_4_bits_pdst,
  input         io_wakeup_ports_4_bits_poisoned,
  input         io_pred_wakeup_port_valid,
  input  [4:0]  io_pred_wakeup_port_bits,
  input         io_spec_ld_wakeup_0_valid,
  input  [5:0]  io_spec_ld_wakeup_0_bits,
  input  [9:0]  io_fu_types_0,
  input  [11:0] io_brupdate_b1_resolve_mask,
  input  [11:0] io_brupdate_b1_mispredict_mask,
  input  [6:0]  io_brupdate_b2_uop_uopc,
  input  [31:0] io_brupdate_b2_uop_inst,
  input  [31:0] io_brupdate_b2_uop_debug_inst,
  input         io_brupdate_b2_uop_is_rvc,
  input  [39:0] io_brupdate_b2_uop_debug_pc,
  input  [2:0]  io_brupdate_b2_uop_iq_type,
  input  [9:0]  io_brupdate_b2_uop_fu_code,
  input  [3:0]  io_brupdate_b2_uop_ctrl_br_type,
  input  [1:0]  io_brupdate_b2_uop_ctrl_op1_sel,
  input  [2:0]  io_brupdate_b2_uop_ctrl_op2_sel,
  input  [2:0]  io_brupdate_b2_uop_ctrl_imm_sel,
  input  [3:0]  io_brupdate_b2_uop_ctrl_op_fcn,
  input         io_brupdate_b2_uop_ctrl_fcn_dw,
  input  [2:0]  io_brupdate_b2_uop_ctrl_csr_cmd,
  input         io_brupdate_b2_uop_ctrl_is_load,
  input         io_brupdate_b2_uop_ctrl_is_sta,
  input         io_brupdate_b2_uop_ctrl_is_std,
  input  [1:0]  io_brupdate_b2_uop_iw_state,
  input         io_brupdate_b2_uop_iw_p1_poisoned,
  input         io_brupdate_b2_uop_iw_p2_poisoned,
  input         io_brupdate_b2_uop_is_br,
  input         io_brupdate_b2_uop_is_jalr,
  input         io_brupdate_b2_uop_is_jal,
  input         io_brupdate_b2_uop_is_sfb,
  input  [11:0] io_brupdate_b2_uop_br_mask,
  input  [3:0]  io_brupdate_b2_uop_br_tag,
  input  [4:0]  io_brupdate_b2_uop_ftq_idx,
  input         io_brupdate_b2_uop_edge_inst,
  input  [5:0]  io_brupdate_b2_uop_pc_lob,
  input         io_brupdate_b2_uop_taken,
  input  [19:0] io_brupdate_b2_uop_imm_packed,
  input  [11:0] io_brupdate_b2_uop_csr_addr,
  input  [5:0]  io_brupdate_b2_uop_rob_idx,
  input  [3:0]  io_brupdate_b2_uop_ldq_idx,
  input  [3:0]  io_brupdate_b2_uop_stq_idx,
  input  [1:0]  io_brupdate_b2_uop_rxq_idx,
  input  [5:0]  io_brupdate_b2_uop_pdst,
  input  [5:0]  io_brupdate_b2_uop_prs1,
  input  [5:0]  io_brupdate_b2_uop_prs2,
  input  [5:0]  io_brupdate_b2_uop_prs3,
  input  [4:0]  io_brupdate_b2_uop_ppred,
  input         io_brupdate_b2_uop_prs1_busy,
  input         io_brupdate_b2_uop_prs2_busy,
  input         io_brupdate_b2_uop_prs3_busy,
  input         io_brupdate_b2_uop_ppred_busy,
  input  [5:0]  io_brupdate_b2_uop_stale_pdst,
  input         io_brupdate_b2_uop_exception,
  input  [63:0] io_brupdate_b2_uop_exc_cause,
  input         io_brupdate_b2_uop_bypassable,
  input  [4:0]  io_brupdate_b2_uop_mem_cmd,
  input  [1:0]  io_brupdate_b2_uop_mem_size,
  input         io_brupdate_b2_uop_mem_signed,
  input         io_brupdate_b2_uop_is_fence,
  input         io_brupdate_b2_uop_is_fencei,
  input         io_brupdate_b2_uop_is_amo,
  input         io_brupdate_b2_uop_uses_ldq,
  input         io_brupdate_b2_uop_uses_stq,
  input         io_brupdate_b2_uop_is_sys_pc2epc,
  input         io_brupdate_b2_uop_is_unique,
  input         io_brupdate_b2_uop_flush_on_commit,
  input         io_brupdate_b2_uop_ldst_is_rs1,
  input  [5:0]  io_brupdate_b2_uop_ldst,
  input  [5:0]  io_brupdate_b2_uop_lrs1,
  input  [5:0]  io_brupdate_b2_uop_lrs2,
  input  [5:0]  io_brupdate_b2_uop_lrs3,
  input         io_brupdate_b2_uop_ldst_val,
  input  [1:0]  io_brupdate_b2_uop_dst_rtype,
  input  [1:0]  io_brupdate_b2_uop_lrs1_rtype,
  input  [1:0]  io_brupdate_b2_uop_lrs2_rtype,
  input         io_brupdate_b2_uop_frs3_en,
  input         io_brupdate_b2_uop_fp_val,
  input         io_brupdate_b2_uop_fp_single,
  input         io_brupdate_b2_uop_xcpt_pf_if,
  input         io_brupdate_b2_uop_xcpt_ae_if,
  input         io_brupdate_b2_uop_xcpt_ma_if,
  input         io_brupdate_b2_uop_bp_debug_if,
  input         io_brupdate_b2_uop_bp_xcpt_if,
  input  [1:0]  io_brupdate_b2_uop_debug_fsrc,
  input  [1:0]  io_brupdate_b2_uop_debug_tsrc,
  input         io_brupdate_b2_valid,
  input         io_brupdate_b2_mispredict,
  input         io_brupdate_b2_taken,
  input  [2:0]  io_brupdate_b2_cfi_type,
  input  [1:0]  io_brupdate_b2_pc_sel,
  input  [39:0] io_brupdate_b2_jalr_target,
  input  [20:0] io_brupdate_b2_target_offset,
  input         io_flush_pipeline,
  input         io_ld_miss,
  output        io_event_empty,
  input  [63:0] io_tsc_reg
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  slots_0_clock; // @[issue-unit.scala 153:73]
  wire  slots_0_reset; // @[issue-unit.scala 153:73]
  wire  slots_0_io_valid; // @[issue-unit.scala 153:73]
  wire  slots_0_io_will_be_valid; // @[issue-unit.scala 153:73]
  wire  slots_0_io_request; // @[issue-unit.scala 153:73]
  wire  slots_0_io_request_hp; // @[issue-unit.scala 153:73]
  wire  slots_0_io_grant; // @[issue-unit.scala 153:73]
  wire [11:0] slots_0_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 153:73]
  wire [11:0] slots_0_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 153:73]
  wire [6:0] slots_0_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_0_io_brupdate_b2_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_0_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_0_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_0_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_0_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_0_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_0_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_0_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_0_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_0_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_0_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_0_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_0_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_0_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_0_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_0_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_0_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_0_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_0_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_0_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_valid; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_mispredict; // @[issue-unit.scala 153:73]
  wire  slots_0_io_brupdate_b2_taken; // @[issue-unit.scala 153:73]
  wire [2:0] slots_0_io_brupdate_b2_cfi_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_brupdate_b2_pc_sel; // @[issue-unit.scala 153:73]
  wire [39:0] slots_0_io_brupdate_b2_jalr_target; // @[issue-unit.scala 153:73]
  wire [20:0] slots_0_io_brupdate_b2_target_offset; // @[issue-unit.scala 153:73]
  wire  slots_0_io_kill; // @[issue-unit.scala 153:73]
  wire  slots_0_io_clear; // @[issue-unit.scala 153:73]
  wire  slots_0_io_ldspec_miss; // @[issue-unit.scala 153:73]
  wire  slots_0_io_wakeup_ports_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_0_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_0_io_wakeup_ports_1_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_0_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_0_io_wakeup_ports_2_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_0_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_0_io_wakeup_ports_3_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_0_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_0_io_wakeup_ports_4_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_0_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_0_io_pred_wakeup_port_valid; // @[issue-unit.scala 153:73]
  wire [4:0] slots_0_io_pred_wakeup_port_bits; // @[issue-unit.scala 153:73]
  wire  slots_0_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_valid; // @[issue-unit.scala 153:73]
  wire [6:0] slots_0_io_in_uop_bits_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_0_io_in_uop_bits_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_0_io_in_uop_bits_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_0_io_in_uop_bits_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_0_io_in_uop_bits_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_0_io_in_uop_bits_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_0_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_0_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_0_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_0_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_0_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_in_uop_bits_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_is_br; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_0_io_in_uop_bits_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_0_io_in_uop_bits_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_0_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_in_uop_bits_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_0_io_in_uop_bits_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_0_io_in_uop_bits_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_in_uop_bits_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_0_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_0_io_in_uop_bits_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_in_uop_bits_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_in_uop_bits_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_in_uop_bits_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_in_uop_bits_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_0_io_in_uop_bits_ppred; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_0_io_in_uop_bits_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_0_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_in_uop_bits_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_in_uop_bits_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_in_uop_bits_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_in_uop_bits_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_in_uop_bits_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_0_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_0_io_out_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_0_io_out_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_0_io_out_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_0_io_out_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_0_io_out_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_0_io_out_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_0_io_out_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_0_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_0_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_0_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_0_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_out_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_0_io_out_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_0_io_out_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_0_io_out_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_out_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_0_io_out_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_0_io_out_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_out_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_0_io_out_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_0_io_out_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_out_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_out_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_out_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_out_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_out_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_0_io_out_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_out_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_0_io_out_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_0_io_out_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_out_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_out_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_out_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_out_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_out_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_out_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_out_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_out_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_0_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_out_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_out_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_0_io_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_0_io_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_0_io_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_0_io_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_0_io_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_0_io_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_0_io_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_0_io_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_0_io_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_0_io_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_0_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_0_io_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_0_io_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_0_io_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_0_io_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_0_io_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_0_io_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_0_io_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_0_io_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_0_io_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_0_io_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_0_io_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_0_io_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_0_io_debug_p1; // @[issue-unit.scala 153:73]
  wire  slots_0_io_debug_p2; // @[issue-unit.scala 153:73]
  wire  slots_0_io_debug_p3; // @[issue-unit.scala 153:73]
  wire  slots_0_io_debug_ppred; // @[issue-unit.scala 153:73]
  wire [1:0] slots_0_io_debug_state; // @[issue-unit.scala 153:73]
  wire  slots_1_clock; // @[issue-unit.scala 153:73]
  wire  slots_1_reset; // @[issue-unit.scala 153:73]
  wire  slots_1_io_valid; // @[issue-unit.scala 153:73]
  wire  slots_1_io_will_be_valid; // @[issue-unit.scala 153:73]
  wire  slots_1_io_request; // @[issue-unit.scala 153:73]
  wire  slots_1_io_request_hp; // @[issue-unit.scala 153:73]
  wire  slots_1_io_grant; // @[issue-unit.scala 153:73]
  wire [11:0] slots_1_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 153:73]
  wire [11:0] slots_1_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 153:73]
  wire [6:0] slots_1_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_1_io_brupdate_b2_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_1_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_1_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_1_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_1_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_1_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_1_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_1_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_1_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_1_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_1_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_1_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_1_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_1_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_1_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_1_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_1_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_1_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_1_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_1_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_valid; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_mispredict; // @[issue-unit.scala 153:73]
  wire  slots_1_io_brupdate_b2_taken; // @[issue-unit.scala 153:73]
  wire [2:0] slots_1_io_brupdate_b2_cfi_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_brupdate_b2_pc_sel; // @[issue-unit.scala 153:73]
  wire [39:0] slots_1_io_brupdate_b2_jalr_target; // @[issue-unit.scala 153:73]
  wire [20:0] slots_1_io_brupdate_b2_target_offset; // @[issue-unit.scala 153:73]
  wire  slots_1_io_kill; // @[issue-unit.scala 153:73]
  wire  slots_1_io_clear; // @[issue-unit.scala 153:73]
  wire  slots_1_io_ldspec_miss; // @[issue-unit.scala 153:73]
  wire  slots_1_io_wakeup_ports_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_1_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_1_io_wakeup_ports_1_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_1_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_1_io_wakeup_ports_2_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_1_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_1_io_wakeup_ports_3_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_1_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_1_io_wakeup_ports_4_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_1_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_1_io_pred_wakeup_port_valid; // @[issue-unit.scala 153:73]
  wire [4:0] slots_1_io_pred_wakeup_port_bits; // @[issue-unit.scala 153:73]
  wire  slots_1_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_valid; // @[issue-unit.scala 153:73]
  wire [6:0] slots_1_io_in_uop_bits_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_1_io_in_uop_bits_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_1_io_in_uop_bits_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_1_io_in_uop_bits_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_1_io_in_uop_bits_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_1_io_in_uop_bits_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_1_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_1_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_1_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_1_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_1_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_in_uop_bits_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_is_br; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_1_io_in_uop_bits_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_1_io_in_uop_bits_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_1_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_in_uop_bits_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_1_io_in_uop_bits_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_1_io_in_uop_bits_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_in_uop_bits_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_1_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_1_io_in_uop_bits_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_in_uop_bits_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_in_uop_bits_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_in_uop_bits_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_in_uop_bits_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_1_io_in_uop_bits_ppred; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_1_io_in_uop_bits_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_1_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_in_uop_bits_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_in_uop_bits_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_in_uop_bits_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_in_uop_bits_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_in_uop_bits_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_1_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_1_io_out_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_1_io_out_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_1_io_out_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_1_io_out_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_1_io_out_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_1_io_out_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_1_io_out_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_1_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_1_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_1_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_1_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_out_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_1_io_out_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_1_io_out_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_1_io_out_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_out_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_1_io_out_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_1_io_out_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_out_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_1_io_out_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_1_io_out_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_out_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_out_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_out_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_out_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_out_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_1_io_out_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_out_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_1_io_out_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_1_io_out_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_out_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_out_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_out_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_out_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_out_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_out_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_out_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_out_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_1_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_out_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_out_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_1_io_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_1_io_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_1_io_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_1_io_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_1_io_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_1_io_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_1_io_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_1_io_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_1_io_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_1_io_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_1_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_1_io_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_1_io_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_1_io_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_1_io_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_1_io_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_1_io_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_1_io_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_1_io_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_1_io_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_1_io_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_1_io_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_1_io_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_1_io_debug_p1; // @[issue-unit.scala 153:73]
  wire  slots_1_io_debug_p2; // @[issue-unit.scala 153:73]
  wire  slots_1_io_debug_p3; // @[issue-unit.scala 153:73]
  wire  slots_1_io_debug_ppred; // @[issue-unit.scala 153:73]
  wire [1:0] slots_1_io_debug_state; // @[issue-unit.scala 153:73]
  wire  slots_2_clock; // @[issue-unit.scala 153:73]
  wire  slots_2_reset; // @[issue-unit.scala 153:73]
  wire  slots_2_io_valid; // @[issue-unit.scala 153:73]
  wire  slots_2_io_will_be_valid; // @[issue-unit.scala 153:73]
  wire  slots_2_io_request; // @[issue-unit.scala 153:73]
  wire  slots_2_io_request_hp; // @[issue-unit.scala 153:73]
  wire  slots_2_io_grant; // @[issue-unit.scala 153:73]
  wire [11:0] slots_2_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 153:73]
  wire [11:0] slots_2_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 153:73]
  wire [6:0] slots_2_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_2_io_brupdate_b2_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_2_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_2_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_2_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_2_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_2_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_2_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_2_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_2_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_2_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_2_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_2_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_2_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_2_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_2_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_2_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_2_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_2_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_2_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_2_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_valid; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_mispredict; // @[issue-unit.scala 153:73]
  wire  slots_2_io_brupdate_b2_taken; // @[issue-unit.scala 153:73]
  wire [2:0] slots_2_io_brupdate_b2_cfi_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_brupdate_b2_pc_sel; // @[issue-unit.scala 153:73]
  wire [39:0] slots_2_io_brupdate_b2_jalr_target; // @[issue-unit.scala 153:73]
  wire [20:0] slots_2_io_brupdate_b2_target_offset; // @[issue-unit.scala 153:73]
  wire  slots_2_io_kill; // @[issue-unit.scala 153:73]
  wire  slots_2_io_clear; // @[issue-unit.scala 153:73]
  wire  slots_2_io_ldspec_miss; // @[issue-unit.scala 153:73]
  wire  slots_2_io_wakeup_ports_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_2_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_2_io_wakeup_ports_1_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_2_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_2_io_wakeup_ports_2_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_2_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_2_io_wakeup_ports_3_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_2_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_2_io_wakeup_ports_4_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_2_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_2_io_pred_wakeup_port_valid; // @[issue-unit.scala 153:73]
  wire [4:0] slots_2_io_pred_wakeup_port_bits; // @[issue-unit.scala 153:73]
  wire  slots_2_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_valid; // @[issue-unit.scala 153:73]
  wire [6:0] slots_2_io_in_uop_bits_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_2_io_in_uop_bits_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_2_io_in_uop_bits_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_2_io_in_uop_bits_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_2_io_in_uop_bits_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_2_io_in_uop_bits_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_2_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_2_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_2_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_2_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_2_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_in_uop_bits_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_is_br; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_2_io_in_uop_bits_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_2_io_in_uop_bits_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_2_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_in_uop_bits_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_2_io_in_uop_bits_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_2_io_in_uop_bits_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_in_uop_bits_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_2_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_2_io_in_uop_bits_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_in_uop_bits_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_in_uop_bits_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_in_uop_bits_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_in_uop_bits_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_2_io_in_uop_bits_ppred; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_2_io_in_uop_bits_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_2_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_in_uop_bits_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_in_uop_bits_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_in_uop_bits_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_in_uop_bits_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_in_uop_bits_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_2_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_2_io_out_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_2_io_out_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_2_io_out_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_2_io_out_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_2_io_out_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_2_io_out_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_2_io_out_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_2_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_2_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_2_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_2_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_out_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_2_io_out_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_2_io_out_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_2_io_out_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_out_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_2_io_out_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_2_io_out_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_out_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_2_io_out_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_2_io_out_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_out_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_out_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_out_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_out_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_out_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_2_io_out_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_out_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_2_io_out_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_2_io_out_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_out_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_out_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_out_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_out_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_out_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_out_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_out_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_out_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_2_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_out_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_out_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_2_io_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_2_io_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_2_io_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_2_io_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_2_io_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_2_io_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_2_io_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_2_io_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_2_io_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_2_io_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_2_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_2_io_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_2_io_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_2_io_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_2_io_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_2_io_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_2_io_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_2_io_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_2_io_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_2_io_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_2_io_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_2_io_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_2_io_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_2_io_debug_p1; // @[issue-unit.scala 153:73]
  wire  slots_2_io_debug_p2; // @[issue-unit.scala 153:73]
  wire  slots_2_io_debug_p3; // @[issue-unit.scala 153:73]
  wire  slots_2_io_debug_ppred; // @[issue-unit.scala 153:73]
  wire [1:0] slots_2_io_debug_state; // @[issue-unit.scala 153:73]
  wire  slots_3_clock; // @[issue-unit.scala 153:73]
  wire  slots_3_reset; // @[issue-unit.scala 153:73]
  wire  slots_3_io_valid; // @[issue-unit.scala 153:73]
  wire  slots_3_io_will_be_valid; // @[issue-unit.scala 153:73]
  wire  slots_3_io_request; // @[issue-unit.scala 153:73]
  wire  slots_3_io_request_hp; // @[issue-unit.scala 153:73]
  wire  slots_3_io_grant; // @[issue-unit.scala 153:73]
  wire [11:0] slots_3_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 153:73]
  wire [11:0] slots_3_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 153:73]
  wire [6:0] slots_3_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_3_io_brupdate_b2_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_3_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_3_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_3_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_3_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_3_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_3_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_3_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_3_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_3_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_3_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_3_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_3_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_3_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_3_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_3_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_3_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_3_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_3_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_3_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_valid; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_mispredict; // @[issue-unit.scala 153:73]
  wire  slots_3_io_brupdate_b2_taken; // @[issue-unit.scala 153:73]
  wire [2:0] slots_3_io_brupdate_b2_cfi_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_brupdate_b2_pc_sel; // @[issue-unit.scala 153:73]
  wire [39:0] slots_3_io_brupdate_b2_jalr_target; // @[issue-unit.scala 153:73]
  wire [20:0] slots_3_io_brupdate_b2_target_offset; // @[issue-unit.scala 153:73]
  wire  slots_3_io_kill; // @[issue-unit.scala 153:73]
  wire  slots_3_io_clear; // @[issue-unit.scala 153:73]
  wire  slots_3_io_ldspec_miss; // @[issue-unit.scala 153:73]
  wire  slots_3_io_wakeup_ports_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_3_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_3_io_wakeup_ports_1_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_3_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_3_io_wakeup_ports_2_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_3_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_3_io_wakeup_ports_3_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_3_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_3_io_wakeup_ports_4_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_3_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_3_io_pred_wakeup_port_valid; // @[issue-unit.scala 153:73]
  wire [4:0] slots_3_io_pred_wakeup_port_bits; // @[issue-unit.scala 153:73]
  wire  slots_3_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_valid; // @[issue-unit.scala 153:73]
  wire [6:0] slots_3_io_in_uop_bits_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_3_io_in_uop_bits_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_3_io_in_uop_bits_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_3_io_in_uop_bits_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_3_io_in_uop_bits_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_3_io_in_uop_bits_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_3_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_3_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_3_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_3_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_3_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_in_uop_bits_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_is_br; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_3_io_in_uop_bits_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_3_io_in_uop_bits_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_3_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_in_uop_bits_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_3_io_in_uop_bits_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_3_io_in_uop_bits_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_in_uop_bits_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_3_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_3_io_in_uop_bits_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_in_uop_bits_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_in_uop_bits_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_in_uop_bits_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_in_uop_bits_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_3_io_in_uop_bits_ppred; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_3_io_in_uop_bits_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_3_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_in_uop_bits_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_in_uop_bits_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_in_uop_bits_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_in_uop_bits_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_in_uop_bits_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_3_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_3_io_out_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_3_io_out_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_3_io_out_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_3_io_out_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_3_io_out_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_3_io_out_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_3_io_out_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_3_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_3_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_3_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_3_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_out_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_3_io_out_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_3_io_out_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_3_io_out_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_out_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_3_io_out_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_3_io_out_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_out_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_3_io_out_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_3_io_out_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_out_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_out_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_out_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_out_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_out_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_3_io_out_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_out_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_3_io_out_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_3_io_out_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_out_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_out_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_out_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_out_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_out_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_out_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_out_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_out_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_3_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_out_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_out_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_3_io_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_3_io_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_3_io_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_3_io_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_3_io_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_3_io_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_3_io_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_3_io_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_3_io_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_3_io_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_3_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_3_io_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_3_io_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_3_io_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_3_io_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_3_io_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_3_io_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_3_io_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_3_io_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_3_io_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_3_io_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_3_io_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_3_io_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_3_io_debug_p1; // @[issue-unit.scala 153:73]
  wire  slots_3_io_debug_p2; // @[issue-unit.scala 153:73]
  wire  slots_3_io_debug_p3; // @[issue-unit.scala 153:73]
  wire  slots_3_io_debug_ppred; // @[issue-unit.scala 153:73]
  wire [1:0] slots_3_io_debug_state; // @[issue-unit.scala 153:73]
  wire  slots_4_clock; // @[issue-unit.scala 153:73]
  wire  slots_4_reset; // @[issue-unit.scala 153:73]
  wire  slots_4_io_valid; // @[issue-unit.scala 153:73]
  wire  slots_4_io_will_be_valid; // @[issue-unit.scala 153:73]
  wire  slots_4_io_request; // @[issue-unit.scala 153:73]
  wire  slots_4_io_request_hp; // @[issue-unit.scala 153:73]
  wire  slots_4_io_grant; // @[issue-unit.scala 153:73]
  wire [11:0] slots_4_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 153:73]
  wire [11:0] slots_4_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 153:73]
  wire [6:0] slots_4_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_4_io_brupdate_b2_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_4_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_4_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_4_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_4_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_4_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_4_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_4_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_4_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_4_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_4_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_4_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_4_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_4_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_4_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_4_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_4_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_4_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_4_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_4_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_valid; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_mispredict; // @[issue-unit.scala 153:73]
  wire  slots_4_io_brupdate_b2_taken; // @[issue-unit.scala 153:73]
  wire [2:0] slots_4_io_brupdate_b2_cfi_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_brupdate_b2_pc_sel; // @[issue-unit.scala 153:73]
  wire [39:0] slots_4_io_brupdate_b2_jalr_target; // @[issue-unit.scala 153:73]
  wire [20:0] slots_4_io_brupdate_b2_target_offset; // @[issue-unit.scala 153:73]
  wire  slots_4_io_kill; // @[issue-unit.scala 153:73]
  wire  slots_4_io_clear; // @[issue-unit.scala 153:73]
  wire  slots_4_io_ldspec_miss; // @[issue-unit.scala 153:73]
  wire  slots_4_io_wakeup_ports_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_4_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_4_io_wakeup_ports_1_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_4_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_4_io_wakeup_ports_2_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_4_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_4_io_wakeup_ports_3_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_4_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_4_io_wakeup_ports_4_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_4_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_4_io_pred_wakeup_port_valid; // @[issue-unit.scala 153:73]
  wire [4:0] slots_4_io_pred_wakeup_port_bits; // @[issue-unit.scala 153:73]
  wire  slots_4_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_valid; // @[issue-unit.scala 153:73]
  wire [6:0] slots_4_io_in_uop_bits_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_4_io_in_uop_bits_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_4_io_in_uop_bits_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_4_io_in_uop_bits_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_4_io_in_uop_bits_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_4_io_in_uop_bits_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_4_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_4_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_4_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_4_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_4_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_in_uop_bits_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_is_br; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_4_io_in_uop_bits_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_4_io_in_uop_bits_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_4_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_in_uop_bits_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_4_io_in_uop_bits_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_4_io_in_uop_bits_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_in_uop_bits_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_4_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_4_io_in_uop_bits_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_in_uop_bits_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_in_uop_bits_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_in_uop_bits_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_in_uop_bits_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_4_io_in_uop_bits_ppred; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_4_io_in_uop_bits_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_4_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_in_uop_bits_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_in_uop_bits_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_in_uop_bits_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_in_uop_bits_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_in_uop_bits_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_4_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_4_io_out_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_4_io_out_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_4_io_out_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_4_io_out_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_4_io_out_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_4_io_out_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_4_io_out_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_4_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_4_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_4_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_4_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_out_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_4_io_out_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_4_io_out_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_4_io_out_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_out_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_4_io_out_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_4_io_out_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_out_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_4_io_out_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_4_io_out_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_out_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_out_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_out_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_out_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_out_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_4_io_out_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_out_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_4_io_out_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_4_io_out_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_out_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_out_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_out_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_out_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_out_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_out_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_out_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_out_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_4_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_out_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_out_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_4_io_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_4_io_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_4_io_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_4_io_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_4_io_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_4_io_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_4_io_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_4_io_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_4_io_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_4_io_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_4_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_4_io_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_4_io_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_4_io_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_4_io_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_4_io_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_4_io_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_4_io_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_4_io_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_4_io_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_4_io_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_4_io_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_4_io_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_4_io_debug_p1; // @[issue-unit.scala 153:73]
  wire  slots_4_io_debug_p2; // @[issue-unit.scala 153:73]
  wire  slots_4_io_debug_p3; // @[issue-unit.scala 153:73]
  wire  slots_4_io_debug_ppred; // @[issue-unit.scala 153:73]
  wire [1:0] slots_4_io_debug_state; // @[issue-unit.scala 153:73]
  wire  slots_5_clock; // @[issue-unit.scala 153:73]
  wire  slots_5_reset; // @[issue-unit.scala 153:73]
  wire  slots_5_io_valid; // @[issue-unit.scala 153:73]
  wire  slots_5_io_will_be_valid; // @[issue-unit.scala 153:73]
  wire  slots_5_io_request; // @[issue-unit.scala 153:73]
  wire  slots_5_io_request_hp; // @[issue-unit.scala 153:73]
  wire  slots_5_io_grant; // @[issue-unit.scala 153:73]
  wire [11:0] slots_5_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 153:73]
  wire [11:0] slots_5_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 153:73]
  wire [6:0] slots_5_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_5_io_brupdate_b2_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_5_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_5_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_5_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_5_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_5_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_5_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_5_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_5_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_5_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_5_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_5_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_5_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_5_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_5_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_5_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_5_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_5_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_5_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_5_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_valid; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_mispredict; // @[issue-unit.scala 153:73]
  wire  slots_5_io_brupdate_b2_taken; // @[issue-unit.scala 153:73]
  wire [2:0] slots_5_io_brupdate_b2_cfi_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_brupdate_b2_pc_sel; // @[issue-unit.scala 153:73]
  wire [39:0] slots_5_io_brupdate_b2_jalr_target; // @[issue-unit.scala 153:73]
  wire [20:0] slots_5_io_brupdate_b2_target_offset; // @[issue-unit.scala 153:73]
  wire  slots_5_io_kill; // @[issue-unit.scala 153:73]
  wire  slots_5_io_clear; // @[issue-unit.scala 153:73]
  wire  slots_5_io_ldspec_miss; // @[issue-unit.scala 153:73]
  wire  slots_5_io_wakeup_ports_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_5_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_5_io_wakeup_ports_1_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_5_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_5_io_wakeup_ports_2_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_5_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_5_io_wakeup_ports_3_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_5_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_5_io_wakeup_ports_4_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_5_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_5_io_pred_wakeup_port_valid; // @[issue-unit.scala 153:73]
  wire [4:0] slots_5_io_pred_wakeup_port_bits; // @[issue-unit.scala 153:73]
  wire  slots_5_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_valid; // @[issue-unit.scala 153:73]
  wire [6:0] slots_5_io_in_uop_bits_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_5_io_in_uop_bits_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_5_io_in_uop_bits_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_5_io_in_uop_bits_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_5_io_in_uop_bits_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_5_io_in_uop_bits_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_5_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_5_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_5_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_5_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_5_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_in_uop_bits_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_is_br; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_5_io_in_uop_bits_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_5_io_in_uop_bits_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_5_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_in_uop_bits_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_5_io_in_uop_bits_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_5_io_in_uop_bits_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_in_uop_bits_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_5_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_5_io_in_uop_bits_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_in_uop_bits_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_in_uop_bits_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_in_uop_bits_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_in_uop_bits_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_5_io_in_uop_bits_ppred; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_5_io_in_uop_bits_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_5_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_in_uop_bits_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_in_uop_bits_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_in_uop_bits_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_in_uop_bits_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_in_uop_bits_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_5_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_5_io_out_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_5_io_out_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_5_io_out_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_5_io_out_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_5_io_out_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_5_io_out_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_5_io_out_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_5_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_5_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_5_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_5_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_out_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_5_io_out_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_5_io_out_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_5_io_out_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_out_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_5_io_out_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_5_io_out_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_out_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_5_io_out_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_5_io_out_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_out_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_out_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_out_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_out_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_out_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_5_io_out_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_out_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_5_io_out_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_5_io_out_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_out_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_out_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_out_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_out_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_out_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_out_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_out_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_out_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_5_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_out_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_out_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_5_io_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_5_io_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_5_io_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_5_io_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_5_io_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_5_io_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_5_io_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_5_io_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_5_io_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_5_io_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_5_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_5_io_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_5_io_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_5_io_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_5_io_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_5_io_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_5_io_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_5_io_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_5_io_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_5_io_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_5_io_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_5_io_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_5_io_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_5_io_debug_p1; // @[issue-unit.scala 153:73]
  wire  slots_5_io_debug_p2; // @[issue-unit.scala 153:73]
  wire  slots_5_io_debug_p3; // @[issue-unit.scala 153:73]
  wire  slots_5_io_debug_ppred; // @[issue-unit.scala 153:73]
  wire [1:0] slots_5_io_debug_state; // @[issue-unit.scala 153:73]
  wire  slots_6_clock; // @[issue-unit.scala 153:73]
  wire  slots_6_reset; // @[issue-unit.scala 153:73]
  wire  slots_6_io_valid; // @[issue-unit.scala 153:73]
  wire  slots_6_io_will_be_valid; // @[issue-unit.scala 153:73]
  wire  slots_6_io_request; // @[issue-unit.scala 153:73]
  wire  slots_6_io_request_hp; // @[issue-unit.scala 153:73]
  wire  slots_6_io_grant; // @[issue-unit.scala 153:73]
  wire [11:0] slots_6_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 153:73]
  wire [11:0] slots_6_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 153:73]
  wire [6:0] slots_6_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_6_io_brupdate_b2_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_6_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_6_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_6_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_6_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_6_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_6_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_6_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_6_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_6_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_6_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_6_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_6_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_6_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_6_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_6_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_6_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_6_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_6_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_6_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_valid; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_mispredict; // @[issue-unit.scala 153:73]
  wire  slots_6_io_brupdate_b2_taken; // @[issue-unit.scala 153:73]
  wire [2:0] slots_6_io_brupdate_b2_cfi_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_brupdate_b2_pc_sel; // @[issue-unit.scala 153:73]
  wire [39:0] slots_6_io_brupdate_b2_jalr_target; // @[issue-unit.scala 153:73]
  wire [20:0] slots_6_io_brupdate_b2_target_offset; // @[issue-unit.scala 153:73]
  wire  slots_6_io_kill; // @[issue-unit.scala 153:73]
  wire  slots_6_io_clear; // @[issue-unit.scala 153:73]
  wire  slots_6_io_ldspec_miss; // @[issue-unit.scala 153:73]
  wire  slots_6_io_wakeup_ports_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_6_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_6_io_wakeup_ports_1_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_6_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_6_io_wakeup_ports_2_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_6_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_6_io_wakeup_ports_3_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_6_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_6_io_wakeup_ports_4_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_6_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_6_io_pred_wakeup_port_valid; // @[issue-unit.scala 153:73]
  wire [4:0] slots_6_io_pred_wakeup_port_bits; // @[issue-unit.scala 153:73]
  wire  slots_6_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_valid; // @[issue-unit.scala 153:73]
  wire [6:0] slots_6_io_in_uop_bits_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_6_io_in_uop_bits_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_6_io_in_uop_bits_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_6_io_in_uop_bits_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_6_io_in_uop_bits_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_6_io_in_uop_bits_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_6_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_6_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_6_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_6_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_6_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_in_uop_bits_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_is_br; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_6_io_in_uop_bits_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_6_io_in_uop_bits_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_6_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_in_uop_bits_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_6_io_in_uop_bits_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_6_io_in_uop_bits_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_in_uop_bits_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_6_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_6_io_in_uop_bits_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_in_uop_bits_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_in_uop_bits_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_in_uop_bits_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_in_uop_bits_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_6_io_in_uop_bits_ppred; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_6_io_in_uop_bits_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_6_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_in_uop_bits_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_in_uop_bits_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_in_uop_bits_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_in_uop_bits_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_in_uop_bits_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_6_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_6_io_out_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_6_io_out_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_6_io_out_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_6_io_out_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_6_io_out_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_6_io_out_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_6_io_out_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_6_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_6_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_6_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_6_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_out_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_6_io_out_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_6_io_out_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_6_io_out_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_out_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_6_io_out_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_6_io_out_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_out_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_6_io_out_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_6_io_out_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_out_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_out_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_out_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_out_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_out_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_6_io_out_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_out_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_6_io_out_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_6_io_out_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_out_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_out_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_out_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_out_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_out_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_out_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_out_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_out_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_6_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_out_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_out_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_6_io_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_6_io_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_6_io_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_6_io_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_6_io_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_6_io_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_6_io_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_6_io_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_6_io_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_6_io_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_6_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_6_io_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_6_io_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_6_io_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_6_io_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_6_io_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_6_io_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_6_io_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_6_io_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_6_io_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_6_io_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_6_io_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_6_io_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_6_io_debug_p1; // @[issue-unit.scala 153:73]
  wire  slots_6_io_debug_p2; // @[issue-unit.scala 153:73]
  wire  slots_6_io_debug_p3; // @[issue-unit.scala 153:73]
  wire  slots_6_io_debug_ppred; // @[issue-unit.scala 153:73]
  wire [1:0] slots_6_io_debug_state; // @[issue-unit.scala 153:73]
  wire  slots_7_clock; // @[issue-unit.scala 153:73]
  wire  slots_7_reset; // @[issue-unit.scala 153:73]
  wire  slots_7_io_valid; // @[issue-unit.scala 153:73]
  wire  slots_7_io_will_be_valid; // @[issue-unit.scala 153:73]
  wire  slots_7_io_request; // @[issue-unit.scala 153:73]
  wire  slots_7_io_request_hp; // @[issue-unit.scala 153:73]
  wire  slots_7_io_grant; // @[issue-unit.scala 153:73]
  wire [11:0] slots_7_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 153:73]
  wire [11:0] slots_7_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 153:73]
  wire [6:0] slots_7_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_7_io_brupdate_b2_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_7_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_7_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_7_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_7_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_7_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_7_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_7_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_7_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_7_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_7_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_7_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_7_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_7_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_7_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_7_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_7_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_7_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_7_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_7_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_valid; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_mispredict; // @[issue-unit.scala 153:73]
  wire  slots_7_io_brupdate_b2_taken; // @[issue-unit.scala 153:73]
  wire [2:0] slots_7_io_brupdate_b2_cfi_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_brupdate_b2_pc_sel; // @[issue-unit.scala 153:73]
  wire [39:0] slots_7_io_brupdate_b2_jalr_target; // @[issue-unit.scala 153:73]
  wire [20:0] slots_7_io_brupdate_b2_target_offset; // @[issue-unit.scala 153:73]
  wire  slots_7_io_kill; // @[issue-unit.scala 153:73]
  wire  slots_7_io_clear; // @[issue-unit.scala 153:73]
  wire  slots_7_io_ldspec_miss; // @[issue-unit.scala 153:73]
  wire  slots_7_io_wakeup_ports_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_7_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_7_io_wakeup_ports_1_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_7_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_7_io_wakeup_ports_2_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_7_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_7_io_wakeup_ports_3_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_7_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_7_io_wakeup_ports_4_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_7_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_7_io_pred_wakeup_port_valid; // @[issue-unit.scala 153:73]
  wire [4:0] slots_7_io_pred_wakeup_port_bits; // @[issue-unit.scala 153:73]
  wire  slots_7_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_valid; // @[issue-unit.scala 153:73]
  wire [6:0] slots_7_io_in_uop_bits_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_7_io_in_uop_bits_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_7_io_in_uop_bits_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_7_io_in_uop_bits_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_7_io_in_uop_bits_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_7_io_in_uop_bits_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_7_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_7_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_7_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_7_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_7_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_in_uop_bits_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_is_br; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_7_io_in_uop_bits_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_7_io_in_uop_bits_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_7_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_in_uop_bits_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_7_io_in_uop_bits_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_7_io_in_uop_bits_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_in_uop_bits_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_7_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_7_io_in_uop_bits_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_in_uop_bits_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_in_uop_bits_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_in_uop_bits_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_in_uop_bits_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_7_io_in_uop_bits_ppred; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_7_io_in_uop_bits_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_7_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_in_uop_bits_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_in_uop_bits_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_in_uop_bits_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_in_uop_bits_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_in_uop_bits_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_7_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_7_io_out_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_7_io_out_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_7_io_out_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_7_io_out_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_7_io_out_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_7_io_out_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_7_io_out_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_7_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_7_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_7_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_7_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_out_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_7_io_out_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_7_io_out_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_7_io_out_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_out_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_7_io_out_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_7_io_out_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_out_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_7_io_out_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_7_io_out_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_out_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_out_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_out_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_out_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_out_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_7_io_out_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_out_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_7_io_out_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_7_io_out_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_out_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_out_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_out_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_out_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_out_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_out_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_out_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_out_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_7_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_out_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_out_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_7_io_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_7_io_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_7_io_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_7_io_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_7_io_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_7_io_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_7_io_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_7_io_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_7_io_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_7_io_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_7_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_7_io_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_7_io_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_7_io_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_7_io_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_7_io_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_7_io_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_7_io_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_7_io_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_7_io_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_7_io_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_7_io_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_7_io_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_7_io_debug_p1; // @[issue-unit.scala 153:73]
  wire  slots_7_io_debug_p2; // @[issue-unit.scala 153:73]
  wire  slots_7_io_debug_p3; // @[issue-unit.scala 153:73]
  wire  slots_7_io_debug_ppred; // @[issue-unit.scala 153:73]
  wire [1:0] slots_7_io_debug_state; // @[issue-unit.scala 153:73]
  wire  slots_8_clock; // @[issue-unit.scala 153:73]
  wire  slots_8_reset; // @[issue-unit.scala 153:73]
  wire  slots_8_io_valid; // @[issue-unit.scala 153:73]
  wire  slots_8_io_will_be_valid; // @[issue-unit.scala 153:73]
  wire  slots_8_io_request; // @[issue-unit.scala 153:73]
  wire  slots_8_io_request_hp; // @[issue-unit.scala 153:73]
  wire  slots_8_io_grant; // @[issue-unit.scala 153:73]
  wire [11:0] slots_8_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 153:73]
  wire [11:0] slots_8_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 153:73]
  wire [6:0] slots_8_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_8_io_brupdate_b2_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_8_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_8_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_8_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_8_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_8_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_8_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_8_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_8_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_8_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_8_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_8_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_8_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_8_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_8_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_8_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_8_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_8_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_8_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_8_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_valid; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_mispredict; // @[issue-unit.scala 153:73]
  wire  slots_8_io_brupdate_b2_taken; // @[issue-unit.scala 153:73]
  wire [2:0] slots_8_io_brupdate_b2_cfi_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_brupdate_b2_pc_sel; // @[issue-unit.scala 153:73]
  wire [39:0] slots_8_io_brupdate_b2_jalr_target; // @[issue-unit.scala 153:73]
  wire [20:0] slots_8_io_brupdate_b2_target_offset; // @[issue-unit.scala 153:73]
  wire  slots_8_io_kill; // @[issue-unit.scala 153:73]
  wire  slots_8_io_clear; // @[issue-unit.scala 153:73]
  wire  slots_8_io_ldspec_miss; // @[issue-unit.scala 153:73]
  wire  slots_8_io_wakeup_ports_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_8_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_8_io_wakeup_ports_1_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_8_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_8_io_wakeup_ports_2_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_8_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_8_io_wakeup_ports_3_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_8_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_8_io_wakeup_ports_4_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_8_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_8_io_pred_wakeup_port_valid; // @[issue-unit.scala 153:73]
  wire [4:0] slots_8_io_pred_wakeup_port_bits; // @[issue-unit.scala 153:73]
  wire  slots_8_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_valid; // @[issue-unit.scala 153:73]
  wire [6:0] slots_8_io_in_uop_bits_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_8_io_in_uop_bits_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_8_io_in_uop_bits_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_8_io_in_uop_bits_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_8_io_in_uop_bits_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_8_io_in_uop_bits_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_8_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_8_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_8_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_8_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_8_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_in_uop_bits_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_is_br; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_8_io_in_uop_bits_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_8_io_in_uop_bits_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_8_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_in_uop_bits_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_8_io_in_uop_bits_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_8_io_in_uop_bits_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_in_uop_bits_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_8_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_8_io_in_uop_bits_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_in_uop_bits_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_in_uop_bits_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_in_uop_bits_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_in_uop_bits_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_8_io_in_uop_bits_ppred; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_8_io_in_uop_bits_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_8_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_in_uop_bits_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_in_uop_bits_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_in_uop_bits_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_in_uop_bits_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_in_uop_bits_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_8_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_8_io_out_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_8_io_out_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_8_io_out_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_8_io_out_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_8_io_out_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_8_io_out_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_8_io_out_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_8_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_8_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_8_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_8_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_out_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_8_io_out_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_8_io_out_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_8_io_out_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_out_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_8_io_out_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_8_io_out_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_out_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_8_io_out_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_8_io_out_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_out_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_out_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_out_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_out_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_out_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_8_io_out_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_out_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_8_io_out_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_8_io_out_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_out_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_out_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_out_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_out_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_out_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_out_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_out_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_out_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_8_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_out_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_out_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_8_io_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_8_io_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_8_io_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_8_io_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_8_io_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_8_io_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_8_io_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_8_io_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_8_io_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_8_io_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_8_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_8_io_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_8_io_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_8_io_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_8_io_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_8_io_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_8_io_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_8_io_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_8_io_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_8_io_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_8_io_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_8_io_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_8_io_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_8_io_debug_p1; // @[issue-unit.scala 153:73]
  wire  slots_8_io_debug_p2; // @[issue-unit.scala 153:73]
  wire  slots_8_io_debug_p3; // @[issue-unit.scala 153:73]
  wire  slots_8_io_debug_ppred; // @[issue-unit.scala 153:73]
  wire [1:0] slots_8_io_debug_state; // @[issue-unit.scala 153:73]
  wire  slots_9_clock; // @[issue-unit.scala 153:73]
  wire  slots_9_reset; // @[issue-unit.scala 153:73]
  wire  slots_9_io_valid; // @[issue-unit.scala 153:73]
  wire  slots_9_io_will_be_valid; // @[issue-unit.scala 153:73]
  wire  slots_9_io_request; // @[issue-unit.scala 153:73]
  wire  slots_9_io_request_hp; // @[issue-unit.scala 153:73]
  wire  slots_9_io_grant; // @[issue-unit.scala 153:73]
  wire [11:0] slots_9_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 153:73]
  wire [11:0] slots_9_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 153:73]
  wire [6:0] slots_9_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_9_io_brupdate_b2_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_9_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_9_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_9_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_9_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_9_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_9_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_9_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_9_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_9_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_9_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_9_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_9_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_9_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_9_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_9_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_9_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_9_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_9_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_9_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_valid; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_mispredict; // @[issue-unit.scala 153:73]
  wire  slots_9_io_brupdate_b2_taken; // @[issue-unit.scala 153:73]
  wire [2:0] slots_9_io_brupdate_b2_cfi_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_brupdate_b2_pc_sel; // @[issue-unit.scala 153:73]
  wire [39:0] slots_9_io_brupdate_b2_jalr_target; // @[issue-unit.scala 153:73]
  wire [20:0] slots_9_io_brupdate_b2_target_offset; // @[issue-unit.scala 153:73]
  wire  slots_9_io_kill; // @[issue-unit.scala 153:73]
  wire  slots_9_io_clear; // @[issue-unit.scala 153:73]
  wire  slots_9_io_ldspec_miss; // @[issue-unit.scala 153:73]
  wire  slots_9_io_wakeup_ports_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_9_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_9_io_wakeup_ports_1_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_9_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_9_io_wakeup_ports_2_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_9_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_9_io_wakeup_ports_3_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_9_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_9_io_wakeup_ports_4_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_9_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_9_io_pred_wakeup_port_valid; // @[issue-unit.scala 153:73]
  wire [4:0] slots_9_io_pred_wakeup_port_bits; // @[issue-unit.scala 153:73]
  wire  slots_9_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_valid; // @[issue-unit.scala 153:73]
  wire [6:0] slots_9_io_in_uop_bits_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_9_io_in_uop_bits_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_9_io_in_uop_bits_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_9_io_in_uop_bits_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_9_io_in_uop_bits_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_9_io_in_uop_bits_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_9_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_9_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_9_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_9_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_9_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_in_uop_bits_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_is_br; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_9_io_in_uop_bits_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_9_io_in_uop_bits_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_9_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_in_uop_bits_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_9_io_in_uop_bits_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_9_io_in_uop_bits_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_in_uop_bits_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_9_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_9_io_in_uop_bits_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_in_uop_bits_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_in_uop_bits_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_in_uop_bits_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_in_uop_bits_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_9_io_in_uop_bits_ppred; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_9_io_in_uop_bits_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_9_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_in_uop_bits_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_in_uop_bits_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_in_uop_bits_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_in_uop_bits_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_in_uop_bits_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_9_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_9_io_out_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_9_io_out_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_9_io_out_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_9_io_out_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_9_io_out_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_9_io_out_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_9_io_out_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_9_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_9_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_9_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_9_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_out_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_9_io_out_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_9_io_out_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_9_io_out_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_out_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_9_io_out_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_9_io_out_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_out_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_9_io_out_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_9_io_out_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_out_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_out_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_out_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_out_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_out_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_9_io_out_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_out_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_9_io_out_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_9_io_out_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_out_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_out_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_out_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_out_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_out_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_out_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_out_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_out_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_9_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_out_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_out_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_9_io_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_9_io_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_9_io_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_9_io_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_9_io_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_9_io_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_9_io_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_9_io_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_9_io_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_9_io_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_9_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_9_io_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_9_io_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_9_io_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_9_io_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_9_io_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_9_io_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_9_io_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_9_io_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_9_io_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_9_io_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_9_io_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_9_io_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_9_io_debug_p1; // @[issue-unit.scala 153:73]
  wire  slots_9_io_debug_p2; // @[issue-unit.scala 153:73]
  wire  slots_9_io_debug_p3; // @[issue-unit.scala 153:73]
  wire  slots_9_io_debug_ppred; // @[issue-unit.scala 153:73]
  wire [1:0] slots_9_io_debug_state; // @[issue-unit.scala 153:73]
  wire  slots_10_clock; // @[issue-unit.scala 153:73]
  wire  slots_10_reset; // @[issue-unit.scala 153:73]
  wire  slots_10_io_valid; // @[issue-unit.scala 153:73]
  wire  slots_10_io_will_be_valid; // @[issue-unit.scala 153:73]
  wire  slots_10_io_request; // @[issue-unit.scala 153:73]
  wire  slots_10_io_request_hp; // @[issue-unit.scala 153:73]
  wire  slots_10_io_grant; // @[issue-unit.scala 153:73]
  wire [11:0] slots_10_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 153:73]
  wire [11:0] slots_10_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 153:73]
  wire [6:0] slots_10_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_10_io_brupdate_b2_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_10_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_10_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_10_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_10_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_10_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_10_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_10_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_10_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_10_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_10_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_10_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_10_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_10_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_10_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_10_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_10_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_10_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_10_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_10_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_valid; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_mispredict; // @[issue-unit.scala 153:73]
  wire  slots_10_io_brupdate_b2_taken; // @[issue-unit.scala 153:73]
  wire [2:0] slots_10_io_brupdate_b2_cfi_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_brupdate_b2_pc_sel; // @[issue-unit.scala 153:73]
  wire [39:0] slots_10_io_brupdate_b2_jalr_target; // @[issue-unit.scala 153:73]
  wire [20:0] slots_10_io_brupdate_b2_target_offset; // @[issue-unit.scala 153:73]
  wire  slots_10_io_kill; // @[issue-unit.scala 153:73]
  wire  slots_10_io_clear; // @[issue-unit.scala 153:73]
  wire  slots_10_io_ldspec_miss; // @[issue-unit.scala 153:73]
  wire  slots_10_io_wakeup_ports_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_10_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_10_io_wakeup_ports_1_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_10_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_10_io_wakeup_ports_2_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_10_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_10_io_wakeup_ports_3_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_10_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_10_io_wakeup_ports_4_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_10_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_10_io_pred_wakeup_port_valid; // @[issue-unit.scala 153:73]
  wire [4:0] slots_10_io_pred_wakeup_port_bits; // @[issue-unit.scala 153:73]
  wire  slots_10_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_valid; // @[issue-unit.scala 153:73]
  wire [6:0] slots_10_io_in_uop_bits_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_10_io_in_uop_bits_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_10_io_in_uop_bits_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_10_io_in_uop_bits_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_10_io_in_uop_bits_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_10_io_in_uop_bits_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_10_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_10_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_10_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_10_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_10_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_in_uop_bits_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_is_br; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_10_io_in_uop_bits_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_10_io_in_uop_bits_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_10_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_in_uop_bits_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_10_io_in_uop_bits_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_10_io_in_uop_bits_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_in_uop_bits_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_10_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_10_io_in_uop_bits_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_in_uop_bits_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_in_uop_bits_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_in_uop_bits_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_in_uop_bits_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_10_io_in_uop_bits_ppred; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_10_io_in_uop_bits_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_10_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_in_uop_bits_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_in_uop_bits_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_in_uop_bits_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_in_uop_bits_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_in_uop_bits_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_10_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_10_io_out_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_10_io_out_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_10_io_out_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_10_io_out_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_10_io_out_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_10_io_out_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_10_io_out_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_10_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_10_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_10_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_10_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_out_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_10_io_out_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_10_io_out_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_10_io_out_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_out_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_10_io_out_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_10_io_out_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_out_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_10_io_out_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_10_io_out_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_out_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_out_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_out_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_out_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_out_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_10_io_out_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_out_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_10_io_out_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_10_io_out_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_out_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_out_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_out_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_out_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_out_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_out_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_out_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_out_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_10_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_out_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_out_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_10_io_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_10_io_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_10_io_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_10_io_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_10_io_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_10_io_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_10_io_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_10_io_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_10_io_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_10_io_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_10_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_10_io_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_10_io_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_10_io_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_10_io_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_10_io_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_10_io_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_10_io_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_10_io_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_10_io_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_10_io_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_10_io_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_10_io_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_10_io_debug_p1; // @[issue-unit.scala 153:73]
  wire  slots_10_io_debug_p2; // @[issue-unit.scala 153:73]
  wire  slots_10_io_debug_p3; // @[issue-unit.scala 153:73]
  wire  slots_10_io_debug_ppred; // @[issue-unit.scala 153:73]
  wire [1:0] slots_10_io_debug_state; // @[issue-unit.scala 153:73]
  wire  slots_11_clock; // @[issue-unit.scala 153:73]
  wire  slots_11_reset; // @[issue-unit.scala 153:73]
  wire  slots_11_io_valid; // @[issue-unit.scala 153:73]
  wire  slots_11_io_will_be_valid; // @[issue-unit.scala 153:73]
  wire  slots_11_io_request; // @[issue-unit.scala 153:73]
  wire  slots_11_io_request_hp; // @[issue-unit.scala 153:73]
  wire  slots_11_io_grant; // @[issue-unit.scala 153:73]
  wire [11:0] slots_11_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 153:73]
  wire [11:0] slots_11_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 153:73]
  wire [6:0] slots_11_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_11_io_brupdate_b2_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_11_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_11_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_11_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_11_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_11_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_11_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_11_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_11_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_11_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_11_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_11_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_11_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_11_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_11_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_11_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_11_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_11_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_11_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_11_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_valid; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_mispredict; // @[issue-unit.scala 153:73]
  wire  slots_11_io_brupdate_b2_taken; // @[issue-unit.scala 153:73]
  wire [2:0] slots_11_io_brupdate_b2_cfi_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_brupdate_b2_pc_sel; // @[issue-unit.scala 153:73]
  wire [39:0] slots_11_io_brupdate_b2_jalr_target; // @[issue-unit.scala 153:73]
  wire [20:0] slots_11_io_brupdate_b2_target_offset; // @[issue-unit.scala 153:73]
  wire  slots_11_io_kill; // @[issue-unit.scala 153:73]
  wire  slots_11_io_clear; // @[issue-unit.scala 153:73]
  wire  slots_11_io_ldspec_miss; // @[issue-unit.scala 153:73]
  wire  slots_11_io_wakeup_ports_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_11_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_11_io_wakeup_ports_1_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_11_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_11_io_wakeup_ports_2_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_11_io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_11_io_wakeup_ports_3_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_11_io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_11_io_wakeup_ports_4_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 153:73]
  wire  slots_11_io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_11_io_pred_wakeup_port_valid; // @[issue-unit.scala 153:73]
  wire [4:0] slots_11_io_pred_wakeup_port_bits; // @[issue-unit.scala 153:73]
  wire  slots_11_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_valid; // @[issue-unit.scala 153:73]
  wire [6:0] slots_11_io_in_uop_bits_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_11_io_in_uop_bits_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_11_io_in_uop_bits_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_11_io_in_uop_bits_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_11_io_in_uop_bits_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_11_io_in_uop_bits_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_11_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_11_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_11_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_11_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_11_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_in_uop_bits_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_is_br; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_11_io_in_uop_bits_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_11_io_in_uop_bits_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_11_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_in_uop_bits_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_11_io_in_uop_bits_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_11_io_in_uop_bits_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_in_uop_bits_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_11_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_11_io_in_uop_bits_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_in_uop_bits_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_in_uop_bits_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_in_uop_bits_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_in_uop_bits_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_11_io_in_uop_bits_ppred; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_11_io_in_uop_bits_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_11_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_in_uop_bits_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_in_uop_bits_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_in_uop_bits_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_in_uop_bits_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_in_uop_bits_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_11_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_11_io_out_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_11_io_out_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_11_io_out_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_11_io_out_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_11_io_out_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_11_io_out_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_11_io_out_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_11_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_11_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_11_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_11_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_out_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_11_io_out_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_11_io_out_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_11_io_out_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_out_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_11_io_out_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_11_io_out_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_out_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_11_io_out_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_11_io_out_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_out_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_out_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_out_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_out_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_out_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_11_io_out_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_out_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_11_io_out_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_11_io_out_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_out_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_out_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_out_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_out_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_out_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_out_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_out_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_out_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_11_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_out_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_out_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire [6:0] slots_11_io_uop_uopc; // @[issue-unit.scala 153:73]
  wire [31:0] slots_11_io_uop_inst; // @[issue-unit.scala 153:73]
  wire [31:0] slots_11_io_uop_debug_inst; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_is_rvc; // @[issue-unit.scala 153:73]
  wire [39:0] slots_11_io_uop_debug_pc; // @[issue-unit.scala 153:73]
  wire [2:0] slots_11_io_uop_iq_type; // @[issue-unit.scala 153:73]
  wire [9:0] slots_11_io_uop_fu_code; // @[issue-unit.scala 153:73]
  wire [3:0] slots_11_io_uop_ctrl_br_type; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_uop_ctrl_op1_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_11_io_uop_ctrl_op2_sel; // @[issue-unit.scala 153:73]
  wire [2:0] slots_11_io_uop_ctrl_imm_sel; // @[issue-unit.scala 153:73]
  wire [3:0] slots_11_io_uop_ctrl_op_fcn; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 153:73]
  wire [2:0] slots_11_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_ctrl_is_load; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_ctrl_is_sta; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_ctrl_is_std; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_uop_iw_state; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_iw_p1_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_iw_p2_poisoned; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_is_br; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_is_jalr; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_is_jal; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_is_sfb; // @[issue-unit.scala 153:73]
  wire [11:0] slots_11_io_uop_br_mask; // @[issue-unit.scala 153:73]
  wire [3:0] slots_11_io_uop_br_tag; // @[issue-unit.scala 153:73]
  wire [4:0] slots_11_io_uop_ftq_idx; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_edge_inst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_uop_pc_lob; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_taken; // @[issue-unit.scala 153:73]
  wire [19:0] slots_11_io_uop_imm_packed; // @[issue-unit.scala 153:73]
  wire [11:0] slots_11_io_uop_csr_addr; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_uop_rob_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_11_io_uop_ldq_idx; // @[issue-unit.scala 153:73]
  wire [3:0] slots_11_io_uop_stq_idx; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_uop_rxq_idx; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_uop_pdst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_uop_prs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_uop_prs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_uop_prs3; // @[issue-unit.scala 153:73]
  wire [4:0] slots_11_io_uop_ppred; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_prs1_busy; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_prs2_busy; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_prs3_busy; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_ppred_busy; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_uop_stale_pdst; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_exception; // @[issue-unit.scala 153:73]
  wire [63:0] slots_11_io_uop_exc_cause; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_bypassable; // @[issue-unit.scala 153:73]
  wire [4:0] slots_11_io_uop_mem_cmd; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_uop_mem_size; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_mem_signed; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_is_fence; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_is_fencei; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_is_amo; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_uses_ldq; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_uses_stq; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_is_sys_pc2epc; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_is_unique; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_flush_on_commit; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_ldst_is_rs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_uop_ldst; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_uop_lrs1; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_uop_lrs2; // @[issue-unit.scala 153:73]
  wire [5:0] slots_11_io_uop_lrs3; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_ldst_val; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_uop_dst_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_uop_lrs1_rtype; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_uop_lrs2_rtype; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_frs3_en; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_fp_val; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_fp_single; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_xcpt_pf_if; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_xcpt_ae_if; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_xcpt_ma_if; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_bp_debug_if; // @[issue-unit.scala 153:73]
  wire  slots_11_io_uop_bp_xcpt_if; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_uop_debug_fsrc; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_uop_debug_tsrc; // @[issue-unit.scala 153:73]
  wire  slots_11_io_debug_p1; // @[issue-unit.scala 153:73]
  wire  slots_11_io_debug_p2; // @[issue-unit.scala 153:73]
  wire  slots_11_io_debug_p3; // @[issue-unit.scala 153:73]
  wire  slots_11_io_debug_ppred; // @[issue-unit.scala 153:73]
  wire [1:0] slots_11_io_debug_state; // @[issue-unit.scala 153:73]
  wire  _T = io_dis_uops_0_bits_uopc == 7'h2; // @[issue-unit.scala 127:39]
  wire  _T_3 = io_dis_uops_0_bits_uopc == 7'h43; // @[issue-unit.scala 128:39]
  wire  _T_4 = io_dis_uops_0_bits_uopc == 7'h2 & io_dis_uops_0_bits_lrs2_rtype == 2'h0 | _T_3; // @[issue-unit.scala 127:96]
  wire [1:0] _GEN_0 = _T & io_dis_uops_0_bits_lrs2_rtype != 2'h0 ? 2'h2 : io_dis_uops_0_bits_lrs2_rtype; // @[issue-unit.scala 131:102 issue-unit.scala 132:32 issue-unit.scala 120:17]
  wire  _GEN_1 = _T & io_dis_uops_0_bits_lrs2_rtype != 2'h0 ? 1'h0 : io_dis_uops_0_bits_prs2_busy; // @[issue-unit.scala 131:102 issue-unit.scala 133:32 issue-unit.scala 120:17]
  wire [1:0] uops_12_iw_state = _T_4 ? 2'h2 : 2'h1; // @[issue-unit.scala 128:54 issue-unit.scala 129:30 issue-unit.scala 123:26]
  wire [1:0] uops_12_lrs2_rtype = _T_4 ? io_dis_uops_0_bits_lrs2_rtype : _GEN_0; // @[issue-unit.scala 128:54 issue-unit.scala 120:17]
  wire  uops_12_prs2_busy = _T_4 ? io_dis_uops_0_bits_prs2_busy : _GEN_1; // @[issue-unit.scala 128:54 issue-unit.scala 120:17]
  wire  _T_13 = io_dis_uops_1_bits_uopc == 7'h2; // @[issue-unit.scala 127:39]
  wire  _T_16 = io_dis_uops_1_bits_uopc == 7'h43; // @[issue-unit.scala 128:39]
  wire  _T_17 = io_dis_uops_1_bits_uopc == 7'h2 & io_dis_uops_1_bits_lrs2_rtype == 2'h0 | _T_16; // @[issue-unit.scala 127:96]
  wire [1:0] _GEN_5 = _T_13 & io_dis_uops_1_bits_lrs2_rtype != 2'h0 ? 2'h2 : io_dis_uops_1_bits_lrs2_rtype; // @[issue-unit.scala 131:102 issue-unit.scala 132:32 issue-unit.scala 120:17]
  wire  _GEN_6 = _T_13 & io_dis_uops_1_bits_lrs2_rtype != 2'h0 ? 1'h0 : io_dis_uops_1_bits_prs2_busy; // @[issue-unit.scala 131:102 issue-unit.scala 133:32 issue-unit.scala 120:17]
  wire [1:0] uops_13_iw_state = _T_17 ? 2'h2 : 2'h1; // @[issue-unit.scala 128:54 issue-unit.scala 129:30 issue-unit.scala 123:26]
  wire [1:0] uops_13_lrs2_rtype = _T_17 ? io_dis_uops_1_bits_lrs2_rtype : _GEN_5; // @[issue-unit.scala 128:54 issue-unit.scala 120:17]
  wire  uops_13_prs2_busy = _T_17 ? io_dis_uops_1_bits_prs2_busy : _GEN_6; // @[issue-unit.scala 128:54 issue-unit.scala 120:17]
  wire  issue_slots_0_valid = slots_0_io_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_valid = slots_1_io_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_valid = slots_2_io_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_valid = slots_3_io_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_valid = slots_4_io_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_valid = slots_5_io_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_valid = slots_6_io_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_valid = slots_7_io_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_valid = slots_8_io_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_valid = slots_9_io_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_valid = slots_10_io_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_valid = slots_11_io_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_request = slots_1_io_request; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_1_uop_fu_code = slots_1_io_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] _T_285 = issue_slots_1_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 116:54]
  wire  _T_286 = _T_285 != 10'h0; // @[issue-unit-age-ordered.scala 116:72]
  wire  _T_289 = issue_slots_1_request & _T_286; // @[issue-unit-age-ordered.scala 118:40]
  wire  issue_slots_0_request = slots_0_io_request; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_0_uop_fu_code = slots_0_io_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] _T_270 = issue_slots_0_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 116:54]
  wire  _T_271 = _T_270 != 10'h0; // @[issue-unit-age-ordered.scala 116:72]
  wire  _T_279 = issue_slots_0_request & _T_271; // @[issue-unit-age-ordered.scala 124:52]
  wire  issue_slots_1_grant = issue_slots_1_request & _T_286 & ~_T_279; // @[issue-unit-age-ordered.scala 118:56]
  wire  issue_slots_2_request = slots_2_io_request; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_2_uop_fu_code = slots_2_io_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] _T_300 = issue_slots_2_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 116:54]
  wire  _T_301 = _T_300 != 10'h0; // @[issue-unit-age-ordered.scala 116:72]
  wire  _T_304 = issue_slots_2_request & _T_301; // @[issue-unit-age-ordered.scala 118:40]
  wire  _T_295 = _T_289 | issue_slots_0_request & _T_271; // @[issue-unit-age-ordered.scala 124:69]
  wire  issue_slots_2_grant = issue_slots_2_request & _T_301 & ~_T_295; // @[issue-unit-age-ordered.scala 118:56]
  wire [1:0] _T_59 = issue_slots_1_grant + issue_slots_2_grant; // @[Bitwise.scala 47:55]
  wire [1:0] _GEN_2931 = {{1'd0}, _T_279}; // @[Bitwise.scala 47:55]
  wire [2:0] _T_61 = _GEN_2931 + _T_59; // @[Bitwise.scala 47:55]
  wire  issue_slots_4_request = slots_4_io_request; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_4_uop_fu_code = slots_4_io_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] _T_330 = issue_slots_4_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 116:54]
  wire  _T_331 = _T_330 != 10'h0; // @[issue-unit-age-ordered.scala 116:72]
  wire  _T_334 = issue_slots_4_request & _T_331; // @[issue-unit-age-ordered.scala 118:40]
  wire  issue_slots_3_request = slots_3_io_request; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_3_uop_fu_code = slots_3_io_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] _T_315 = issue_slots_3_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 116:54]
  wire  _T_316 = _T_315 != 10'h0; // @[issue-unit-age-ordered.scala 116:72]
  wire  _T_324 = issue_slots_3_request & _T_316; // @[issue-unit-age-ordered.scala 124:52]
  wire  _T_310 = _T_304 | (_T_289 | issue_slots_0_request & _T_271); // @[issue-unit-age-ordered.scala 124:69]
  wire  _T_325 = issue_slots_3_request & _T_316 | (_T_304 | (_T_289 | issue_slots_0_request & _T_271)); // @[issue-unit-age-ordered.scala 124:69]
  wire  issue_slots_4_grant = issue_slots_4_request & _T_331 & ~_T_325; // @[issue-unit-age-ordered.scala 118:56]
  wire  issue_slots_5_request = slots_5_io_request; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_5_uop_fu_code = slots_5_io_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] _T_345 = issue_slots_5_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 116:54]
  wire  _T_346 = _T_345 != 10'h0; // @[issue-unit-age-ordered.scala 116:72]
  wire  _T_349 = issue_slots_5_request & _T_346; // @[issue-unit-age-ordered.scala 118:40]
  wire  _T_340 = _T_334 | (issue_slots_3_request & _T_316 | (_T_304 | (_T_289 | issue_slots_0_request & _T_271))); // @[issue-unit-age-ordered.scala 124:69]
  wire  issue_slots_5_grant = issue_slots_5_request & _T_346 & ~_T_340; // @[issue-unit-age-ordered.scala 118:56]
  wire [1:0] _T_63 = issue_slots_4_grant + issue_slots_5_grant; // @[Bitwise.scala 47:55]
  wire  issue_slots_3_grant = _T_324 & ~_T_310; // @[issue-unit-age-ordered.scala 118:56]
  wire [1:0] _GEN_2932 = {{1'd0}, issue_slots_3_grant}; // @[Bitwise.scala 47:55]
  wire [2:0] _T_65 = _GEN_2932 + _T_63; // @[Bitwise.scala 47:55]
  wire [2:0] _T_67 = _T_61[1:0] + _T_65[1:0]; // @[Bitwise.scala 47:55]
  wire  issue_slots_7_request = slots_7_io_request; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_7_uop_fu_code = slots_7_io_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] _T_375 = issue_slots_7_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 116:54]
  wire  _T_376 = _T_375 != 10'h0; // @[issue-unit-age-ordered.scala 116:72]
  wire  _T_379 = issue_slots_7_request & _T_376; // @[issue-unit-age-ordered.scala 118:40]
  wire  issue_slots_6_request = slots_6_io_request; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_6_uop_fu_code = slots_6_io_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] _T_360 = issue_slots_6_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 116:54]
  wire  _T_361 = _T_360 != 10'h0; // @[issue-unit-age-ordered.scala 116:72]
  wire  _T_369 = issue_slots_6_request & _T_361; // @[issue-unit-age-ordered.scala 124:52]
  wire  _T_355 = _T_349 | (_T_334 | (issue_slots_3_request & _T_316 | (_T_304 | (_T_289 | issue_slots_0_request & _T_271
    )))); // @[issue-unit-age-ordered.scala 124:69]
  wire  _T_370 = issue_slots_6_request & _T_361 | (_T_349 | (_T_334 | (issue_slots_3_request & _T_316 | (_T_304 | (
    _T_289 | issue_slots_0_request & _T_271))))); // @[issue-unit-age-ordered.scala 124:69]
  wire  issue_slots_7_grant = issue_slots_7_request & _T_376 & ~_T_370; // @[issue-unit-age-ordered.scala 118:56]
  wire  issue_slots_8_request = slots_8_io_request; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_8_uop_fu_code = slots_8_io_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] _T_390 = issue_slots_8_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 116:54]
  wire  _T_391 = _T_390 != 10'h0; // @[issue-unit-age-ordered.scala 116:72]
  wire  _T_394 = issue_slots_8_request & _T_391; // @[issue-unit-age-ordered.scala 118:40]
  wire  _T_385 = _T_379 | (issue_slots_6_request & _T_361 | (_T_349 | (_T_334 | (issue_slots_3_request & _T_316 | (
    _T_304 | (_T_289 | issue_slots_0_request & _T_271)))))); // @[issue-unit-age-ordered.scala 124:69]
  wire  issue_slots_8_grant = issue_slots_8_request & _T_391 & ~_T_385; // @[issue-unit-age-ordered.scala 118:56]
  wire [1:0] _T_69 = issue_slots_7_grant + issue_slots_8_grant; // @[Bitwise.scala 47:55]
  wire  issue_slots_6_grant = _T_369 & ~_T_355; // @[issue-unit-age-ordered.scala 118:56]
  wire [1:0] _GEN_2933 = {{1'd0}, issue_slots_6_grant}; // @[Bitwise.scala 47:55]
  wire [2:0] _T_71 = _GEN_2933 + _T_69; // @[Bitwise.scala 47:55]
  wire  issue_slots_10_request = slots_10_io_request; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_10_uop_fu_code = slots_10_io_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] _T_420 = issue_slots_10_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 116:54]
  wire  _T_421 = _T_420 != 10'h0; // @[issue-unit-age-ordered.scala 116:72]
  wire  _T_424 = issue_slots_10_request & _T_421; // @[issue-unit-age-ordered.scala 118:40]
  wire  issue_slots_9_request = slots_9_io_request; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_9_uop_fu_code = slots_9_io_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] _T_405 = issue_slots_9_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 116:54]
  wire  _T_406 = _T_405 != 10'h0; // @[issue-unit-age-ordered.scala 116:72]
  wire  _T_414 = issue_slots_9_request & _T_406; // @[issue-unit-age-ordered.scala 124:52]
  wire  _T_400 = _T_394 | (_T_379 | (issue_slots_6_request & _T_361 | (_T_349 | (_T_334 | (issue_slots_3_request &
    _T_316 | (_T_304 | (_T_289 | issue_slots_0_request & _T_271))))))); // @[issue-unit-age-ordered.scala 124:69]
  wire  _T_415 = issue_slots_9_request & _T_406 | (_T_394 | (_T_379 | (issue_slots_6_request & _T_361 | (_T_349 | (
    _T_334 | (issue_slots_3_request & _T_316 | (_T_304 | (_T_289 | issue_slots_0_request & _T_271)))))))); // @[issue-unit-age-ordered.scala 124:69]
  wire  issue_slots_10_grant = issue_slots_10_request & _T_421 & ~_T_415; // @[issue-unit-age-ordered.scala 118:56]
  wire  issue_slots_11_request = slots_11_io_request; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_11_uop_fu_code = slots_11_io_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] _T_435 = issue_slots_11_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 116:54]
  wire  _T_436 = _T_435 != 10'h0; // @[issue-unit-age-ordered.scala 116:72]
  wire  _T_430 = _T_424 | (issue_slots_9_request & _T_406 | (_T_394 | (_T_379 | (issue_slots_6_request & _T_361 | (
    _T_349 | (_T_334 | (issue_slots_3_request & _T_316 | (_T_304 | (_T_289 | issue_slots_0_request & _T_271))))))))); // @[issue-unit-age-ordered.scala 124:69]
  wire  issue_slots_11_grant = issue_slots_11_request & _T_436 & ~_T_430; // @[issue-unit-age-ordered.scala 118:56]
  wire [1:0] _T_73 = issue_slots_10_grant + issue_slots_11_grant; // @[Bitwise.scala 47:55]
  wire  issue_slots_9_grant = _T_414 & ~_T_400; // @[issue-unit-age-ordered.scala 118:56]
  wire [1:0] _GEN_2934 = {{1'd0}, issue_slots_9_grant}; // @[Bitwise.scala 47:55]
  wire [2:0] _T_75 = _GEN_2934 + _T_73; // @[Bitwise.scala 47:55]
  wire [2:0] _T_77 = _T_71[1:0] + _T_75[1:0]; // @[Bitwise.scala 47:55]
  wire [3:0] _T_79 = _T_67 + _T_77; // @[Bitwise.scala 47:55]
  wire  vacants_0 = ~issue_slots_0_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_1 = ~issue_slots_1_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_2 = ~issue_slots_2_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_3 = ~issue_slots_3_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_4 = ~issue_slots_4_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_5 = ~issue_slots_5_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_6 = ~issue_slots_6_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_7 = ~issue_slots_7_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_8 = ~issue_slots_8_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_9 = ~issue_slots_9_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_10 = ~issue_slots_10_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_11 = ~issue_slots_11_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_12 = ~io_dis_uops_0_valid; // @[issue-unit-age-ordered.scala 39:82]
  wire [2:0] _GEN_11 = vacants_0 ? 3'h1 : 3'h0; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_98 = {_GEN_11[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_12 = ~_GEN_11[1] & vacants_1 ? _T_98 : {{1'd0}, _GEN_11[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_13 = _GEN_11[1:0] == 2'h0 & vacants_1 ? 3'h1 : _GEN_12; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_104 = {_GEN_13[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_14 = ~_GEN_13[1] & vacants_2 ? _T_104 : {{1'd0}, _GEN_13[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_15 = _GEN_13[1:0] == 2'h0 & vacants_2 ? 3'h1 : _GEN_14; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_110 = {_GEN_15[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_16 = ~_GEN_15[1] & vacants_3 ? _T_110 : {{1'd0}, _GEN_15[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_17 = _GEN_15[1:0] == 2'h0 & vacants_3 ? 3'h1 : _GEN_16; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_116 = {_GEN_17[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_18 = ~_GEN_17[1] & vacants_4 ? _T_116 : {{1'd0}, _GEN_17[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_19 = _GEN_17[1:0] == 2'h0 & vacants_4 ? 3'h1 : _GEN_18; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_122 = {_GEN_19[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_20 = ~_GEN_19[1] & vacants_5 ? _T_122 : {{1'd0}, _GEN_19[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_21 = _GEN_19[1:0] == 2'h0 & vacants_5 ? 3'h1 : _GEN_20; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_128 = {_GEN_21[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_22 = ~_GEN_21[1] & vacants_6 ? _T_128 : {{1'd0}, _GEN_21[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_23 = _GEN_21[1:0] == 2'h0 & vacants_6 ? 3'h1 : _GEN_22; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_134 = {_GEN_23[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_24 = ~_GEN_23[1] & vacants_7 ? _T_134 : {{1'd0}, _GEN_23[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_25 = _GEN_23[1:0] == 2'h0 & vacants_7 ? 3'h1 : _GEN_24; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_140 = {_GEN_25[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_26 = ~_GEN_25[1] & vacants_8 ? _T_140 : {{1'd0}, _GEN_25[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_27 = _GEN_25[1:0] == 2'h0 & vacants_8 ? 3'h1 : _GEN_26; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_146 = {_GEN_27[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_28 = ~_GEN_27[1] & vacants_9 ? _T_146 : {{1'd0}, _GEN_27[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_29 = _GEN_27[1:0] == 2'h0 & vacants_9 ? 3'h1 : _GEN_28; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_152 = {_GEN_29[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_30 = ~_GEN_29[1] & vacants_10 ? _T_152 : {{1'd0}, _GEN_29[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_31 = _GEN_29[1:0] == 2'h0 & vacants_10 ? 3'h1 : _GEN_30; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_158 = {_GEN_31[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_32 = ~_GEN_31[1] & vacants_11 ? _T_158 : {{1'd0}, _GEN_31[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_33 = _GEN_31[1:0] == 2'h0 & vacants_11 ? 3'h1 : _GEN_32; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_164 = {_GEN_33[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_34 = ~_GEN_33[1] & vacants_12 ? _T_164 : {{1'd0}, _GEN_33[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_35 = _GEN_33[1:0] == 2'h0 & vacants_12 ? 3'h1 : _GEN_34; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire  _T_165 = ~io_dis_uops_0_bits_exception; // @[issue-unit-age-ordered.scala 62:57]
  wire  _T_166 = io_dis_uops_0_valid & _T_165; // @[issue-unit-age-ordered.scala 61:77]
  wire  _T_167 = ~io_dis_uops_0_bits_is_fence; // @[issue-unit-age-ordered.scala 63:57]
  wire  _T_168 = _T_166 & _T_167; // @[issue-unit-age-ordered.scala 62:80]
  wire  _T_169 = ~io_dis_uops_0_bits_is_fencei; // @[issue-unit-age-ordered.scala 64:57]
  wire  will_be_valid_12 = _T_168 & _T_169; // @[issue-unit-age-ordered.scala 63:79]
  wire  _T_170 = ~io_dis_uops_1_bits_exception; // @[issue-unit-age-ordered.scala 62:57]
  wire  _T_171 = io_dis_uops_1_valid & _T_170; // @[issue-unit-age-ordered.scala 61:77]
  wire  _T_172 = ~io_dis_uops_1_bits_is_fence; // @[issue-unit-age-ordered.scala 63:57]
  wire  _T_173 = _T_171 & _T_172; // @[issue-unit-age-ordered.scala 62:80]
  wire  _T_174 = ~io_dis_uops_1_bits_is_fencei; // @[issue-unit-age-ordered.scala 64:57]
  wire  will_be_valid_13 = _T_173 & _T_174; // @[issue-unit-age-ordered.scala 63:79]
  wire  issue_slots_1_will_be_valid = slots_1_io_will_be_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_36 = _GEN_11[1:0] == 2'h1 & issue_slots_1_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire [1:0] issue_slots_1_out_uop_debug_tsrc = slots_1_io_out_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_1_out_uop_debug_fsrc = slots_1_io_out_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_bp_xcpt_if = slots_1_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_bp_debug_if = slots_1_io_out_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_xcpt_ma_if = slots_1_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_xcpt_ae_if = slots_1_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_xcpt_pf_if = slots_1_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_fp_single = slots_1_io_out_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_fp_val = slots_1_io_out_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_frs3_en = slots_1_io_out_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_1_out_uop_lrs2_rtype = slots_1_io_out_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_1_out_uop_lrs1_rtype = slots_1_io_out_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_1_out_uop_dst_rtype = slots_1_io_out_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_ldst_val = slots_1_io_out_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_1_out_uop_lrs3 = slots_1_io_out_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_1_out_uop_lrs2 = slots_1_io_out_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_1_out_uop_lrs1 = slots_1_io_out_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_1_out_uop_ldst = slots_1_io_out_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_ldst_is_rs1 = slots_1_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_flush_on_commit = slots_1_io_out_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_is_unique = slots_1_io_out_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_is_sys_pc2epc = slots_1_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_uses_stq = slots_1_io_out_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_uses_ldq = slots_1_io_out_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_is_amo = slots_1_io_out_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_is_fencei = slots_1_io_out_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_is_fence = slots_1_io_out_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_mem_signed = slots_1_io_out_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_1_out_uop_mem_size = slots_1_io_out_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_1_out_uop_mem_cmd = slots_1_io_out_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_bypassable = slots_1_io_out_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] issue_slots_1_out_uop_exc_cause = slots_1_io_out_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_exception = slots_1_io_out_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_1_out_uop_stale_pdst = slots_1_io_out_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_ppred_busy = slots_1_io_out_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_prs3_busy = slots_1_io_out_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_prs2_busy = slots_1_io_out_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_prs1_busy = slots_1_io_out_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_1_out_uop_ppred = slots_1_io_out_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_1_out_uop_prs3 = slots_1_io_out_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_1_out_uop_prs2 = slots_1_io_out_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_1_out_uop_prs1 = slots_1_io_out_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_1_out_uop_pdst = slots_1_io_out_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_1_out_uop_rxq_idx = slots_1_io_out_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_1_out_uop_stq_idx = slots_1_io_out_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_1_out_uop_ldq_idx = slots_1_io_out_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_1_out_uop_rob_idx = slots_1_io_out_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_1_out_uop_csr_addr = slots_1_io_out_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] issue_slots_1_out_uop_imm_packed = slots_1_io_out_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_taken = slots_1_io_out_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_1_out_uop_pc_lob = slots_1_io_out_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_edge_inst = slots_1_io_out_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_1_out_uop_ftq_idx = slots_1_io_out_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_1_out_uop_br_tag = slots_1_io_out_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_1_out_uop_br_mask = slots_1_io_out_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_is_sfb = slots_1_io_out_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_is_jal = slots_1_io_out_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_is_jalr = slots_1_io_out_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_is_br = slots_1_io_out_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_iw_p2_poisoned = slots_1_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_iw_p1_poisoned = slots_1_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_1_out_uop_iw_state = slots_1_io_out_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_ctrl_is_std = slots_1_io_out_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_ctrl_is_sta = slots_1_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_ctrl_is_load = slots_1_io_out_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_1_out_uop_ctrl_csr_cmd = slots_1_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_ctrl_fcn_dw = slots_1_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_1_out_uop_ctrl_op_fcn = slots_1_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_1_out_uop_ctrl_imm_sel = slots_1_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_1_out_uop_ctrl_op2_sel = slots_1_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_1_out_uop_ctrl_op1_sel = slots_1_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_1_out_uop_ctrl_br_type = slots_1_io_out_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_1_out_uop_fu_code = slots_1_io_out_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_1_out_uop_iq_type = slots_1_io_out_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] issue_slots_1_out_uop_debug_pc = slots_1_io_out_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_out_uop_is_rvc = slots_1_io_out_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_1_out_uop_debug_inst = slots_1_io_out_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_1_out_uop_inst = slots_1_io_out_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] issue_slots_1_out_uop_uopc = slots_1_io_out_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_will_be_valid = slots_2_io_will_be_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_0_in_uop_valid = _GEN_13[1:0] == 2'h2 ? issue_slots_2_will_be_valid : _GEN_36; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_2_out_uop_debug_tsrc = slots_2_io_out_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_2_out_uop_debug_fsrc = slots_2_io_out_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_bp_xcpt_if = slots_2_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_bp_debug_if = slots_2_io_out_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_xcpt_ma_if = slots_2_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_xcpt_ae_if = slots_2_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_xcpt_pf_if = slots_2_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_fp_single = slots_2_io_out_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_fp_val = slots_2_io_out_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_frs3_en = slots_2_io_out_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_2_out_uop_lrs2_rtype = slots_2_io_out_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_2_out_uop_lrs1_rtype = slots_2_io_out_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_2_out_uop_dst_rtype = slots_2_io_out_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_ldst_val = slots_2_io_out_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_2_out_uop_lrs3 = slots_2_io_out_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_2_out_uop_lrs2 = slots_2_io_out_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_2_out_uop_lrs1 = slots_2_io_out_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_2_out_uop_ldst = slots_2_io_out_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_ldst_is_rs1 = slots_2_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_flush_on_commit = slots_2_io_out_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_is_unique = slots_2_io_out_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_is_sys_pc2epc = slots_2_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_uses_stq = slots_2_io_out_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_uses_ldq = slots_2_io_out_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_is_amo = slots_2_io_out_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_is_fencei = slots_2_io_out_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_is_fence = slots_2_io_out_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_mem_signed = slots_2_io_out_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_2_out_uop_mem_size = slots_2_io_out_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_2_out_uop_mem_cmd = slots_2_io_out_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_bypassable = slots_2_io_out_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] issue_slots_2_out_uop_exc_cause = slots_2_io_out_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_exception = slots_2_io_out_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_2_out_uop_stale_pdst = slots_2_io_out_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_ppred_busy = slots_2_io_out_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_prs3_busy = slots_2_io_out_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_prs2_busy = slots_2_io_out_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_prs1_busy = slots_2_io_out_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_2_out_uop_ppred = slots_2_io_out_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_2_out_uop_prs3 = slots_2_io_out_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_2_out_uop_prs2 = slots_2_io_out_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_2_out_uop_prs1 = slots_2_io_out_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_2_out_uop_pdst = slots_2_io_out_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_2_out_uop_rxq_idx = slots_2_io_out_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_2_out_uop_stq_idx = slots_2_io_out_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_2_out_uop_ldq_idx = slots_2_io_out_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_2_out_uop_rob_idx = slots_2_io_out_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_2_out_uop_csr_addr = slots_2_io_out_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] issue_slots_2_out_uop_imm_packed = slots_2_io_out_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_taken = slots_2_io_out_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_2_out_uop_pc_lob = slots_2_io_out_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_edge_inst = slots_2_io_out_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_2_out_uop_ftq_idx = slots_2_io_out_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_2_out_uop_br_tag = slots_2_io_out_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_2_out_uop_br_mask = slots_2_io_out_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_is_sfb = slots_2_io_out_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_is_jal = slots_2_io_out_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_is_jalr = slots_2_io_out_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_is_br = slots_2_io_out_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_iw_p2_poisoned = slots_2_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_iw_p1_poisoned = slots_2_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_2_out_uop_iw_state = slots_2_io_out_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_ctrl_is_std = slots_2_io_out_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_ctrl_is_sta = slots_2_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_ctrl_is_load = slots_2_io_out_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_2_out_uop_ctrl_csr_cmd = slots_2_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_ctrl_fcn_dw = slots_2_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_2_out_uop_ctrl_op_fcn = slots_2_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_2_out_uop_ctrl_imm_sel = slots_2_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_2_out_uop_ctrl_op2_sel = slots_2_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_2_out_uop_ctrl_op1_sel = slots_2_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_2_out_uop_ctrl_br_type = slots_2_io_out_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_2_out_uop_fu_code = slots_2_io_out_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_2_out_uop_iq_type = slots_2_io_out_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] issue_slots_2_out_uop_debug_pc = slots_2_io_out_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_out_uop_is_rvc = slots_2_io_out_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_2_out_uop_debug_inst = slots_2_io_out_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_2_out_uop_inst = slots_2_io_out_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] issue_slots_2_out_uop_uopc = slots_2_io_out_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_196 = _GEN_13[1:0] == 2'h1 & issue_slots_2_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_3_will_be_valid = slots_3_io_will_be_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_in_uop_valid = _GEN_15[1:0] == 2'h2 ? issue_slots_3_will_be_valid : _GEN_196; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_3_out_uop_debug_tsrc = slots_3_io_out_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_3_out_uop_debug_fsrc = slots_3_io_out_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_bp_xcpt_if = slots_3_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_bp_debug_if = slots_3_io_out_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_xcpt_ma_if = slots_3_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_xcpt_ae_if = slots_3_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_xcpt_pf_if = slots_3_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_fp_single = slots_3_io_out_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_fp_val = slots_3_io_out_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_frs3_en = slots_3_io_out_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_3_out_uop_lrs2_rtype = slots_3_io_out_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_3_out_uop_lrs1_rtype = slots_3_io_out_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_3_out_uop_dst_rtype = slots_3_io_out_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_ldst_val = slots_3_io_out_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_3_out_uop_lrs3 = slots_3_io_out_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_3_out_uop_lrs2 = slots_3_io_out_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_3_out_uop_lrs1 = slots_3_io_out_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_3_out_uop_ldst = slots_3_io_out_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_ldst_is_rs1 = slots_3_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_flush_on_commit = slots_3_io_out_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_is_unique = slots_3_io_out_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_is_sys_pc2epc = slots_3_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_uses_stq = slots_3_io_out_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_uses_ldq = slots_3_io_out_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_is_amo = slots_3_io_out_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_is_fencei = slots_3_io_out_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_is_fence = slots_3_io_out_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_mem_signed = slots_3_io_out_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_3_out_uop_mem_size = slots_3_io_out_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_3_out_uop_mem_cmd = slots_3_io_out_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_bypassable = slots_3_io_out_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] issue_slots_3_out_uop_exc_cause = slots_3_io_out_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_exception = slots_3_io_out_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_3_out_uop_stale_pdst = slots_3_io_out_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_ppred_busy = slots_3_io_out_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_prs3_busy = slots_3_io_out_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_prs2_busy = slots_3_io_out_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_prs1_busy = slots_3_io_out_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_3_out_uop_ppred = slots_3_io_out_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_3_out_uop_prs3 = slots_3_io_out_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_3_out_uop_prs2 = slots_3_io_out_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_3_out_uop_prs1 = slots_3_io_out_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_3_out_uop_pdst = slots_3_io_out_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_3_out_uop_rxq_idx = slots_3_io_out_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_3_out_uop_stq_idx = slots_3_io_out_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_3_out_uop_ldq_idx = slots_3_io_out_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_3_out_uop_rob_idx = slots_3_io_out_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_3_out_uop_csr_addr = slots_3_io_out_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] issue_slots_3_out_uop_imm_packed = slots_3_io_out_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_taken = slots_3_io_out_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_3_out_uop_pc_lob = slots_3_io_out_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_edge_inst = slots_3_io_out_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_3_out_uop_ftq_idx = slots_3_io_out_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_3_out_uop_br_tag = slots_3_io_out_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_3_out_uop_br_mask = slots_3_io_out_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_is_sfb = slots_3_io_out_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_is_jal = slots_3_io_out_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_is_jalr = slots_3_io_out_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_is_br = slots_3_io_out_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_iw_p2_poisoned = slots_3_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_iw_p1_poisoned = slots_3_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_3_out_uop_iw_state = slots_3_io_out_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_ctrl_is_std = slots_3_io_out_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_ctrl_is_sta = slots_3_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_ctrl_is_load = slots_3_io_out_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_3_out_uop_ctrl_csr_cmd = slots_3_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_ctrl_fcn_dw = slots_3_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_3_out_uop_ctrl_op_fcn = slots_3_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_3_out_uop_ctrl_imm_sel = slots_3_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_3_out_uop_ctrl_op2_sel = slots_3_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_3_out_uop_ctrl_op1_sel = slots_3_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_3_out_uop_ctrl_br_type = slots_3_io_out_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_3_out_uop_fu_code = slots_3_io_out_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_3_out_uop_iq_type = slots_3_io_out_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] issue_slots_3_out_uop_debug_pc = slots_3_io_out_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_out_uop_is_rvc = slots_3_io_out_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_3_out_uop_debug_inst = slots_3_io_out_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_3_out_uop_inst = slots_3_io_out_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] issue_slots_3_out_uop_uopc = slots_3_io_out_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_1_clear = _GEN_11[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_356 = _GEN_15[1:0] == 2'h1 & issue_slots_3_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_4_will_be_valid = slots_4_io_will_be_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_in_uop_valid = _GEN_17[1:0] == 2'h2 ? issue_slots_4_will_be_valid : _GEN_356; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_4_out_uop_debug_tsrc = slots_4_io_out_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_4_out_uop_debug_fsrc = slots_4_io_out_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_bp_xcpt_if = slots_4_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_bp_debug_if = slots_4_io_out_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_xcpt_ma_if = slots_4_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_xcpt_ae_if = slots_4_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_xcpt_pf_if = slots_4_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_fp_single = slots_4_io_out_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_fp_val = slots_4_io_out_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_frs3_en = slots_4_io_out_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_4_out_uop_lrs2_rtype = slots_4_io_out_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_4_out_uop_lrs1_rtype = slots_4_io_out_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_4_out_uop_dst_rtype = slots_4_io_out_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_ldst_val = slots_4_io_out_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_4_out_uop_lrs3 = slots_4_io_out_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_4_out_uop_lrs2 = slots_4_io_out_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_4_out_uop_lrs1 = slots_4_io_out_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_4_out_uop_ldst = slots_4_io_out_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_ldst_is_rs1 = slots_4_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_flush_on_commit = slots_4_io_out_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_is_unique = slots_4_io_out_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_is_sys_pc2epc = slots_4_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_uses_stq = slots_4_io_out_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_uses_ldq = slots_4_io_out_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_is_amo = slots_4_io_out_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_is_fencei = slots_4_io_out_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_is_fence = slots_4_io_out_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_mem_signed = slots_4_io_out_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_4_out_uop_mem_size = slots_4_io_out_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_4_out_uop_mem_cmd = slots_4_io_out_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_bypassable = slots_4_io_out_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] issue_slots_4_out_uop_exc_cause = slots_4_io_out_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_exception = slots_4_io_out_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_4_out_uop_stale_pdst = slots_4_io_out_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_ppred_busy = slots_4_io_out_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_prs3_busy = slots_4_io_out_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_prs2_busy = slots_4_io_out_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_prs1_busy = slots_4_io_out_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_4_out_uop_ppred = slots_4_io_out_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_4_out_uop_prs3 = slots_4_io_out_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_4_out_uop_prs2 = slots_4_io_out_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_4_out_uop_prs1 = slots_4_io_out_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_4_out_uop_pdst = slots_4_io_out_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_4_out_uop_rxq_idx = slots_4_io_out_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_4_out_uop_stq_idx = slots_4_io_out_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_4_out_uop_ldq_idx = slots_4_io_out_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_4_out_uop_rob_idx = slots_4_io_out_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_4_out_uop_csr_addr = slots_4_io_out_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] issue_slots_4_out_uop_imm_packed = slots_4_io_out_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_taken = slots_4_io_out_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_4_out_uop_pc_lob = slots_4_io_out_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_edge_inst = slots_4_io_out_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_4_out_uop_ftq_idx = slots_4_io_out_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_4_out_uop_br_tag = slots_4_io_out_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_4_out_uop_br_mask = slots_4_io_out_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_is_sfb = slots_4_io_out_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_is_jal = slots_4_io_out_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_is_jalr = slots_4_io_out_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_is_br = slots_4_io_out_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_iw_p2_poisoned = slots_4_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_iw_p1_poisoned = slots_4_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_4_out_uop_iw_state = slots_4_io_out_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_ctrl_is_std = slots_4_io_out_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_ctrl_is_sta = slots_4_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_ctrl_is_load = slots_4_io_out_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_4_out_uop_ctrl_csr_cmd = slots_4_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_ctrl_fcn_dw = slots_4_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_4_out_uop_ctrl_op_fcn = slots_4_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_4_out_uop_ctrl_imm_sel = slots_4_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_4_out_uop_ctrl_op2_sel = slots_4_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_4_out_uop_ctrl_op1_sel = slots_4_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_4_out_uop_ctrl_br_type = slots_4_io_out_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_4_out_uop_fu_code = slots_4_io_out_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_4_out_uop_iq_type = slots_4_io_out_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] issue_slots_4_out_uop_debug_pc = slots_4_io_out_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_out_uop_is_rvc = slots_4_io_out_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_4_out_uop_debug_inst = slots_4_io_out_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_4_out_uop_inst = slots_4_io_out_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] issue_slots_4_out_uop_uopc = slots_4_io_out_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_2_clear = _GEN_13[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_516 = _GEN_17[1:0] == 2'h1 & issue_slots_4_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_5_will_be_valid = slots_5_io_will_be_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_in_uop_valid = _GEN_19[1:0] == 2'h2 ? issue_slots_5_will_be_valid : _GEN_516; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_5_out_uop_debug_tsrc = slots_5_io_out_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_5_out_uop_debug_fsrc = slots_5_io_out_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_bp_xcpt_if = slots_5_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_bp_debug_if = slots_5_io_out_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_xcpt_ma_if = slots_5_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_xcpt_ae_if = slots_5_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_xcpt_pf_if = slots_5_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_fp_single = slots_5_io_out_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_fp_val = slots_5_io_out_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_frs3_en = slots_5_io_out_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_5_out_uop_lrs2_rtype = slots_5_io_out_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_5_out_uop_lrs1_rtype = slots_5_io_out_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_5_out_uop_dst_rtype = slots_5_io_out_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_ldst_val = slots_5_io_out_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_5_out_uop_lrs3 = slots_5_io_out_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_5_out_uop_lrs2 = slots_5_io_out_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_5_out_uop_lrs1 = slots_5_io_out_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_5_out_uop_ldst = slots_5_io_out_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_ldst_is_rs1 = slots_5_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_flush_on_commit = slots_5_io_out_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_is_unique = slots_5_io_out_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_is_sys_pc2epc = slots_5_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_uses_stq = slots_5_io_out_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_uses_ldq = slots_5_io_out_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_is_amo = slots_5_io_out_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_is_fencei = slots_5_io_out_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_is_fence = slots_5_io_out_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_mem_signed = slots_5_io_out_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_5_out_uop_mem_size = slots_5_io_out_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_5_out_uop_mem_cmd = slots_5_io_out_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_bypassable = slots_5_io_out_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] issue_slots_5_out_uop_exc_cause = slots_5_io_out_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_exception = slots_5_io_out_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_5_out_uop_stale_pdst = slots_5_io_out_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_ppred_busy = slots_5_io_out_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_prs3_busy = slots_5_io_out_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_prs2_busy = slots_5_io_out_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_prs1_busy = slots_5_io_out_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_5_out_uop_ppred = slots_5_io_out_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_5_out_uop_prs3 = slots_5_io_out_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_5_out_uop_prs2 = slots_5_io_out_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_5_out_uop_prs1 = slots_5_io_out_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_5_out_uop_pdst = slots_5_io_out_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_5_out_uop_rxq_idx = slots_5_io_out_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_5_out_uop_stq_idx = slots_5_io_out_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_5_out_uop_ldq_idx = slots_5_io_out_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_5_out_uop_rob_idx = slots_5_io_out_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_5_out_uop_csr_addr = slots_5_io_out_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] issue_slots_5_out_uop_imm_packed = slots_5_io_out_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_taken = slots_5_io_out_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_5_out_uop_pc_lob = slots_5_io_out_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_edge_inst = slots_5_io_out_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_5_out_uop_ftq_idx = slots_5_io_out_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_5_out_uop_br_tag = slots_5_io_out_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_5_out_uop_br_mask = slots_5_io_out_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_is_sfb = slots_5_io_out_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_is_jal = slots_5_io_out_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_is_jalr = slots_5_io_out_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_is_br = slots_5_io_out_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_iw_p2_poisoned = slots_5_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_iw_p1_poisoned = slots_5_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_5_out_uop_iw_state = slots_5_io_out_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_ctrl_is_std = slots_5_io_out_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_ctrl_is_sta = slots_5_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_ctrl_is_load = slots_5_io_out_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_5_out_uop_ctrl_csr_cmd = slots_5_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_ctrl_fcn_dw = slots_5_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_5_out_uop_ctrl_op_fcn = slots_5_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_5_out_uop_ctrl_imm_sel = slots_5_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_5_out_uop_ctrl_op2_sel = slots_5_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_5_out_uop_ctrl_op1_sel = slots_5_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_5_out_uop_ctrl_br_type = slots_5_io_out_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_5_out_uop_fu_code = slots_5_io_out_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_5_out_uop_iq_type = slots_5_io_out_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] issue_slots_5_out_uop_debug_pc = slots_5_io_out_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_out_uop_is_rvc = slots_5_io_out_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_5_out_uop_debug_inst = slots_5_io_out_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_5_out_uop_inst = slots_5_io_out_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] issue_slots_5_out_uop_uopc = slots_5_io_out_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_3_clear = _GEN_15[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_676 = _GEN_19[1:0] == 2'h1 & issue_slots_5_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_6_will_be_valid = slots_6_io_will_be_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_in_uop_valid = _GEN_21[1:0] == 2'h2 ? issue_slots_6_will_be_valid : _GEN_676; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_6_out_uop_debug_tsrc = slots_6_io_out_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_6_out_uop_debug_fsrc = slots_6_io_out_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_bp_xcpt_if = slots_6_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_bp_debug_if = slots_6_io_out_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_xcpt_ma_if = slots_6_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_xcpt_ae_if = slots_6_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_xcpt_pf_if = slots_6_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_fp_single = slots_6_io_out_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_fp_val = slots_6_io_out_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_frs3_en = slots_6_io_out_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_6_out_uop_lrs2_rtype = slots_6_io_out_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_6_out_uop_lrs1_rtype = slots_6_io_out_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_6_out_uop_dst_rtype = slots_6_io_out_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_ldst_val = slots_6_io_out_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_6_out_uop_lrs3 = slots_6_io_out_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_6_out_uop_lrs2 = slots_6_io_out_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_6_out_uop_lrs1 = slots_6_io_out_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_6_out_uop_ldst = slots_6_io_out_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_ldst_is_rs1 = slots_6_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_flush_on_commit = slots_6_io_out_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_is_unique = slots_6_io_out_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_is_sys_pc2epc = slots_6_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_uses_stq = slots_6_io_out_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_uses_ldq = slots_6_io_out_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_is_amo = slots_6_io_out_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_is_fencei = slots_6_io_out_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_is_fence = slots_6_io_out_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_mem_signed = slots_6_io_out_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_6_out_uop_mem_size = slots_6_io_out_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_6_out_uop_mem_cmd = slots_6_io_out_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_bypassable = slots_6_io_out_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] issue_slots_6_out_uop_exc_cause = slots_6_io_out_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_exception = slots_6_io_out_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_6_out_uop_stale_pdst = slots_6_io_out_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_ppred_busy = slots_6_io_out_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_prs3_busy = slots_6_io_out_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_prs2_busy = slots_6_io_out_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_prs1_busy = slots_6_io_out_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_6_out_uop_ppred = slots_6_io_out_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_6_out_uop_prs3 = slots_6_io_out_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_6_out_uop_prs2 = slots_6_io_out_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_6_out_uop_prs1 = slots_6_io_out_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_6_out_uop_pdst = slots_6_io_out_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_6_out_uop_rxq_idx = slots_6_io_out_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_6_out_uop_stq_idx = slots_6_io_out_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_6_out_uop_ldq_idx = slots_6_io_out_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_6_out_uop_rob_idx = slots_6_io_out_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_6_out_uop_csr_addr = slots_6_io_out_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] issue_slots_6_out_uop_imm_packed = slots_6_io_out_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_taken = slots_6_io_out_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_6_out_uop_pc_lob = slots_6_io_out_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_edge_inst = slots_6_io_out_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_6_out_uop_ftq_idx = slots_6_io_out_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_6_out_uop_br_tag = slots_6_io_out_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_6_out_uop_br_mask = slots_6_io_out_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_is_sfb = slots_6_io_out_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_is_jal = slots_6_io_out_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_is_jalr = slots_6_io_out_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_is_br = slots_6_io_out_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_iw_p2_poisoned = slots_6_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_iw_p1_poisoned = slots_6_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_6_out_uop_iw_state = slots_6_io_out_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_ctrl_is_std = slots_6_io_out_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_ctrl_is_sta = slots_6_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_ctrl_is_load = slots_6_io_out_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_6_out_uop_ctrl_csr_cmd = slots_6_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_ctrl_fcn_dw = slots_6_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_6_out_uop_ctrl_op_fcn = slots_6_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_6_out_uop_ctrl_imm_sel = slots_6_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_6_out_uop_ctrl_op2_sel = slots_6_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_6_out_uop_ctrl_op1_sel = slots_6_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_6_out_uop_ctrl_br_type = slots_6_io_out_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_6_out_uop_fu_code = slots_6_io_out_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_6_out_uop_iq_type = slots_6_io_out_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] issue_slots_6_out_uop_debug_pc = slots_6_io_out_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_out_uop_is_rvc = slots_6_io_out_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_6_out_uop_debug_inst = slots_6_io_out_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_6_out_uop_inst = slots_6_io_out_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] issue_slots_6_out_uop_uopc = slots_6_io_out_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_4_clear = _GEN_17[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_836 = _GEN_21[1:0] == 2'h1 & issue_slots_6_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_7_will_be_valid = slots_7_io_will_be_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_in_uop_valid = _GEN_23[1:0] == 2'h2 ? issue_slots_7_will_be_valid : _GEN_836; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_7_out_uop_debug_tsrc = slots_7_io_out_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_7_out_uop_debug_fsrc = slots_7_io_out_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_bp_xcpt_if = slots_7_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_bp_debug_if = slots_7_io_out_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_xcpt_ma_if = slots_7_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_xcpt_ae_if = slots_7_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_xcpt_pf_if = slots_7_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_fp_single = slots_7_io_out_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_fp_val = slots_7_io_out_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_frs3_en = slots_7_io_out_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_7_out_uop_lrs2_rtype = slots_7_io_out_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_7_out_uop_lrs1_rtype = slots_7_io_out_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_7_out_uop_dst_rtype = slots_7_io_out_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_ldst_val = slots_7_io_out_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_7_out_uop_lrs3 = slots_7_io_out_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_7_out_uop_lrs2 = slots_7_io_out_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_7_out_uop_lrs1 = slots_7_io_out_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_7_out_uop_ldst = slots_7_io_out_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_ldst_is_rs1 = slots_7_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_flush_on_commit = slots_7_io_out_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_is_unique = slots_7_io_out_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_is_sys_pc2epc = slots_7_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_uses_stq = slots_7_io_out_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_uses_ldq = slots_7_io_out_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_is_amo = slots_7_io_out_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_is_fencei = slots_7_io_out_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_is_fence = slots_7_io_out_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_mem_signed = slots_7_io_out_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_7_out_uop_mem_size = slots_7_io_out_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_7_out_uop_mem_cmd = slots_7_io_out_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_bypassable = slots_7_io_out_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] issue_slots_7_out_uop_exc_cause = slots_7_io_out_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_exception = slots_7_io_out_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_7_out_uop_stale_pdst = slots_7_io_out_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_ppred_busy = slots_7_io_out_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_prs3_busy = slots_7_io_out_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_prs2_busy = slots_7_io_out_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_prs1_busy = slots_7_io_out_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_7_out_uop_ppred = slots_7_io_out_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_7_out_uop_prs3 = slots_7_io_out_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_7_out_uop_prs2 = slots_7_io_out_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_7_out_uop_prs1 = slots_7_io_out_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_7_out_uop_pdst = slots_7_io_out_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_7_out_uop_rxq_idx = slots_7_io_out_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_7_out_uop_stq_idx = slots_7_io_out_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_7_out_uop_ldq_idx = slots_7_io_out_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_7_out_uop_rob_idx = slots_7_io_out_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_7_out_uop_csr_addr = slots_7_io_out_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] issue_slots_7_out_uop_imm_packed = slots_7_io_out_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_taken = slots_7_io_out_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_7_out_uop_pc_lob = slots_7_io_out_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_edge_inst = slots_7_io_out_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_7_out_uop_ftq_idx = slots_7_io_out_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_7_out_uop_br_tag = slots_7_io_out_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_7_out_uop_br_mask = slots_7_io_out_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_is_sfb = slots_7_io_out_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_is_jal = slots_7_io_out_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_is_jalr = slots_7_io_out_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_is_br = slots_7_io_out_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_iw_p2_poisoned = slots_7_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_iw_p1_poisoned = slots_7_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_7_out_uop_iw_state = slots_7_io_out_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_ctrl_is_std = slots_7_io_out_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_ctrl_is_sta = slots_7_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_ctrl_is_load = slots_7_io_out_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_7_out_uop_ctrl_csr_cmd = slots_7_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_ctrl_fcn_dw = slots_7_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_7_out_uop_ctrl_op_fcn = slots_7_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_7_out_uop_ctrl_imm_sel = slots_7_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_7_out_uop_ctrl_op2_sel = slots_7_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_7_out_uop_ctrl_op1_sel = slots_7_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_7_out_uop_ctrl_br_type = slots_7_io_out_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_7_out_uop_fu_code = slots_7_io_out_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_7_out_uop_iq_type = slots_7_io_out_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] issue_slots_7_out_uop_debug_pc = slots_7_io_out_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_out_uop_is_rvc = slots_7_io_out_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_7_out_uop_debug_inst = slots_7_io_out_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_7_out_uop_inst = slots_7_io_out_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] issue_slots_7_out_uop_uopc = slots_7_io_out_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_5_clear = _GEN_19[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_996 = _GEN_23[1:0] == 2'h1 & issue_slots_7_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_8_will_be_valid = slots_8_io_will_be_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_in_uop_valid = _GEN_25[1:0] == 2'h2 ? issue_slots_8_will_be_valid : _GEN_996; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_8_out_uop_debug_tsrc = slots_8_io_out_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_8_out_uop_debug_fsrc = slots_8_io_out_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_bp_xcpt_if = slots_8_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_bp_debug_if = slots_8_io_out_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_xcpt_ma_if = slots_8_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_xcpt_ae_if = slots_8_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_xcpt_pf_if = slots_8_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_fp_single = slots_8_io_out_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_fp_val = slots_8_io_out_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_frs3_en = slots_8_io_out_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_8_out_uop_lrs2_rtype = slots_8_io_out_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_8_out_uop_lrs1_rtype = slots_8_io_out_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_8_out_uop_dst_rtype = slots_8_io_out_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_ldst_val = slots_8_io_out_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_8_out_uop_lrs3 = slots_8_io_out_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_8_out_uop_lrs2 = slots_8_io_out_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_8_out_uop_lrs1 = slots_8_io_out_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_8_out_uop_ldst = slots_8_io_out_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_ldst_is_rs1 = slots_8_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_flush_on_commit = slots_8_io_out_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_is_unique = slots_8_io_out_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_is_sys_pc2epc = slots_8_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_uses_stq = slots_8_io_out_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_uses_ldq = slots_8_io_out_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_is_amo = slots_8_io_out_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_is_fencei = slots_8_io_out_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_is_fence = slots_8_io_out_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_mem_signed = slots_8_io_out_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_8_out_uop_mem_size = slots_8_io_out_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_8_out_uop_mem_cmd = slots_8_io_out_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_bypassable = slots_8_io_out_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] issue_slots_8_out_uop_exc_cause = slots_8_io_out_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_exception = slots_8_io_out_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_8_out_uop_stale_pdst = slots_8_io_out_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_ppred_busy = slots_8_io_out_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_prs3_busy = slots_8_io_out_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_prs2_busy = slots_8_io_out_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_prs1_busy = slots_8_io_out_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_8_out_uop_ppred = slots_8_io_out_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_8_out_uop_prs3 = slots_8_io_out_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_8_out_uop_prs2 = slots_8_io_out_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_8_out_uop_prs1 = slots_8_io_out_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_8_out_uop_pdst = slots_8_io_out_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_8_out_uop_rxq_idx = slots_8_io_out_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_8_out_uop_stq_idx = slots_8_io_out_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_8_out_uop_ldq_idx = slots_8_io_out_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_8_out_uop_rob_idx = slots_8_io_out_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_8_out_uop_csr_addr = slots_8_io_out_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] issue_slots_8_out_uop_imm_packed = slots_8_io_out_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_taken = slots_8_io_out_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_8_out_uop_pc_lob = slots_8_io_out_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_edge_inst = slots_8_io_out_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_8_out_uop_ftq_idx = slots_8_io_out_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_8_out_uop_br_tag = slots_8_io_out_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_8_out_uop_br_mask = slots_8_io_out_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_is_sfb = slots_8_io_out_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_is_jal = slots_8_io_out_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_is_jalr = slots_8_io_out_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_is_br = slots_8_io_out_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_iw_p2_poisoned = slots_8_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_iw_p1_poisoned = slots_8_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_8_out_uop_iw_state = slots_8_io_out_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_ctrl_is_std = slots_8_io_out_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_ctrl_is_sta = slots_8_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_ctrl_is_load = slots_8_io_out_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_8_out_uop_ctrl_csr_cmd = slots_8_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_ctrl_fcn_dw = slots_8_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_8_out_uop_ctrl_op_fcn = slots_8_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_8_out_uop_ctrl_imm_sel = slots_8_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_8_out_uop_ctrl_op2_sel = slots_8_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_8_out_uop_ctrl_op1_sel = slots_8_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_8_out_uop_ctrl_br_type = slots_8_io_out_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_8_out_uop_fu_code = slots_8_io_out_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_8_out_uop_iq_type = slots_8_io_out_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] issue_slots_8_out_uop_debug_pc = slots_8_io_out_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_out_uop_is_rvc = slots_8_io_out_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_8_out_uop_debug_inst = slots_8_io_out_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_8_out_uop_inst = slots_8_io_out_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] issue_slots_8_out_uop_uopc = slots_8_io_out_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_6_clear = _GEN_21[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_1156 = _GEN_25[1:0] == 2'h1 & issue_slots_8_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_9_will_be_valid = slots_9_io_will_be_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_in_uop_valid = _GEN_27[1:0] == 2'h2 ? issue_slots_9_will_be_valid : _GEN_1156; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_9_out_uop_debug_tsrc = slots_9_io_out_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_9_out_uop_debug_fsrc = slots_9_io_out_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_bp_xcpt_if = slots_9_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_bp_debug_if = slots_9_io_out_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_xcpt_ma_if = slots_9_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_xcpt_ae_if = slots_9_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_xcpt_pf_if = slots_9_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_fp_single = slots_9_io_out_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_fp_val = slots_9_io_out_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_frs3_en = slots_9_io_out_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_9_out_uop_lrs2_rtype = slots_9_io_out_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_9_out_uop_lrs1_rtype = slots_9_io_out_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_9_out_uop_dst_rtype = slots_9_io_out_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_ldst_val = slots_9_io_out_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_9_out_uop_lrs3 = slots_9_io_out_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_9_out_uop_lrs2 = slots_9_io_out_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_9_out_uop_lrs1 = slots_9_io_out_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_9_out_uop_ldst = slots_9_io_out_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_ldst_is_rs1 = slots_9_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_flush_on_commit = slots_9_io_out_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_is_unique = slots_9_io_out_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_is_sys_pc2epc = slots_9_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_uses_stq = slots_9_io_out_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_uses_ldq = slots_9_io_out_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_is_amo = slots_9_io_out_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_is_fencei = slots_9_io_out_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_is_fence = slots_9_io_out_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_mem_signed = slots_9_io_out_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_9_out_uop_mem_size = slots_9_io_out_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_9_out_uop_mem_cmd = slots_9_io_out_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_bypassable = slots_9_io_out_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] issue_slots_9_out_uop_exc_cause = slots_9_io_out_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_exception = slots_9_io_out_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_9_out_uop_stale_pdst = slots_9_io_out_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_ppred_busy = slots_9_io_out_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_prs3_busy = slots_9_io_out_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_prs2_busy = slots_9_io_out_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_prs1_busy = slots_9_io_out_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_9_out_uop_ppred = slots_9_io_out_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_9_out_uop_prs3 = slots_9_io_out_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_9_out_uop_prs2 = slots_9_io_out_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_9_out_uop_prs1 = slots_9_io_out_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_9_out_uop_pdst = slots_9_io_out_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_9_out_uop_rxq_idx = slots_9_io_out_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_9_out_uop_stq_idx = slots_9_io_out_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_9_out_uop_ldq_idx = slots_9_io_out_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_9_out_uop_rob_idx = slots_9_io_out_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_9_out_uop_csr_addr = slots_9_io_out_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] issue_slots_9_out_uop_imm_packed = slots_9_io_out_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_taken = slots_9_io_out_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_9_out_uop_pc_lob = slots_9_io_out_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_edge_inst = slots_9_io_out_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_9_out_uop_ftq_idx = slots_9_io_out_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_9_out_uop_br_tag = slots_9_io_out_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_9_out_uop_br_mask = slots_9_io_out_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_is_sfb = slots_9_io_out_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_is_jal = slots_9_io_out_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_is_jalr = slots_9_io_out_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_is_br = slots_9_io_out_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_iw_p2_poisoned = slots_9_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_iw_p1_poisoned = slots_9_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_9_out_uop_iw_state = slots_9_io_out_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_ctrl_is_std = slots_9_io_out_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_ctrl_is_sta = slots_9_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_ctrl_is_load = slots_9_io_out_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_9_out_uop_ctrl_csr_cmd = slots_9_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_ctrl_fcn_dw = slots_9_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_9_out_uop_ctrl_op_fcn = slots_9_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_9_out_uop_ctrl_imm_sel = slots_9_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_9_out_uop_ctrl_op2_sel = slots_9_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_9_out_uop_ctrl_op1_sel = slots_9_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_9_out_uop_ctrl_br_type = slots_9_io_out_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_9_out_uop_fu_code = slots_9_io_out_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_9_out_uop_iq_type = slots_9_io_out_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] issue_slots_9_out_uop_debug_pc = slots_9_io_out_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_out_uop_is_rvc = slots_9_io_out_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_9_out_uop_debug_inst = slots_9_io_out_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_9_out_uop_inst = slots_9_io_out_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] issue_slots_9_out_uop_uopc = slots_9_io_out_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_7_clear = _GEN_23[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_1316 = _GEN_27[1:0] == 2'h1 & issue_slots_9_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_10_will_be_valid = slots_10_io_will_be_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_in_uop_valid = _GEN_29[1:0] == 2'h2 ? issue_slots_10_will_be_valid : _GEN_1316; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_10_out_uop_debug_tsrc = slots_10_io_out_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_10_out_uop_debug_fsrc = slots_10_io_out_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_bp_xcpt_if = slots_10_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_bp_debug_if = slots_10_io_out_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_xcpt_ma_if = slots_10_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_xcpt_ae_if = slots_10_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_xcpt_pf_if = slots_10_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_fp_single = slots_10_io_out_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_fp_val = slots_10_io_out_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_frs3_en = slots_10_io_out_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_10_out_uop_lrs2_rtype = slots_10_io_out_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_10_out_uop_lrs1_rtype = slots_10_io_out_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_10_out_uop_dst_rtype = slots_10_io_out_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_ldst_val = slots_10_io_out_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_10_out_uop_lrs3 = slots_10_io_out_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_10_out_uop_lrs2 = slots_10_io_out_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_10_out_uop_lrs1 = slots_10_io_out_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_10_out_uop_ldst = slots_10_io_out_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_ldst_is_rs1 = slots_10_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_flush_on_commit = slots_10_io_out_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_is_unique = slots_10_io_out_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_is_sys_pc2epc = slots_10_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_uses_stq = slots_10_io_out_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_uses_ldq = slots_10_io_out_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_is_amo = slots_10_io_out_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_is_fencei = slots_10_io_out_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_is_fence = slots_10_io_out_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_mem_signed = slots_10_io_out_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_10_out_uop_mem_size = slots_10_io_out_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_10_out_uop_mem_cmd = slots_10_io_out_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_bypassable = slots_10_io_out_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] issue_slots_10_out_uop_exc_cause = slots_10_io_out_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_exception = slots_10_io_out_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_10_out_uop_stale_pdst = slots_10_io_out_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_ppred_busy = slots_10_io_out_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_prs3_busy = slots_10_io_out_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_prs2_busy = slots_10_io_out_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_prs1_busy = slots_10_io_out_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_10_out_uop_ppred = slots_10_io_out_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_10_out_uop_prs3 = slots_10_io_out_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_10_out_uop_prs2 = slots_10_io_out_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_10_out_uop_prs1 = slots_10_io_out_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_10_out_uop_pdst = slots_10_io_out_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_10_out_uop_rxq_idx = slots_10_io_out_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_10_out_uop_stq_idx = slots_10_io_out_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_10_out_uop_ldq_idx = slots_10_io_out_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_10_out_uop_rob_idx = slots_10_io_out_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_10_out_uop_csr_addr = slots_10_io_out_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] issue_slots_10_out_uop_imm_packed = slots_10_io_out_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_taken = slots_10_io_out_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_10_out_uop_pc_lob = slots_10_io_out_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_edge_inst = slots_10_io_out_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_10_out_uop_ftq_idx = slots_10_io_out_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_10_out_uop_br_tag = slots_10_io_out_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_10_out_uop_br_mask = slots_10_io_out_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_is_sfb = slots_10_io_out_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_is_jal = slots_10_io_out_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_is_jalr = slots_10_io_out_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_is_br = slots_10_io_out_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_iw_p2_poisoned = slots_10_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_iw_p1_poisoned = slots_10_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_10_out_uop_iw_state = slots_10_io_out_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_ctrl_is_std = slots_10_io_out_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_ctrl_is_sta = slots_10_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_ctrl_is_load = slots_10_io_out_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_10_out_uop_ctrl_csr_cmd = slots_10_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_ctrl_fcn_dw = slots_10_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_10_out_uop_ctrl_op_fcn = slots_10_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_10_out_uop_ctrl_imm_sel = slots_10_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_10_out_uop_ctrl_op2_sel = slots_10_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_10_out_uop_ctrl_op1_sel = slots_10_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_10_out_uop_ctrl_br_type = slots_10_io_out_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_10_out_uop_fu_code = slots_10_io_out_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_10_out_uop_iq_type = slots_10_io_out_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] issue_slots_10_out_uop_debug_pc = slots_10_io_out_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_10_out_uop_is_rvc = slots_10_io_out_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_10_out_uop_debug_inst = slots_10_io_out_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_10_out_uop_inst = slots_10_io_out_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] issue_slots_10_out_uop_uopc = slots_10_io_out_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_8_clear = _GEN_25[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_1476 = _GEN_29[1:0] == 2'h1 & issue_slots_10_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_11_will_be_valid = slots_11_io_will_be_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_in_uop_valid = _GEN_31[1:0] == 2'h2 ? issue_slots_11_will_be_valid : _GEN_1476; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_11_out_uop_debug_tsrc = slots_11_io_out_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_11_out_uop_debug_fsrc = slots_11_io_out_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_bp_xcpt_if = slots_11_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_bp_debug_if = slots_11_io_out_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_xcpt_ma_if = slots_11_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_xcpt_ae_if = slots_11_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_xcpt_pf_if = slots_11_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_fp_single = slots_11_io_out_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_fp_val = slots_11_io_out_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_frs3_en = slots_11_io_out_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_11_out_uop_lrs2_rtype = slots_11_io_out_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_11_out_uop_lrs1_rtype = slots_11_io_out_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_11_out_uop_dst_rtype = slots_11_io_out_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_ldst_val = slots_11_io_out_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_out_uop_lrs3 = slots_11_io_out_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_out_uop_lrs2 = slots_11_io_out_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_out_uop_lrs1 = slots_11_io_out_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_out_uop_ldst = slots_11_io_out_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_ldst_is_rs1 = slots_11_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_flush_on_commit = slots_11_io_out_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_is_unique = slots_11_io_out_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_is_sys_pc2epc = slots_11_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_uses_stq = slots_11_io_out_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_uses_ldq = slots_11_io_out_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_is_amo = slots_11_io_out_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_is_fencei = slots_11_io_out_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_is_fence = slots_11_io_out_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_mem_signed = slots_11_io_out_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_11_out_uop_mem_size = slots_11_io_out_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_11_out_uop_mem_cmd = slots_11_io_out_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_bypassable = slots_11_io_out_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] issue_slots_11_out_uop_exc_cause = slots_11_io_out_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_exception = slots_11_io_out_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_out_uop_stale_pdst = slots_11_io_out_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_ppred_busy = slots_11_io_out_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_prs3_busy = slots_11_io_out_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_prs2_busy = slots_11_io_out_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_prs1_busy = slots_11_io_out_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_11_out_uop_ppred = slots_11_io_out_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_out_uop_prs3 = slots_11_io_out_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_out_uop_prs2 = slots_11_io_out_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_out_uop_prs1 = slots_11_io_out_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_out_uop_pdst = slots_11_io_out_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_11_out_uop_rxq_idx = slots_11_io_out_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_11_out_uop_stq_idx = slots_11_io_out_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_11_out_uop_ldq_idx = slots_11_io_out_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_out_uop_rob_idx = slots_11_io_out_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_11_out_uop_csr_addr = slots_11_io_out_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] issue_slots_11_out_uop_imm_packed = slots_11_io_out_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_taken = slots_11_io_out_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_out_uop_pc_lob = slots_11_io_out_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_edge_inst = slots_11_io_out_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_11_out_uop_ftq_idx = slots_11_io_out_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_11_out_uop_br_tag = slots_11_io_out_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_11_out_uop_br_mask = slots_11_io_out_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_is_sfb = slots_11_io_out_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_is_jal = slots_11_io_out_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_is_jalr = slots_11_io_out_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_is_br = slots_11_io_out_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_iw_p2_poisoned = slots_11_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_iw_p1_poisoned = slots_11_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_11_out_uop_iw_state = slots_11_io_out_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_ctrl_is_std = slots_11_io_out_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_ctrl_is_sta = slots_11_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_ctrl_is_load = slots_11_io_out_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_11_out_uop_ctrl_csr_cmd = slots_11_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_ctrl_fcn_dw = slots_11_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_11_out_uop_ctrl_op_fcn = slots_11_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_11_out_uop_ctrl_imm_sel = slots_11_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_11_out_uop_ctrl_op2_sel = slots_11_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_11_out_uop_ctrl_op1_sel = slots_11_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_11_out_uop_ctrl_br_type = slots_11_io_out_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [9:0] issue_slots_11_out_uop_fu_code = slots_11_io_out_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_11_out_uop_iq_type = slots_11_io_out_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] issue_slots_11_out_uop_debug_pc = slots_11_io_out_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_out_uop_is_rvc = slots_11_io_out_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_11_out_uop_debug_inst = slots_11_io_out_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_11_out_uop_inst = slots_11_io_out_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] issue_slots_11_out_uop_uopc = slots_11_io_out_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_9_clear = _GEN_27[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_1636 = _GEN_31[1:0] == 2'h1 & issue_slots_11_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_10_in_uop_valid = _GEN_33[1:0] == 2'h2 ? will_be_valid_12 : _GEN_1636; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire  issue_slots_10_clear = _GEN_29[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_1796 = _GEN_33[1:0] == 2'h1 & will_be_valid_12; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_11_in_uop_valid = _GEN_35[1:0] == 2'h2 ? will_be_valid_13 : _GEN_1796; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire  issue_slots_11_clear = _GEN_31[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  issue_slots_0_will_be_valid = slots_0_io_will_be_valid; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  will_be_available_0 = ~issue_slots_0_will_be_valid & ~issue_slots_0_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_1 = (~issue_slots_1_will_be_valid | issue_slots_1_clear) & ~issue_slots_1_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_2 = (~issue_slots_2_will_be_valid | issue_slots_2_clear) & ~issue_slots_2_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_3 = (~issue_slots_3_will_be_valid | issue_slots_3_clear) & ~issue_slots_3_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_4 = (~issue_slots_4_will_be_valid | issue_slots_4_clear) & ~issue_slots_4_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_5 = (~issue_slots_5_will_be_valid | issue_slots_5_clear) & ~issue_slots_5_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_6 = (~issue_slots_6_will_be_valid | issue_slots_6_clear) & ~issue_slots_6_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_7 = (~issue_slots_7_will_be_valid | issue_slots_7_clear) & ~issue_slots_7_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_8 = (~issue_slots_8_will_be_valid | issue_slots_8_clear) & ~issue_slots_8_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_9 = (~issue_slots_9_will_be_valid | issue_slots_9_clear) & ~issue_slots_9_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_10 = (~issue_slots_10_will_be_valid | issue_slots_10_clear) & ~issue_slots_10_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_11 = (~issue_slots_11_will_be_valid | issue_slots_11_clear) & ~issue_slots_11_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire [1:0] _T_247 = will_be_available_1 + will_be_available_2; // @[Bitwise.scala 47:55]
  wire [1:0] _GEN_2935 = {{1'd0}, will_be_available_0}; // @[Bitwise.scala 47:55]
  wire [2:0] _T_249 = _GEN_2935 + _T_247; // @[Bitwise.scala 47:55]
  wire [1:0] _T_251 = will_be_available_4 + will_be_available_5; // @[Bitwise.scala 47:55]
  wire [1:0] _GEN_2936 = {{1'd0}, will_be_available_3}; // @[Bitwise.scala 47:55]
  wire [2:0] _T_253 = _GEN_2936 + _T_251; // @[Bitwise.scala 47:55]
  wire [2:0] _T_255 = _T_249[1:0] + _T_253[1:0]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_257 = will_be_available_7 + will_be_available_8; // @[Bitwise.scala 47:55]
  wire [1:0] _GEN_2937 = {{1'd0}, will_be_available_6}; // @[Bitwise.scala 47:55]
  wire [2:0] _T_259 = _GEN_2937 + _T_257; // @[Bitwise.scala 47:55]
  wire [1:0] _T_261 = will_be_available_10 + will_be_available_11; // @[Bitwise.scala 47:55]
  wire [1:0] _GEN_2938 = {{1'd0}, will_be_available_9}; // @[Bitwise.scala 47:55]
  wire [2:0] _T_263 = _GEN_2938 + _T_261; // @[Bitwise.scala 47:55]
  wire [2:0] _T_265 = _T_259[1:0] + _T_263[1:0]; // @[Bitwise.scala 47:55]
  wire [3:0] num_available = _T_255 + _T_265; // @[Bitwise.scala 47:55]
  reg  REG; // @[issue-unit-age-ordered.scala 87:36]
  reg  REG_1; // @[issue-unit-age-ordered.scala 87:36]
  wire [1:0] issue_slots_0_uop_debug_tsrc = slots_0_io_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_1957 = _T_279 ? issue_slots_0_uop_debug_tsrc : 2'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_0_uop_debug_fsrc = slots_0_io_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_1958 = _T_279 ? issue_slots_0_uop_debug_fsrc : 2'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_bp_xcpt_if = slots_0_io_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1959 = _T_279 & issue_slots_0_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_bp_debug_if = slots_0_io_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1960 = _T_279 & issue_slots_0_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_xcpt_ma_if = slots_0_io_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1961 = _T_279 & issue_slots_0_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_xcpt_ae_if = slots_0_io_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1962 = _T_279 & issue_slots_0_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_xcpt_pf_if = slots_0_io_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1963 = _T_279 & issue_slots_0_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_fp_single = slots_0_io_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1964 = _T_279 & issue_slots_0_uop_fp_single; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_fp_val = slots_0_io_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1965 = _T_279 & issue_slots_0_uop_fp_val; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_frs3_en = slots_0_io_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1966 = _T_279 & issue_slots_0_uop_frs3_en; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_0_uop_lrs2_rtype = slots_0_io_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_1967 = _T_279 ? issue_slots_0_uop_lrs2_rtype : 2'h2; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 102:31]
  wire [1:0] issue_slots_0_uop_lrs1_rtype = slots_0_io_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_1968 = _T_279 ? issue_slots_0_uop_lrs1_rtype : 2'h2; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 101:31]
  wire [1:0] issue_slots_0_uop_dst_rtype = slots_0_io_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_1969 = _T_279 ? issue_slots_0_uop_dst_rtype : 2'h2; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_ldst_val = slots_0_io_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1970 = _T_279 & issue_slots_0_uop_ldst_val; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_lrs3 = slots_0_io_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_1971 = _T_279 ? issue_slots_0_uop_lrs3 : 6'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_lrs2 = slots_0_io_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_1972 = _T_279 ? issue_slots_0_uop_lrs2 : 6'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_lrs1 = slots_0_io_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_1973 = _T_279 ? issue_slots_0_uop_lrs1 : 6'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_ldst = slots_0_io_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_1974 = _T_279 ? issue_slots_0_uop_ldst : 6'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_ldst_is_rs1 = slots_0_io_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1975 = _T_279 & issue_slots_0_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_flush_on_commit = slots_0_io_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1976 = _T_279 & issue_slots_0_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_unique = slots_0_io_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1977 = _T_279 & issue_slots_0_uop_is_unique; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_sys_pc2epc = slots_0_io_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1978 = _T_279 & issue_slots_0_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_uses_stq = slots_0_io_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1979 = _T_279 & issue_slots_0_uop_uses_stq; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_uses_ldq = slots_0_io_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1980 = _T_279 & issue_slots_0_uop_uses_ldq; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_amo = slots_0_io_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1981 = _T_279 & issue_slots_0_uop_is_amo; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_fencei = slots_0_io_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1982 = _T_279 & issue_slots_0_uop_is_fencei; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_fence = slots_0_io_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1983 = _T_279 & issue_slots_0_uop_is_fence; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_mem_signed = slots_0_io_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1984 = _T_279 & issue_slots_0_uop_mem_signed; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_0_uop_mem_size = slots_0_io_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_1985 = _T_279 ? issue_slots_0_uop_mem_size : 2'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [4:0] issue_slots_0_uop_mem_cmd = slots_0_io_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_1986 = _T_279 ? issue_slots_0_uop_mem_cmd : 5'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_bypassable = slots_0_io_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1987 = _T_279 & issue_slots_0_uop_bypassable; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [63:0] issue_slots_0_uop_exc_cause = slots_0_io_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] _GEN_1988 = _T_279 ? issue_slots_0_uop_exc_cause : 64'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_exception = slots_0_io_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1989 = _T_279 & issue_slots_0_uop_exception; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_stale_pdst = slots_0_io_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_1990 = _T_279 ? issue_slots_0_uop_stale_pdst : 6'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_ppred_busy = slots_0_io_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1991 = _T_279 & issue_slots_0_uop_ppred_busy; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_prs3_busy = slots_0_io_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1992 = _T_279 & issue_slots_0_uop_prs3_busy; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_prs2_busy = slots_0_io_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1993 = _T_279 & issue_slots_0_uop_prs2_busy; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_prs1_busy = slots_0_io_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_1994 = _T_279 & issue_slots_0_uop_prs1_busy; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [4:0] issue_slots_0_uop_ppred = slots_0_io_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_1995 = _T_279 ? issue_slots_0_uop_ppred : 5'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_prs3 = slots_0_io_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_1996 = _T_279 ? issue_slots_0_uop_prs3 : 6'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 100:25]
  wire [5:0] issue_slots_0_uop_prs2 = slots_0_io_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_1997 = _T_279 ? issue_slots_0_uop_prs2 : 6'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 99:25]
  wire [5:0] issue_slots_0_uop_prs1 = slots_0_io_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_1998 = _T_279 ? issue_slots_0_uop_prs1 : 6'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 98:25]
  wire [5:0] issue_slots_0_uop_pdst = slots_0_io_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_1999 = _T_279 ? issue_slots_0_uop_pdst : 6'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_0_uop_rxq_idx = slots_0_io_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2000 = _T_279 ? issue_slots_0_uop_rxq_idx : 2'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] issue_slots_0_uop_stq_idx = slots_0_io_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2001 = _T_279 ? issue_slots_0_uop_stq_idx : 4'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] issue_slots_0_uop_ldq_idx = slots_0_io_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2002 = _T_279 ? issue_slots_0_uop_ldq_idx : 4'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_rob_idx = slots_0_io_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2003 = _T_279 ? issue_slots_0_uop_rob_idx : 6'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [11:0] issue_slots_0_uop_csr_addr = slots_0_io_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2004 = _T_279 ? issue_slots_0_uop_csr_addr : 12'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [19:0] issue_slots_0_uop_imm_packed = slots_0_io_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] _GEN_2005 = _T_279 ? issue_slots_0_uop_imm_packed : 20'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_taken = slots_0_io_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2006 = _T_279 & issue_slots_0_uop_taken; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_pc_lob = slots_0_io_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2007 = _T_279 ? issue_slots_0_uop_pc_lob : 6'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_edge_inst = slots_0_io_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2008 = _T_279 & issue_slots_0_uop_edge_inst; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [4:0] issue_slots_0_uop_ftq_idx = slots_0_io_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2009 = _T_279 ? issue_slots_0_uop_ftq_idx : 5'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] issue_slots_0_uop_br_tag = slots_0_io_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2010 = _T_279 ? issue_slots_0_uop_br_tag : 4'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [11:0] issue_slots_0_uop_br_mask = slots_0_io_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2011 = _T_279 ? issue_slots_0_uop_br_mask : 12'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_sfb = slots_0_io_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2012 = _T_279 & issue_slots_0_uop_is_sfb; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_jal = slots_0_io_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2013 = _T_279 & issue_slots_0_uop_is_jal; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_jalr = slots_0_io_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2014 = _T_279 & issue_slots_0_uop_is_jalr; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_br = slots_0_io_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2015 = _T_279 & issue_slots_0_uop_is_br; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_iw_p2_poisoned = slots_0_io_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2016 = _T_279 & issue_slots_0_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_iw_p1_poisoned = slots_0_io_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2017 = _T_279 & issue_slots_0_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_0_uop_iw_state = slots_0_io_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2018 = _T_279 ? issue_slots_0_uop_iw_state : 2'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_ctrl_is_std = slots_0_io_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2019 = _T_279 & issue_slots_0_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_ctrl_is_sta = slots_0_io_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2020 = _T_279 & issue_slots_0_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_ctrl_is_load = slots_0_io_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2021 = _T_279 & issue_slots_0_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [2:0] issue_slots_0_uop_ctrl_csr_cmd = slots_0_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2022 = _T_279 ? issue_slots_0_uop_ctrl_csr_cmd : 3'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_ctrl_fcn_dw = slots_0_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2023 = _T_279 & issue_slots_0_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] issue_slots_0_uop_ctrl_op_fcn = slots_0_io_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2024 = _T_279 ? issue_slots_0_uop_ctrl_op_fcn : 4'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [2:0] issue_slots_0_uop_ctrl_imm_sel = slots_0_io_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2025 = _T_279 ? issue_slots_0_uop_ctrl_imm_sel : 3'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [2:0] issue_slots_0_uop_ctrl_op2_sel = slots_0_io_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2026 = _T_279 ? issue_slots_0_uop_ctrl_op2_sel : 3'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_0_uop_ctrl_op1_sel = slots_0_io_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2027 = _T_279 ? issue_slots_0_uop_ctrl_op1_sel : 2'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] issue_slots_0_uop_ctrl_br_type = slots_0_io_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2028 = _T_279 ? issue_slots_0_uop_ctrl_br_type : 4'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [9:0] _GEN_2029 = _T_279 ? issue_slots_0_uop_fu_code : 10'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [2:0] issue_slots_0_uop_iq_type = slots_0_io_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2030 = _T_279 ? issue_slots_0_uop_iq_type : 3'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [39:0] issue_slots_0_uop_debug_pc = slots_0_io_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] _GEN_2031 = _T_279 ? issue_slots_0_uop_debug_pc : 40'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_rvc = slots_0_io_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2032 = _T_279 & issue_slots_0_uop_is_rvc; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [31:0] issue_slots_0_uop_debug_inst = slots_0_io_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2033 = _T_279 ? issue_slots_0_uop_debug_inst : 32'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [31:0] issue_slots_0_uop_inst = slots_0_io_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2034 = _T_279 ? issue_slots_0_uop_inst : 32'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [6:0] issue_slots_0_uop_uopc = slots_0_io_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] _GEN_2035 = _T_279 ? issue_slots_0_uop_uopc : 7'h0; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_1_uop_debug_tsrc = slots_1_io_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2038 = issue_slots_1_grant ? issue_slots_1_uop_debug_tsrc : _GEN_1957; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_1_uop_debug_fsrc = slots_1_io_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2039 = issue_slots_1_grant ? issue_slots_1_uop_debug_fsrc : _GEN_1958; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_bp_xcpt_if = slots_1_io_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2040 = issue_slots_1_grant ? issue_slots_1_uop_bp_xcpt_if : _GEN_1959; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_bp_debug_if = slots_1_io_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2041 = issue_slots_1_grant ? issue_slots_1_uop_bp_debug_if : _GEN_1960; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_xcpt_ma_if = slots_1_io_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2042 = issue_slots_1_grant ? issue_slots_1_uop_xcpt_ma_if : _GEN_1961; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_xcpt_ae_if = slots_1_io_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2043 = issue_slots_1_grant ? issue_slots_1_uop_xcpt_ae_if : _GEN_1962; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_xcpt_pf_if = slots_1_io_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2044 = issue_slots_1_grant ? issue_slots_1_uop_xcpt_pf_if : _GEN_1963; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_fp_single = slots_1_io_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2045 = issue_slots_1_grant ? issue_slots_1_uop_fp_single : _GEN_1964; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_fp_val = slots_1_io_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2046 = issue_slots_1_grant ? issue_slots_1_uop_fp_val : _GEN_1965; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_frs3_en = slots_1_io_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2047 = issue_slots_1_grant ? issue_slots_1_uop_frs3_en : _GEN_1966; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_1_uop_lrs2_rtype = slots_1_io_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2048 = issue_slots_1_grant ? issue_slots_1_uop_lrs2_rtype : _GEN_1967; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_1_uop_lrs1_rtype = slots_1_io_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2049 = issue_slots_1_grant ? issue_slots_1_uop_lrs1_rtype : _GEN_1968; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_1_uop_dst_rtype = slots_1_io_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2050 = issue_slots_1_grant ? issue_slots_1_uop_dst_rtype : _GEN_1969; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_ldst_val = slots_1_io_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2051 = issue_slots_1_grant ? issue_slots_1_uop_ldst_val : _GEN_1970; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_1_uop_lrs3 = slots_1_io_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2052 = issue_slots_1_grant ? issue_slots_1_uop_lrs3 : _GEN_1971; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_1_uop_lrs2 = slots_1_io_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2053 = issue_slots_1_grant ? issue_slots_1_uop_lrs2 : _GEN_1972; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_1_uop_lrs1 = slots_1_io_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2054 = issue_slots_1_grant ? issue_slots_1_uop_lrs1 : _GEN_1973; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_1_uop_ldst = slots_1_io_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2055 = issue_slots_1_grant ? issue_slots_1_uop_ldst : _GEN_1974; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_ldst_is_rs1 = slots_1_io_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2056 = issue_slots_1_grant ? issue_slots_1_uop_ldst_is_rs1 : _GEN_1975; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_flush_on_commit = slots_1_io_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2057 = issue_slots_1_grant ? issue_slots_1_uop_flush_on_commit : _GEN_1976; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_is_unique = slots_1_io_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2058 = issue_slots_1_grant ? issue_slots_1_uop_is_unique : _GEN_1977; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_is_sys_pc2epc = slots_1_io_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2059 = issue_slots_1_grant ? issue_slots_1_uop_is_sys_pc2epc : _GEN_1978; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_uses_stq = slots_1_io_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2060 = issue_slots_1_grant ? issue_slots_1_uop_uses_stq : _GEN_1979; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_uses_ldq = slots_1_io_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2061 = issue_slots_1_grant ? issue_slots_1_uop_uses_ldq : _GEN_1980; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_is_amo = slots_1_io_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2062 = issue_slots_1_grant ? issue_slots_1_uop_is_amo : _GEN_1981; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_is_fencei = slots_1_io_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2063 = issue_slots_1_grant ? issue_slots_1_uop_is_fencei : _GEN_1982; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_is_fence = slots_1_io_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2064 = issue_slots_1_grant ? issue_slots_1_uop_is_fence : _GEN_1983; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_mem_signed = slots_1_io_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2065 = issue_slots_1_grant ? issue_slots_1_uop_mem_signed : _GEN_1984; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_1_uop_mem_size = slots_1_io_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2066 = issue_slots_1_grant ? issue_slots_1_uop_mem_size : _GEN_1985; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_1_uop_mem_cmd = slots_1_io_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2067 = issue_slots_1_grant ? issue_slots_1_uop_mem_cmd : _GEN_1986; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_bypassable = slots_1_io_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2068 = issue_slots_1_grant ? issue_slots_1_uop_bypassable : _GEN_1987; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [63:0] issue_slots_1_uop_exc_cause = slots_1_io_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] _GEN_2069 = issue_slots_1_grant ? issue_slots_1_uop_exc_cause : _GEN_1988; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_exception = slots_1_io_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2070 = issue_slots_1_grant ? issue_slots_1_uop_exception : _GEN_1989; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_1_uop_stale_pdst = slots_1_io_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2071 = issue_slots_1_grant ? issue_slots_1_uop_stale_pdst : _GEN_1990; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_ppred_busy = slots_1_io_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2072 = issue_slots_1_grant ? issue_slots_1_uop_ppred_busy : _GEN_1991; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_prs3_busy = slots_1_io_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2073 = issue_slots_1_grant ? issue_slots_1_uop_prs3_busy : _GEN_1992; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_prs2_busy = slots_1_io_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2074 = issue_slots_1_grant ? issue_slots_1_uop_prs2_busy : _GEN_1993; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_prs1_busy = slots_1_io_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2075 = issue_slots_1_grant ? issue_slots_1_uop_prs1_busy : _GEN_1994; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_1_uop_ppred = slots_1_io_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2076 = issue_slots_1_grant ? issue_slots_1_uop_ppred : _GEN_1995; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_1_uop_prs3 = slots_1_io_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2077 = issue_slots_1_grant ? issue_slots_1_uop_prs3 : _GEN_1996; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_1_uop_prs2 = slots_1_io_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2078 = issue_slots_1_grant ? issue_slots_1_uop_prs2 : _GEN_1997; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_1_uop_prs1 = slots_1_io_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2079 = issue_slots_1_grant ? issue_slots_1_uop_prs1 : _GEN_1998; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_1_uop_pdst = slots_1_io_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2080 = issue_slots_1_grant ? issue_slots_1_uop_pdst : _GEN_1999; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_1_uop_rxq_idx = slots_1_io_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2081 = issue_slots_1_grant ? issue_slots_1_uop_rxq_idx : _GEN_2000; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_1_uop_stq_idx = slots_1_io_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2082 = issue_slots_1_grant ? issue_slots_1_uop_stq_idx : _GEN_2001; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_1_uop_ldq_idx = slots_1_io_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2083 = issue_slots_1_grant ? issue_slots_1_uop_ldq_idx : _GEN_2002; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_1_uop_rob_idx = slots_1_io_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2084 = issue_slots_1_grant ? issue_slots_1_uop_rob_idx : _GEN_2003; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [11:0] issue_slots_1_uop_csr_addr = slots_1_io_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2085 = issue_slots_1_grant ? issue_slots_1_uop_csr_addr : _GEN_2004; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [19:0] issue_slots_1_uop_imm_packed = slots_1_io_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] _GEN_2086 = issue_slots_1_grant ? issue_slots_1_uop_imm_packed : _GEN_2005; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_taken = slots_1_io_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2087 = issue_slots_1_grant ? issue_slots_1_uop_taken : _GEN_2006; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_1_uop_pc_lob = slots_1_io_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2088 = issue_slots_1_grant ? issue_slots_1_uop_pc_lob : _GEN_2007; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_edge_inst = slots_1_io_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2089 = issue_slots_1_grant ? issue_slots_1_uop_edge_inst : _GEN_2008; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_1_uop_ftq_idx = slots_1_io_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2090 = issue_slots_1_grant ? issue_slots_1_uop_ftq_idx : _GEN_2009; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_1_uop_br_tag = slots_1_io_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2091 = issue_slots_1_grant ? issue_slots_1_uop_br_tag : _GEN_2010; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [11:0] issue_slots_1_uop_br_mask = slots_1_io_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2092 = issue_slots_1_grant ? issue_slots_1_uop_br_mask : _GEN_2011; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_is_sfb = slots_1_io_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2093 = issue_slots_1_grant ? issue_slots_1_uop_is_sfb : _GEN_2012; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_is_jal = slots_1_io_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2094 = issue_slots_1_grant ? issue_slots_1_uop_is_jal : _GEN_2013; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_is_jalr = slots_1_io_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2095 = issue_slots_1_grant ? issue_slots_1_uop_is_jalr : _GEN_2014; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_is_br = slots_1_io_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2096 = issue_slots_1_grant ? issue_slots_1_uop_is_br : _GEN_2015; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_iw_p2_poisoned = slots_1_io_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2097 = issue_slots_1_grant ? issue_slots_1_uop_iw_p2_poisoned : _GEN_2016; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_iw_p1_poisoned = slots_1_io_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2098 = issue_slots_1_grant ? issue_slots_1_uop_iw_p1_poisoned : _GEN_2017; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_1_uop_iw_state = slots_1_io_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2099 = issue_slots_1_grant ? issue_slots_1_uop_iw_state : _GEN_2018; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_ctrl_is_std = slots_1_io_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2100 = issue_slots_1_grant ? issue_slots_1_uop_ctrl_is_std : _GEN_2019; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_ctrl_is_sta = slots_1_io_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2101 = issue_slots_1_grant ? issue_slots_1_uop_ctrl_is_sta : _GEN_2020; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_ctrl_is_load = slots_1_io_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2102 = issue_slots_1_grant ? issue_slots_1_uop_ctrl_is_load : _GEN_2021; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_1_uop_ctrl_csr_cmd = slots_1_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2103 = issue_slots_1_grant ? issue_slots_1_uop_ctrl_csr_cmd : _GEN_2022; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_ctrl_fcn_dw = slots_1_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2104 = issue_slots_1_grant ? issue_slots_1_uop_ctrl_fcn_dw : _GEN_2023; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_1_uop_ctrl_op_fcn = slots_1_io_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2105 = issue_slots_1_grant ? issue_slots_1_uop_ctrl_op_fcn : _GEN_2024; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_1_uop_ctrl_imm_sel = slots_1_io_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2106 = issue_slots_1_grant ? issue_slots_1_uop_ctrl_imm_sel : _GEN_2025; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_1_uop_ctrl_op2_sel = slots_1_io_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2107 = issue_slots_1_grant ? issue_slots_1_uop_ctrl_op2_sel : _GEN_2026; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_1_uop_ctrl_op1_sel = slots_1_io_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2108 = issue_slots_1_grant ? issue_slots_1_uop_ctrl_op1_sel : _GEN_2027; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_1_uop_ctrl_br_type = slots_1_io_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2109 = issue_slots_1_grant ? issue_slots_1_uop_ctrl_br_type : _GEN_2028; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [9:0] _GEN_2110 = issue_slots_1_grant ? issue_slots_1_uop_fu_code : _GEN_2029; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_1_uop_iq_type = slots_1_io_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2111 = issue_slots_1_grant ? issue_slots_1_uop_iq_type : _GEN_2030; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [39:0] issue_slots_1_uop_debug_pc = slots_1_io_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] _GEN_2112 = issue_slots_1_grant ? issue_slots_1_uop_debug_pc : _GEN_2031; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_1_uop_is_rvc = slots_1_io_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2113 = issue_slots_1_grant ? issue_slots_1_uop_is_rvc : _GEN_2032; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [31:0] issue_slots_1_uop_debug_inst = slots_1_io_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2114 = issue_slots_1_grant ? issue_slots_1_uop_debug_inst : _GEN_2033; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [31:0] issue_slots_1_uop_inst = slots_1_io_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2115 = issue_slots_1_grant ? issue_slots_1_uop_inst : _GEN_2034; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [6:0] issue_slots_1_uop_uopc = slots_1_io_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] _GEN_2116 = issue_slots_1_grant ? issue_slots_1_uop_uopc : _GEN_2035; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_2_uop_debug_tsrc = slots_2_io_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2119 = issue_slots_2_grant ? issue_slots_2_uop_debug_tsrc : _GEN_2038; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_2_uop_debug_fsrc = slots_2_io_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2120 = issue_slots_2_grant ? issue_slots_2_uop_debug_fsrc : _GEN_2039; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_bp_xcpt_if = slots_2_io_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2121 = issue_slots_2_grant ? issue_slots_2_uop_bp_xcpt_if : _GEN_2040; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_bp_debug_if = slots_2_io_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2122 = issue_slots_2_grant ? issue_slots_2_uop_bp_debug_if : _GEN_2041; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_xcpt_ma_if = slots_2_io_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2123 = issue_slots_2_grant ? issue_slots_2_uop_xcpt_ma_if : _GEN_2042; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_xcpt_ae_if = slots_2_io_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2124 = issue_slots_2_grant ? issue_slots_2_uop_xcpt_ae_if : _GEN_2043; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_xcpt_pf_if = slots_2_io_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2125 = issue_slots_2_grant ? issue_slots_2_uop_xcpt_pf_if : _GEN_2044; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_fp_single = slots_2_io_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2126 = issue_slots_2_grant ? issue_slots_2_uop_fp_single : _GEN_2045; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_fp_val = slots_2_io_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2127 = issue_slots_2_grant ? issue_slots_2_uop_fp_val : _GEN_2046; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_frs3_en = slots_2_io_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2128 = issue_slots_2_grant ? issue_slots_2_uop_frs3_en : _GEN_2047; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_2_uop_lrs2_rtype = slots_2_io_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2129 = issue_slots_2_grant ? issue_slots_2_uop_lrs2_rtype : _GEN_2048; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_2_uop_lrs1_rtype = slots_2_io_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2130 = issue_slots_2_grant ? issue_slots_2_uop_lrs1_rtype : _GEN_2049; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_2_uop_dst_rtype = slots_2_io_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2131 = issue_slots_2_grant ? issue_slots_2_uop_dst_rtype : _GEN_2050; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_ldst_val = slots_2_io_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2132 = issue_slots_2_grant ? issue_slots_2_uop_ldst_val : _GEN_2051; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_2_uop_lrs3 = slots_2_io_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2133 = issue_slots_2_grant ? issue_slots_2_uop_lrs3 : _GEN_2052; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_2_uop_lrs2 = slots_2_io_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2134 = issue_slots_2_grant ? issue_slots_2_uop_lrs2 : _GEN_2053; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_2_uop_lrs1 = slots_2_io_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2135 = issue_slots_2_grant ? issue_slots_2_uop_lrs1 : _GEN_2054; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_2_uop_ldst = slots_2_io_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2136 = issue_slots_2_grant ? issue_slots_2_uop_ldst : _GEN_2055; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_ldst_is_rs1 = slots_2_io_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2137 = issue_slots_2_grant ? issue_slots_2_uop_ldst_is_rs1 : _GEN_2056; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_flush_on_commit = slots_2_io_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2138 = issue_slots_2_grant ? issue_slots_2_uop_flush_on_commit : _GEN_2057; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_is_unique = slots_2_io_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2139 = issue_slots_2_grant ? issue_slots_2_uop_is_unique : _GEN_2058; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_is_sys_pc2epc = slots_2_io_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2140 = issue_slots_2_grant ? issue_slots_2_uop_is_sys_pc2epc : _GEN_2059; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_uses_stq = slots_2_io_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2141 = issue_slots_2_grant ? issue_slots_2_uop_uses_stq : _GEN_2060; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_uses_ldq = slots_2_io_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2142 = issue_slots_2_grant ? issue_slots_2_uop_uses_ldq : _GEN_2061; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_is_amo = slots_2_io_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2143 = issue_slots_2_grant ? issue_slots_2_uop_is_amo : _GEN_2062; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_is_fencei = slots_2_io_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2144 = issue_slots_2_grant ? issue_slots_2_uop_is_fencei : _GEN_2063; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_is_fence = slots_2_io_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2145 = issue_slots_2_grant ? issue_slots_2_uop_is_fence : _GEN_2064; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_mem_signed = slots_2_io_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2146 = issue_slots_2_grant ? issue_slots_2_uop_mem_signed : _GEN_2065; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_2_uop_mem_size = slots_2_io_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2147 = issue_slots_2_grant ? issue_slots_2_uop_mem_size : _GEN_2066; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_2_uop_mem_cmd = slots_2_io_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2148 = issue_slots_2_grant ? issue_slots_2_uop_mem_cmd : _GEN_2067; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_bypassable = slots_2_io_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2149 = issue_slots_2_grant ? issue_slots_2_uop_bypassable : _GEN_2068; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [63:0] issue_slots_2_uop_exc_cause = slots_2_io_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] _GEN_2150 = issue_slots_2_grant ? issue_slots_2_uop_exc_cause : _GEN_2069; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_exception = slots_2_io_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2151 = issue_slots_2_grant ? issue_slots_2_uop_exception : _GEN_2070; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_2_uop_stale_pdst = slots_2_io_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2152 = issue_slots_2_grant ? issue_slots_2_uop_stale_pdst : _GEN_2071; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_ppred_busy = slots_2_io_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2153 = issue_slots_2_grant ? issue_slots_2_uop_ppred_busy : _GEN_2072; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_prs3_busy = slots_2_io_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2154 = issue_slots_2_grant ? issue_slots_2_uop_prs3_busy : _GEN_2073; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_prs2_busy = slots_2_io_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2155 = issue_slots_2_grant ? issue_slots_2_uop_prs2_busy : _GEN_2074; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_prs1_busy = slots_2_io_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2156 = issue_slots_2_grant ? issue_slots_2_uop_prs1_busy : _GEN_2075; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_2_uop_ppred = slots_2_io_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2157 = issue_slots_2_grant ? issue_slots_2_uop_ppred : _GEN_2076; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_2_uop_prs3 = slots_2_io_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2158 = issue_slots_2_grant ? issue_slots_2_uop_prs3 : _GEN_2077; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_2_uop_prs2 = slots_2_io_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2159 = issue_slots_2_grant ? issue_slots_2_uop_prs2 : _GEN_2078; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_2_uop_prs1 = slots_2_io_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2160 = issue_slots_2_grant ? issue_slots_2_uop_prs1 : _GEN_2079; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_2_uop_pdst = slots_2_io_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2161 = issue_slots_2_grant ? issue_slots_2_uop_pdst : _GEN_2080; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_2_uop_rxq_idx = slots_2_io_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2162 = issue_slots_2_grant ? issue_slots_2_uop_rxq_idx : _GEN_2081; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_2_uop_stq_idx = slots_2_io_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2163 = issue_slots_2_grant ? issue_slots_2_uop_stq_idx : _GEN_2082; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_2_uop_ldq_idx = slots_2_io_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2164 = issue_slots_2_grant ? issue_slots_2_uop_ldq_idx : _GEN_2083; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_2_uop_rob_idx = slots_2_io_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2165 = issue_slots_2_grant ? issue_slots_2_uop_rob_idx : _GEN_2084; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [11:0] issue_slots_2_uop_csr_addr = slots_2_io_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2166 = issue_slots_2_grant ? issue_slots_2_uop_csr_addr : _GEN_2085; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [19:0] issue_slots_2_uop_imm_packed = slots_2_io_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] _GEN_2167 = issue_slots_2_grant ? issue_slots_2_uop_imm_packed : _GEN_2086; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_taken = slots_2_io_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2168 = issue_slots_2_grant ? issue_slots_2_uop_taken : _GEN_2087; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_2_uop_pc_lob = slots_2_io_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2169 = issue_slots_2_grant ? issue_slots_2_uop_pc_lob : _GEN_2088; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_edge_inst = slots_2_io_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2170 = issue_slots_2_grant ? issue_slots_2_uop_edge_inst : _GEN_2089; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_2_uop_ftq_idx = slots_2_io_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2171 = issue_slots_2_grant ? issue_slots_2_uop_ftq_idx : _GEN_2090; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_2_uop_br_tag = slots_2_io_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2172 = issue_slots_2_grant ? issue_slots_2_uop_br_tag : _GEN_2091; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [11:0] issue_slots_2_uop_br_mask = slots_2_io_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2173 = issue_slots_2_grant ? issue_slots_2_uop_br_mask : _GEN_2092; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_is_sfb = slots_2_io_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2174 = issue_slots_2_grant ? issue_slots_2_uop_is_sfb : _GEN_2093; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_is_jal = slots_2_io_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2175 = issue_slots_2_grant ? issue_slots_2_uop_is_jal : _GEN_2094; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_is_jalr = slots_2_io_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2176 = issue_slots_2_grant ? issue_slots_2_uop_is_jalr : _GEN_2095; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_is_br = slots_2_io_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2177 = issue_slots_2_grant ? issue_slots_2_uop_is_br : _GEN_2096; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_iw_p2_poisoned = slots_2_io_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2178 = issue_slots_2_grant ? issue_slots_2_uop_iw_p2_poisoned : _GEN_2097; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_iw_p1_poisoned = slots_2_io_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2179 = issue_slots_2_grant ? issue_slots_2_uop_iw_p1_poisoned : _GEN_2098; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_2_uop_iw_state = slots_2_io_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2180 = issue_slots_2_grant ? issue_slots_2_uop_iw_state : _GEN_2099; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_ctrl_is_std = slots_2_io_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2181 = issue_slots_2_grant ? issue_slots_2_uop_ctrl_is_std : _GEN_2100; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_ctrl_is_sta = slots_2_io_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2182 = issue_slots_2_grant ? issue_slots_2_uop_ctrl_is_sta : _GEN_2101; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_ctrl_is_load = slots_2_io_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2183 = issue_slots_2_grant ? issue_slots_2_uop_ctrl_is_load : _GEN_2102; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_2_uop_ctrl_csr_cmd = slots_2_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2184 = issue_slots_2_grant ? issue_slots_2_uop_ctrl_csr_cmd : _GEN_2103; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_ctrl_fcn_dw = slots_2_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2185 = issue_slots_2_grant ? issue_slots_2_uop_ctrl_fcn_dw : _GEN_2104; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_2_uop_ctrl_op_fcn = slots_2_io_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2186 = issue_slots_2_grant ? issue_slots_2_uop_ctrl_op_fcn : _GEN_2105; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_2_uop_ctrl_imm_sel = slots_2_io_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2187 = issue_slots_2_grant ? issue_slots_2_uop_ctrl_imm_sel : _GEN_2106; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_2_uop_ctrl_op2_sel = slots_2_io_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2188 = issue_slots_2_grant ? issue_slots_2_uop_ctrl_op2_sel : _GEN_2107; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_2_uop_ctrl_op1_sel = slots_2_io_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2189 = issue_slots_2_grant ? issue_slots_2_uop_ctrl_op1_sel : _GEN_2108; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_2_uop_ctrl_br_type = slots_2_io_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2190 = issue_slots_2_grant ? issue_slots_2_uop_ctrl_br_type : _GEN_2109; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [9:0] _GEN_2191 = issue_slots_2_grant ? issue_slots_2_uop_fu_code : _GEN_2110; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_2_uop_iq_type = slots_2_io_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2192 = issue_slots_2_grant ? issue_slots_2_uop_iq_type : _GEN_2111; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [39:0] issue_slots_2_uop_debug_pc = slots_2_io_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] _GEN_2193 = issue_slots_2_grant ? issue_slots_2_uop_debug_pc : _GEN_2112; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_2_uop_is_rvc = slots_2_io_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2194 = issue_slots_2_grant ? issue_slots_2_uop_is_rvc : _GEN_2113; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [31:0] issue_slots_2_uop_debug_inst = slots_2_io_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2195 = issue_slots_2_grant ? issue_slots_2_uop_debug_inst : _GEN_2114; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [31:0] issue_slots_2_uop_inst = slots_2_io_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2196 = issue_slots_2_grant ? issue_slots_2_uop_inst : _GEN_2115; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [6:0] issue_slots_2_uop_uopc = slots_2_io_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] _GEN_2197 = issue_slots_2_grant ? issue_slots_2_uop_uopc : _GEN_2116; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_3_uop_debug_tsrc = slots_3_io_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2200 = issue_slots_3_grant ? issue_slots_3_uop_debug_tsrc : _GEN_2119; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_3_uop_debug_fsrc = slots_3_io_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2201 = issue_slots_3_grant ? issue_slots_3_uop_debug_fsrc : _GEN_2120; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_bp_xcpt_if = slots_3_io_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2202 = issue_slots_3_grant ? issue_slots_3_uop_bp_xcpt_if : _GEN_2121; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_bp_debug_if = slots_3_io_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2203 = issue_slots_3_grant ? issue_slots_3_uop_bp_debug_if : _GEN_2122; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_xcpt_ma_if = slots_3_io_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2204 = issue_slots_3_grant ? issue_slots_3_uop_xcpt_ma_if : _GEN_2123; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_xcpt_ae_if = slots_3_io_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2205 = issue_slots_3_grant ? issue_slots_3_uop_xcpt_ae_if : _GEN_2124; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_xcpt_pf_if = slots_3_io_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2206 = issue_slots_3_grant ? issue_slots_3_uop_xcpt_pf_if : _GEN_2125; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_fp_single = slots_3_io_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2207 = issue_slots_3_grant ? issue_slots_3_uop_fp_single : _GEN_2126; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_fp_val = slots_3_io_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2208 = issue_slots_3_grant ? issue_slots_3_uop_fp_val : _GEN_2127; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_frs3_en = slots_3_io_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2209 = issue_slots_3_grant ? issue_slots_3_uop_frs3_en : _GEN_2128; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_3_uop_lrs2_rtype = slots_3_io_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2210 = issue_slots_3_grant ? issue_slots_3_uop_lrs2_rtype : _GEN_2129; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_3_uop_lrs1_rtype = slots_3_io_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2211 = issue_slots_3_grant ? issue_slots_3_uop_lrs1_rtype : _GEN_2130; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_3_uop_dst_rtype = slots_3_io_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2212 = issue_slots_3_grant ? issue_slots_3_uop_dst_rtype : _GEN_2131; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_ldst_val = slots_3_io_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2213 = issue_slots_3_grant ? issue_slots_3_uop_ldst_val : _GEN_2132; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_3_uop_lrs3 = slots_3_io_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2214 = issue_slots_3_grant ? issue_slots_3_uop_lrs3 : _GEN_2133; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_3_uop_lrs2 = slots_3_io_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2215 = issue_slots_3_grant ? issue_slots_3_uop_lrs2 : _GEN_2134; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_3_uop_lrs1 = slots_3_io_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2216 = issue_slots_3_grant ? issue_slots_3_uop_lrs1 : _GEN_2135; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_3_uop_ldst = slots_3_io_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2217 = issue_slots_3_grant ? issue_slots_3_uop_ldst : _GEN_2136; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_ldst_is_rs1 = slots_3_io_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2218 = issue_slots_3_grant ? issue_slots_3_uop_ldst_is_rs1 : _GEN_2137; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_flush_on_commit = slots_3_io_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2219 = issue_slots_3_grant ? issue_slots_3_uop_flush_on_commit : _GEN_2138; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_is_unique = slots_3_io_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2220 = issue_slots_3_grant ? issue_slots_3_uop_is_unique : _GEN_2139; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_is_sys_pc2epc = slots_3_io_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2221 = issue_slots_3_grant ? issue_slots_3_uop_is_sys_pc2epc : _GEN_2140; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_uses_stq = slots_3_io_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2222 = issue_slots_3_grant ? issue_slots_3_uop_uses_stq : _GEN_2141; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_uses_ldq = slots_3_io_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2223 = issue_slots_3_grant ? issue_slots_3_uop_uses_ldq : _GEN_2142; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_is_amo = slots_3_io_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2224 = issue_slots_3_grant ? issue_slots_3_uop_is_amo : _GEN_2143; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_is_fencei = slots_3_io_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2225 = issue_slots_3_grant ? issue_slots_3_uop_is_fencei : _GEN_2144; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_is_fence = slots_3_io_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2226 = issue_slots_3_grant ? issue_slots_3_uop_is_fence : _GEN_2145; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_mem_signed = slots_3_io_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2227 = issue_slots_3_grant ? issue_slots_3_uop_mem_signed : _GEN_2146; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_3_uop_mem_size = slots_3_io_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2228 = issue_slots_3_grant ? issue_slots_3_uop_mem_size : _GEN_2147; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_3_uop_mem_cmd = slots_3_io_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2229 = issue_slots_3_grant ? issue_slots_3_uop_mem_cmd : _GEN_2148; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_bypassable = slots_3_io_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2230 = issue_slots_3_grant ? issue_slots_3_uop_bypassable : _GEN_2149; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [63:0] issue_slots_3_uop_exc_cause = slots_3_io_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] _GEN_2231 = issue_slots_3_grant ? issue_slots_3_uop_exc_cause : _GEN_2150; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_exception = slots_3_io_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2232 = issue_slots_3_grant ? issue_slots_3_uop_exception : _GEN_2151; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_3_uop_stale_pdst = slots_3_io_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2233 = issue_slots_3_grant ? issue_slots_3_uop_stale_pdst : _GEN_2152; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_ppred_busy = slots_3_io_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2234 = issue_slots_3_grant ? issue_slots_3_uop_ppred_busy : _GEN_2153; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_prs3_busy = slots_3_io_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2235 = issue_slots_3_grant ? issue_slots_3_uop_prs3_busy : _GEN_2154; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_prs2_busy = slots_3_io_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2236 = issue_slots_3_grant ? issue_slots_3_uop_prs2_busy : _GEN_2155; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_prs1_busy = slots_3_io_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2237 = issue_slots_3_grant ? issue_slots_3_uop_prs1_busy : _GEN_2156; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_3_uop_ppred = slots_3_io_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2238 = issue_slots_3_grant ? issue_slots_3_uop_ppred : _GEN_2157; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_3_uop_prs3 = slots_3_io_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2239 = issue_slots_3_grant ? issue_slots_3_uop_prs3 : _GEN_2158; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_3_uop_prs2 = slots_3_io_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2240 = issue_slots_3_grant ? issue_slots_3_uop_prs2 : _GEN_2159; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_3_uop_prs1 = slots_3_io_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2241 = issue_slots_3_grant ? issue_slots_3_uop_prs1 : _GEN_2160; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_3_uop_pdst = slots_3_io_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2242 = issue_slots_3_grant ? issue_slots_3_uop_pdst : _GEN_2161; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_3_uop_rxq_idx = slots_3_io_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2243 = issue_slots_3_grant ? issue_slots_3_uop_rxq_idx : _GEN_2162; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_3_uop_stq_idx = slots_3_io_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2244 = issue_slots_3_grant ? issue_slots_3_uop_stq_idx : _GEN_2163; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_3_uop_ldq_idx = slots_3_io_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2245 = issue_slots_3_grant ? issue_slots_3_uop_ldq_idx : _GEN_2164; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_3_uop_rob_idx = slots_3_io_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2246 = issue_slots_3_grant ? issue_slots_3_uop_rob_idx : _GEN_2165; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [11:0] issue_slots_3_uop_csr_addr = slots_3_io_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2247 = issue_slots_3_grant ? issue_slots_3_uop_csr_addr : _GEN_2166; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [19:0] issue_slots_3_uop_imm_packed = slots_3_io_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] _GEN_2248 = issue_slots_3_grant ? issue_slots_3_uop_imm_packed : _GEN_2167; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_taken = slots_3_io_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2249 = issue_slots_3_grant ? issue_slots_3_uop_taken : _GEN_2168; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_3_uop_pc_lob = slots_3_io_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2250 = issue_slots_3_grant ? issue_slots_3_uop_pc_lob : _GEN_2169; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_edge_inst = slots_3_io_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2251 = issue_slots_3_grant ? issue_slots_3_uop_edge_inst : _GEN_2170; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_3_uop_ftq_idx = slots_3_io_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2252 = issue_slots_3_grant ? issue_slots_3_uop_ftq_idx : _GEN_2171; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_3_uop_br_tag = slots_3_io_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2253 = issue_slots_3_grant ? issue_slots_3_uop_br_tag : _GEN_2172; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [11:0] issue_slots_3_uop_br_mask = slots_3_io_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2254 = issue_slots_3_grant ? issue_slots_3_uop_br_mask : _GEN_2173; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_is_sfb = slots_3_io_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2255 = issue_slots_3_grant ? issue_slots_3_uop_is_sfb : _GEN_2174; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_is_jal = slots_3_io_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2256 = issue_slots_3_grant ? issue_slots_3_uop_is_jal : _GEN_2175; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_is_jalr = slots_3_io_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2257 = issue_slots_3_grant ? issue_slots_3_uop_is_jalr : _GEN_2176; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_is_br = slots_3_io_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2258 = issue_slots_3_grant ? issue_slots_3_uop_is_br : _GEN_2177; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_iw_p2_poisoned = slots_3_io_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2259 = issue_slots_3_grant ? issue_slots_3_uop_iw_p2_poisoned : _GEN_2178; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_iw_p1_poisoned = slots_3_io_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2260 = issue_slots_3_grant ? issue_slots_3_uop_iw_p1_poisoned : _GEN_2179; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_3_uop_iw_state = slots_3_io_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2261 = issue_slots_3_grant ? issue_slots_3_uop_iw_state : _GEN_2180; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_ctrl_is_std = slots_3_io_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2262 = issue_slots_3_grant ? issue_slots_3_uop_ctrl_is_std : _GEN_2181; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_ctrl_is_sta = slots_3_io_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2263 = issue_slots_3_grant ? issue_slots_3_uop_ctrl_is_sta : _GEN_2182; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_ctrl_is_load = slots_3_io_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2264 = issue_slots_3_grant ? issue_slots_3_uop_ctrl_is_load : _GEN_2183; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_3_uop_ctrl_csr_cmd = slots_3_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2265 = issue_slots_3_grant ? issue_slots_3_uop_ctrl_csr_cmd : _GEN_2184; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_ctrl_fcn_dw = slots_3_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2266 = issue_slots_3_grant ? issue_slots_3_uop_ctrl_fcn_dw : _GEN_2185; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_3_uop_ctrl_op_fcn = slots_3_io_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2267 = issue_slots_3_grant ? issue_slots_3_uop_ctrl_op_fcn : _GEN_2186; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_3_uop_ctrl_imm_sel = slots_3_io_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2268 = issue_slots_3_grant ? issue_slots_3_uop_ctrl_imm_sel : _GEN_2187; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_3_uop_ctrl_op2_sel = slots_3_io_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2269 = issue_slots_3_grant ? issue_slots_3_uop_ctrl_op2_sel : _GEN_2188; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_3_uop_ctrl_op1_sel = slots_3_io_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2270 = issue_slots_3_grant ? issue_slots_3_uop_ctrl_op1_sel : _GEN_2189; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_3_uop_ctrl_br_type = slots_3_io_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2271 = issue_slots_3_grant ? issue_slots_3_uop_ctrl_br_type : _GEN_2190; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [9:0] _GEN_2272 = issue_slots_3_grant ? issue_slots_3_uop_fu_code : _GEN_2191; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_3_uop_iq_type = slots_3_io_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2273 = issue_slots_3_grant ? issue_slots_3_uop_iq_type : _GEN_2192; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [39:0] issue_slots_3_uop_debug_pc = slots_3_io_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] _GEN_2274 = issue_slots_3_grant ? issue_slots_3_uop_debug_pc : _GEN_2193; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_3_uop_is_rvc = slots_3_io_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2275 = issue_slots_3_grant ? issue_slots_3_uop_is_rvc : _GEN_2194; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [31:0] issue_slots_3_uop_debug_inst = slots_3_io_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2276 = issue_slots_3_grant ? issue_slots_3_uop_debug_inst : _GEN_2195; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [31:0] issue_slots_3_uop_inst = slots_3_io_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2277 = issue_slots_3_grant ? issue_slots_3_uop_inst : _GEN_2196; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [6:0] issue_slots_3_uop_uopc = slots_3_io_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] _GEN_2278 = issue_slots_3_grant ? issue_slots_3_uop_uopc : _GEN_2197; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_4_uop_debug_tsrc = slots_4_io_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2281 = issue_slots_4_grant ? issue_slots_4_uop_debug_tsrc : _GEN_2200; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_4_uop_debug_fsrc = slots_4_io_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2282 = issue_slots_4_grant ? issue_slots_4_uop_debug_fsrc : _GEN_2201; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_bp_xcpt_if = slots_4_io_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2283 = issue_slots_4_grant ? issue_slots_4_uop_bp_xcpt_if : _GEN_2202; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_bp_debug_if = slots_4_io_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2284 = issue_slots_4_grant ? issue_slots_4_uop_bp_debug_if : _GEN_2203; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_xcpt_ma_if = slots_4_io_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2285 = issue_slots_4_grant ? issue_slots_4_uop_xcpt_ma_if : _GEN_2204; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_xcpt_ae_if = slots_4_io_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2286 = issue_slots_4_grant ? issue_slots_4_uop_xcpt_ae_if : _GEN_2205; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_xcpt_pf_if = slots_4_io_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2287 = issue_slots_4_grant ? issue_slots_4_uop_xcpt_pf_if : _GEN_2206; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_fp_single = slots_4_io_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2288 = issue_slots_4_grant ? issue_slots_4_uop_fp_single : _GEN_2207; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_fp_val = slots_4_io_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2289 = issue_slots_4_grant ? issue_slots_4_uop_fp_val : _GEN_2208; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_frs3_en = slots_4_io_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2290 = issue_slots_4_grant ? issue_slots_4_uop_frs3_en : _GEN_2209; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_4_uop_lrs2_rtype = slots_4_io_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2291 = issue_slots_4_grant ? issue_slots_4_uop_lrs2_rtype : _GEN_2210; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_4_uop_lrs1_rtype = slots_4_io_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2292 = issue_slots_4_grant ? issue_slots_4_uop_lrs1_rtype : _GEN_2211; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_4_uop_dst_rtype = slots_4_io_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2293 = issue_slots_4_grant ? issue_slots_4_uop_dst_rtype : _GEN_2212; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_ldst_val = slots_4_io_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2294 = issue_slots_4_grant ? issue_slots_4_uop_ldst_val : _GEN_2213; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_4_uop_lrs3 = slots_4_io_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2295 = issue_slots_4_grant ? issue_slots_4_uop_lrs3 : _GEN_2214; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_4_uop_lrs2 = slots_4_io_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2296 = issue_slots_4_grant ? issue_slots_4_uop_lrs2 : _GEN_2215; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_4_uop_lrs1 = slots_4_io_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2297 = issue_slots_4_grant ? issue_slots_4_uop_lrs1 : _GEN_2216; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_4_uop_ldst = slots_4_io_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2298 = issue_slots_4_grant ? issue_slots_4_uop_ldst : _GEN_2217; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_ldst_is_rs1 = slots_4_io_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2299 = issue_slots_4_grant ? issue_slots_4_uop_ldst_is_rs1 : _GEN_2218; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_flush_on_commit = slots_4_io_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2300 = issue_slots_4_grant ? issue_slots_4_uop_flush_on_commit : _GEN_2219; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_is_unique = slots_4_io_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2301 = issue_slots_4_grant ? issue_slots_4_uop_is_unique : _GEN_2220; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_is_sys_pc2epc = slots_4_io_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2302 = issue_slots_4_grant ? issue_slots_4_uop_is_sys_pc2epc : _GEN_2221; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_uses_stq = slots_4_io_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2303 = issue_slots_4_grant ? issue_slots_4_uop_uses_stq : _GEN_2222; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_uses_ldq = slots_4_io_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2304 = issue_slots_4_grant ? issue_slots_4_uop_uses_ldq : _GEN_2223; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_is_amo = slots_4_io_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2305 = issue_slots_4_grant ? issue_slots_4_uop_is_amo : _GEN_2224; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_is_fencei = slots_4_io_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2306 = issue_slots_4_grant ? issue_slots_4_uop_is_fencei : _GEN_2225; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_is_fence = slots_4_io_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2307 = issue_slots_4_grant ? issue_slots_4_uop_is_fence : _GEN_2226; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_mem_signed = slots_4_io_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2308 = issue_slots_4_grant ? issue_slots_4_uop_mem_signed : _GEN_2227; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_4_uop_mem_size = slots_4_io_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2309 = issue_slots_4_grant ? issue_slots_4_uop_mem_size : _GEN_2228; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_4_uop_mem_cmd = slots_4_io_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2310 = issue_slots_4_grant ? issue_slots_4_uop_mem_cmd : _GEN_2229; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_bypassable = slots_4_io_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2311 = issue_slots_4_grant ? issue_slots_4_uop_bypassable : _GEN_2230; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [63:0] issue_slots_4_uop_exc_cause = slots_4_io_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] _GEN_2312 = issue_slots_4_grant ? issue_slots_4_uop_exc_cause : _GEN_2231; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_exception = slots_4_io_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2313 = issue_slots_4_grant ? issue_slots_4_uop_exception : _GEN_2232; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_4_uop_stale_pdst = slots_4_io_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2314 = issue_slots_4_grant ? issue_slots_4_uop_stale_pdst : _GEN_2233; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_ppred_busy = slots_4_io_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2315 = issue_slots_4_grant ? issue_slots_4_uop_ppred_busy : _GEN_2234; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_prs3_busy = slots_4_io_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2316 = issue_slots_4_grant ? issue_slots_4_uop_prs3_busy : _GEN_2235; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_prs2_busy = slots_4_io_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2317 = issue_slots_4_grant ? issue_slots_4_uop_prs2_busy : _GEN_2236; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_prs1_busy = slots_4_io_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2318 = issue_slots_4_grant ? issue_slots_4_uop_prs1_busy : _GEN_2237; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_4_uop_ppred = slots_4_io_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2319 = issue_slots_4_grant ? issue_slots_4_uop_ppred : _GEN_2238; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_4_uop_prs3 = slots_4_io_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2320 = issue_slots_4_grant ? issue_slots_4_uop_prs3 : _GEN_2239; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_4_uop_prs2 = slots_4_io_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2321 = issue_slots_4_grant ? issue_slots_4_uop_prs2 : _GEN_2240; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_4_uop_prs1 = slots_4_io_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2322 = issue_slots_4_grant ? issue_slots_4_uop_prs1 : _GEN_2241; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_4_uop_pdst = slots_4_io_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2323 = issue_slots_4_grant ? issue_slots_4_uop_pdst : _GEN_2242; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_4_uop_rxq_idx = slots_4_io_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2324 = issue_slots_4_grant ? issue_slots_4_uop_rxq_idx : _GEN_2243; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_4_uop_stq_idx = slots_4_io_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2325 = issue_slots_4_grant ? issue_slots_4_uop_stq_idx : _GEN_2244; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_4_uop_ldq_idx = slots_4_io_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2326 = issue_slots_4_grant ? issue_slots_4_uop_ldq_idx : _GEN_2245; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_4_uop_rob_idx = slots_4_io_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2327 = issue_slots_4_grant ? issue_slots_4_uop_rob_idx : _GEN_2246; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [11:0] issue_slots_4_uop_csr_addr = slots_4_io_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2328 = issue_slots_4_grant ? issue_slots_4_uop_csr_addr : _GEN_2247; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [19:0] issue_slots_4_uop_imm_packed = slots_4_io_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] _GEN_2329 = issue_slots_4_grant ? issue_slots_4_uop_imm_packed : _GEN_2248; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_taken = slots_4_io_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2330 = issue_slots_4_grant ? issue_slots_4_uop_taken : _GEN_2249; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_4_uop_pc_lob = slots_4_io_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2331 = issue_slots_4_grant ? issue_slots_4_uop_pc_lob : _GEN_2250; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_edge_inst = slots_4_io_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2332 = issue_slots_4_grant ? issue_slots_4_uop_edge_inst : _GEN_2251; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_4_uop_ftq_idx = slots_4_io_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2333 = issue_slots_4_grant ? issue_slots_4_uop_ftq_idx : _GEN_2252; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_4_uop_br_tag = slots_4_io_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2334 = issue_slots_4_grant ? issue_slots_4_uop_br_tag : _GEN_2253; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [11:0] issue_slots_4_uop_br_mask = slots_4_io_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2335 = issue_slots_4_grant ? issue_slots_4_uop_br_mask : _GEN_2254; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_is_sfb = slots_4_io_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2336 = issue_slots_4_grant ? issue_slots_4_uop_is_sfb : _GEN_2255; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_is_jal = slots_4_io_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2337 = issue_slots_4_grant ? issue_slots_4_uop_is_jal : _GEN_2256; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_is_jalr = slots_4_io_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2338 = issue_slots_4_grant ? issue_slots_4_uop_is_jalr : _GEN_2257; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_is_br = slots_4_io_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2339 = issue_slots_4_grant ? issue_slots_4_uop_is_br : _GEN_2258; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_iw_p2_poisoned = slots_4_io_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2340 = issue_slots_4_grant ? issue_slots_4_uop_iw_p2_poisoned : _GEN_2259; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_iw_p1_poisoned = slots_4_io_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2341 = issue_slots_4_grant ? issue_slots_4_uop_iw_p1_poisoned : _GEN_2260; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_4_uop_iw_state = slots_4_io_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2342 = issue_slots_4_grant ? issue_slots_4_uop_iw_state : _GEN_2261; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_ctrl_is_std = slots_4_io_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2343 = issue_slots_4_grant ? issue_slots_4_uop_ctrl_is_std : _GEN_2262; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_ctrl_is_sta = slots_4_io_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2344 = issue_slots_4_grant ? issue_slots_4_uop_ctrl_is_sta : _GEN_2263; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_ctrl_is_load = slots_4_io_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2345 = issue_slots_4_grant ? issue_slots_4_uop_ctrl_is_load : _GEN_2264; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_4_uop_ctrl_csr_cmd = slots_4_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2346 = issue_slots_4_grant ? issue_slots_4_uop_ctrl_csr_cmd : _GEN_2265; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_ctrl_fcn_dw = slots_4_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2347 = issue_slots_4_grant ? issue_slots_4_uop_ctrl_fcn_dw : _GEN_2266; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_4_uop_ctrl_op_fcn = slots_4_io_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2348 = issue_slots_4_grant ? issue_slots_4_uop_ctrl_op_fcn : _GEN_2267; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_4_uop_ctrl_imm_sel = slots_4_io_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2349 = issue_slots_4_grant ? issue_slots_4_uop_ctrl_imm_sel : _GEN_2268; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_4_uop_ctrl_op2_sel = slots_4_io_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2350 = issue_slots_4_grant ? issue_slots_4_uop_ctrl_op2_sel : _GEN_2269; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_4_uop_ctrl_op1_sel = slots_4_io_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2351 = issue_slots_4_grant ? issue_slots_4_uop_ctrl_op1_sel : _GEN_2270; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_4_uop_ctrl_br_type = slots_4_io_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2352 = issue_slots_4_grant ? issue_slots_4_uop_ctrl_br_type : _GEN_2271; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [9:0] _GEN_2353 = issue_slots_4_grant ? issue_slots_4_uop_fu_code : _GEN_2272; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_4_uop_iq_type = slots_4_io_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2354 = issue_slots_4_grant ? issue_slots_4_uop_iq_type : _GEN_2273; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [39:0] issue_slots_4_uop_debug_pc = slots_4_io_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] _GEN_2355 = issue_slots_4_grant ? issue_slots_4_uop_debug_pc : _GEN_2274; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_4_uop_is_rvc = slots_4_io_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2356 = issue_slots_4_grant ? issue_slots_4_uop_is_rvc : _GEN_2275; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [31:0] issue_slots_4_uop_debug_inst = slots_4_io_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2357 = issue_slots_4_grant ? issue_slots_4_uop_debug_inst : _GEN_2276; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [31:0] issue_slots_4_uop_inst = slots_4_io_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2358 = issue_slots_4_grant ? issue_slots_4_uop_inst : _GEN_2277; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [6:0] issue_slots_4_uop_uopc = slots_4_io_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] _GEN_2359 = issue_slots_4_grant ? issue_slots_4_uop_uopc : _GEN_2278; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_5_uop_debug_tsrc = slots_5_io_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2362 = issue_slots_5_grant ? issue_slots_5_uop_debug_tsrc : _GEN_2281; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_5_uop_debug_fsrc = slots_5_io_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2363 = issue_slots_5_grant ? issue_slots_5_uop_debug_fsrc : _GEN_2282; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_bp_xcpt_if = slots_5_io_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2364 = issue_slots_5_grant ? issue_slots_5_uop_bp_xcpt_if : _GEN_2283; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_bp_debug_if = slots_5_io_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2365 = issue_slots_5_grant ? issue_slots_5_uop_bp_debug_if : _GEN_2284; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_xcpt_ma_if = slots_5_io_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2366 = issue_slots_5_grant ? issue_slots_5_uop_xcpt_ma_if : _GEN_2285; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_xcpt_ae_if = slots_5_io_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2367 = issue_slots_5_grant ? issue_slots_5_uop_xcpt_ae_if : _GEN_2286; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_xcpt_pf_if = slots_5_io_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2368 = issue_slots_5_grant ? issue_slots_5_uop_xcpt_pf_if : _GEN_2287; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_fp_single = slots_5_io_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2369 = issue_slots_5_grant ? issue_slots_5_uop_fp_single : _GEN_2288; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_fp_val = slots_5_io_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2370 = issue_slots_5_grant ? issue_slots_5_uop_fp_val : _GEN_2289; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_frs3_en = slots_5_io_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2371 = issue_slots_5_grant ? issue_slots_5_uop_frs3_en : _GEN_2290; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_5_uop_lrs2_rtype = slots_5_io_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2372 = issue_slots_5_grant ? issue_slots_5_uop_lrs2_rtype : _GEN_2291; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_5_uop_lrs1_rtype = slots_5_io_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2373 = issue_slots_5_grant ? issue_slots_5_uop_lrs1_rtype : _GEN_2292; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_5_uop_dst_rtype = slots_5_io_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2374 = issue_slots_5_grant ? issue_slots_5_uop_dst_rtype : _GEN_2293; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_ldst_val = slots_5_io_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2375 = issue_slots_5_grant ? issue_slots_5_uop_ldst_val : _GEN_2294; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_5_uop_lrs3 = slots_5_io_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2376 = issue_slots_5_grant ? issue_slots_5_uop_lrs3 : _GEN_2295; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_5_uop_lrs2 = slots_5_io_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2377 = issue_slots_5_grant ? issue_slots_5_uop_lrs2 : _GEN_2296; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_5_uop_lrs1 = slots_5_io_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2378 = issue_slots_5_grant ? issue_slots_5_uop_lrs1 : _GEN_2297; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_5_uop_ldst = slots_5_io_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2379 = issue_slots_5_grant ? issue_slots_5_uop_ldst : _GEN_2298; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_ldst_is_rs1 = slots_5_io_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2380 = issue_slots_5_grant ? issue_slots_5_uop_ldst_is_rs1 : _GEN_2299; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_flush_on_commit = slots_5_io_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2381 = issue_slots_5_grant ? issue_slots_5_uop_flush_on_commit : _GEN_2300; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_is_unique = slots_5_io_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2382 = issue_slots_5_grant ? issue_slots_5_uop_is_unique : _GEN_2301; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_is_sys_pc2epc = slots_5_io_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2383 = issue_slots_5_grant ? issue_slots_5_uop_is_sys_pc2epc : _GEN_2302; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_uses_stq = slots_5_io_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2384 = issue_slots_5_grant ? issue_slots_5_uop_uses_stq : _GEN_2303; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_uses_ldq = slots_5_io_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2385 = issue_slots_5_grant ? issue_slots_5_uop_uses_ldq : _GEN_2304; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_is_amo = slots_5_io_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2386 = issue_slots_5_grant ? issue_slots_5_uop_is_amo : _GEN_2305; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_is_fencei = slots_5_io_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2387 = issue_slots_5_grant ? issue_slots_5_uop_is_fencei : _GEN_2306; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_is_fence = slots_5_io_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2388 = issue_slots_5_grant ? issue_slots_5_uop_is_fence : _GEN_2307; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_mem_signed = slots_5_io_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2389 = issue_slots_5_grant ? issue_slots_5_uop_mem_signed : _GEN_2308; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_5_uop_mem_size = slots_5_io_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2390 = issue_slots_5_grant ? issue_slots_5_uop_mem_size : _GEN_2309; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_5_uop_mem_cmd = slots_5_io_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2391 = issue_slots_5_grant ? issue_slots_5_uop_mem_cmd : _GEN_2310; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_bypassable = slots_5_io_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2392 = issue_slots_5_grant ? issue_slots_5_uop_bypassable : _GEN_2311; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [63:0] issue_slots_5_uop_exc_cause = slots_5_io_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] _GEN_2393 = issue_slots_5_grant ? issue_slots_5_uop_exc_cause : _GEN_2312; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_exception = slots_5_io_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2394 = issue_slots_5_grant ? issue_slots_5_uop_exception : _GEN_2313; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_5_uop_stale_pdst = slots_5_io_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2395 = issue_slots_5_grant ? issue_slots_5_uop_stale_pdst : _GEN_2314; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_ppred_busy = slots_5_io_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2396 = issue_slots_5_grant ? issue_slots_5_uop_ppred_busy : _GEN_2315; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_prs3_busy = slots_5_io_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2397 = issue_slots_5_grant ? issue_slots_5_uop_prs3_busy : _GEN_2316; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_prs2_busy = slots_5_io_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2398 = issue_slots_5_grant ? issue_slots_5_uop_prs2_busy : _GEN_2317; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_prs1_busy = slots_5_io_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2399 = issue_slots_5_grant ? issue_slots_5_uop_prs1_busy : _GEN_2318; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_5_uop_ppred = slots_5_io_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2400 = issue_slots_5_grant ? issue_slots_5_uop_ppred : _GEN_2319; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_5_uop_prs3 = slots_5_io_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2401 = issue_slots_5_grant ? issue_slots_5_uop_prs3 : _GEN_2320; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_5_uop_prs2 = slots_5_io_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2402 = issue_slots_5_grant ? issue_slots_5_uop_prs2 : _GEN_2321; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_5_uop_prs1 = slots_5_io_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2403 = issue_slots_5_grant ? issue_slots_5_uop_prs1 : _GEN_2322; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_5_uop_pdst = slots_5_io_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2404 = issue_slots_5_grant ? issue_slots_5_uop_pdst : _GEN_2323; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_5_uop_rxq_idx = slots_5_io_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2405 = issue_slots_5_grant ? issue_slots_5_uop_rxq_idx : _GEN_2324; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_5_uop_stq_idx = slots_5_io_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2406 = issue_slots_5_grant ? issue_slots_5_uop_stq_idx : _GEN_2325; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_5_uop_ldq_idx = slots_5_io_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2407 = issue_slots_5_grant ? issue_slots_5_uop_ldq_idx : _GEN_2326; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_5_uop_rob_idx = slots_5_io_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2408 = issue_slots_5_grant ? issue_slots_5_uop_rob_idx : _GEN_2327; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [11:0] issue_slots_5_uop_csr_addr = slots_5_io_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2409 = issue_slots_5_grant ? issue_slots_5_uop_csr_addr : _GEN_2328; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [19:0] issue_slots_5_uop_imm_packed = slots_5_io_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] _GEN_2410 = issue_slots_5_grant ? issue_slots_5_uop_imm_packed : _GEN_2329; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_taken = slots_5_io_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2411 = issue_slots_5_grant ? issue_slots_5_uop_taken : _GEN_2330; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_5_uop_pc_lob = slots_5_io_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2412 = issue_slots_5_grant ? issue_slots_5_uop_pc_lob : _GEN_2331; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_edge_inst = slots_5_io_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2413 = issue_slots_5_grant ? issue_slots_5_uop_edge_inst : _GEN_2332; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_5_uop_ftq_idx = slots_5_io_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2414 = issue_slots_5_grant ? issue_slots_5_uop_ftq_idx : _GEN_2333; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_5_uop_br_tag = slots_5_io_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2415 = issue_slots_5_grant ? issue_slots_5_uop_br_tag : _GEN_2334; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [11:0] issue_slots_5_uop_br_mask = slots_5_io_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2416 = issue_slots_5_grant ? issue_slots_5_uop_br_mask : _GEN_2335; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_is_sfb = slots_5_io_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2417 = issue_slots_5_grant ? issue_slots_5_uop_is_sfb : _GEN_2336; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_is_jal = slots_5_io_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2418 = issue_slots_5_grant ? issue_slots_5_uop_is_jal : _GEN_2337; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_is_jalr = slots_5_io_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2419 = issue_slots_5_grant ? issue_slots_5_uop_is_jalr : _GEN_2338; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_is_br = slots_5_io_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2420 = issue_slots_5_grant ? issue_slots_5_uop_is_br : _GEN_2339; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_iw_p2_poisoned = slots_5_io_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2421 = issue_slots_5_grant ? issue_slots_5_uop_iw_p2_poisoned : _GEN_2340; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_iw_p1_poisoned = slots_5_io_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2422 = issue_slots_5_grant ? issue_slots_5_uop_iw_p1_poisoned : _GEN_2341; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_5_uop_iw_state = slots_5_io_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2423 = issue_slots_5_grant ? issue_slots_5_uop_iw_state : _GEN_2342; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_ctrl_is_std = slots_5_io_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2424 = issue_slots_5_grant ? issue_slots_5_uop_ctrl_is_std : _GEN_2343; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_ctrl_is_sta = slots_5_io_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2425 = issue_slots_5_grant ? issue_slots_5_uop_ctrl_is_sta : _GEN_2344; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_ctrl_is_load = slots_5_io_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2426 = issue_slots_5_grant ? issue_slots_5_uop_ctrl_is_load : _GEN_2345; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_5_uop_ctrl_csr_cmd = slots_5_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2427 = issue_slots_5_grant ? issue_slots_5_uop_ctrl_csr_cmd : _GEN_2346; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_ctrl_fcn_dw = slots_5_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2428 = issue_slots_5_grant ? issue_slots_5_uop_ctrl_fcn_dw : _GEN_2347; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_5_uop_ctrl_op_fcn = slots_5_io_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2429 = issue_slots_5_grant ? issue_slots_5_uop_ctrl_op_fcn : _GEN_2348; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_5_uop_ctrl_imm_sel = slots_5_io_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2430 = issue_slots_5_grant ? issue_slots_5_uop_ctrl_imm_sel : _GEN_2349; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_5_uop_ctrl_op2_sel = slots_5_io_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2431 = issue_slots_5_grant ? issue_slots_5_uop_ctrl_op2_sel : _GEN_2350; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_5_uop_ctrl_op1_sel = slots_5_io_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2432 = issue_slots_5_grant ? issue_slots_5_uop_ctrl_op1_sel : _GEN_2351; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_5_uop_ctrl_br_type = slots_5_io_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2433 = issue_slots_5_grant ? issue_slots_5_uop_ctrl_br_type : _GEN_2352; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [9:0] _GEN_2434 = issue_slots_5_grant ? issue_slots_5_uop_fu_code : _GEN_2353; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_5_uop_iq_type = slots_5_io_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2435 = issue_slots_5_grant ? issue_slots_5_uop_iq_type : _GEN_2354; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [39:0] issue_slots_5_uop_debug_pc = slots_5_io_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] _GEN_2436 = issue_slots_5_grant ? issue_slots_5_uop_debug_pc : _GEN_2355; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_5_uop_is_rvc = slots_5_io_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2437 = issue_slots_5_grant ? issue_slots_5_uop_is_rvc : _GEN_2356; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [31:0] issue_slots_5_uop_debug_inst = slots_5_io_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2438 = issue_slots_5_grant ? issue_slots_5_uop_debug_inst : _GEN_2357; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [31:0] issue_slots_5_uop_inst = slots_5_io_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2439 = issue_slots_5_grant ? issue_slots_5_uop_inst : _GEN_2358; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [6:0] issue_slots_5_uop_uopc = slots_5_io_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] _GEN_2440 = issue_slots_5_grant ? issue_slots_5_uop_uopc : _GEN_2359; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_6_uop_debug_tsrc = slots_6_io_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2443 = issue_slots_6_grant ? issue_slots_6_uop_debug_tsrc : _GEN_2362; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_6_uop_debug_fsrc = slots_6_io_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2444 = issue_slots_6_grant ? issue_slots_6_uop_debug_fsrc : _GEN_2363; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_bp_xcpt_if = slots_6_io_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2445 = issue_slots_6_grant ? issue_slots_6_uop_bp_xcpt_if : _GEN_2364; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_bp_debug_if = slots_6_io_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2446 = issue_slots_6_grant ? issue_slots_6_uop_bp_debug_if : _GEN_2365; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_xcpt_ma_if = slots_6_io_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2447 = issue_slots_6_grant ? issue_slots_6_uop_xcpt_ma_if : _GEN_2366; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_xcpt_ae_if = slots_6_io_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2448 = issue_slots_6_grant ? issue_slots_6_uop_xcpt_ae_if : _GEN_2367; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_xcpt_pf_if = slots_6_io_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2449 = issue_slots_6_grant ? issue_slots_6_uop_xcpt_pf_if : _GEN_2368; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_fp_single = slots_6_io_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2450 = issue_slots_6_grant ? issue_slots_6_uop_fp_single : _GEN_2369; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_fp_val = slots_6_io_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2451 = issue_slots_6_grant ? issue_slots_6_uop_fp_val : _GEN_2370; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_frs3_en = slots_6_io_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2452 = issue_slots_6_grant ? issue_slots_6_uop_frs3_en : _GEN_2371; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_6_uop_lrs2_rtype = slots_6_io_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2453 = issue_slots_6_grant ? issue_slots_6_uop_lrs2_rtype : _GEN_2372; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_6_uop_lrs1_rtype = slots_6_io_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2454 = issue_slots_6_grant ? issue_slots_6_uop_lrs1_rtype : _GEN_2373; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_6_uop_dst_rtype = slots_6_io_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2455 = issue_slots_6_grant ? issue_slots_6_uop_dst_rtype : _GEN_2374; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_ldst_val = slots_6_io_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2456 = issue_slots_6_grant ? issue_slots_6_uop_ldst_val : _GEN_2375; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_6_uop_lrs3 = slots_6_io_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2457 = issue_slots_6_grant ? issue_slots_6_uop_lrs3 : _GEN_2376; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_6_uop_lrs2 = slots_6_io_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2458 = issue_slots_6_grant ? issue_slots_6_uop_lrs2 : _GEN_2377; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_6_uop_lrs1 = slots_6_io_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2459 = issue_slots_6_grant ? issue_slots_6_uop_lrs1 : _GEN_2378; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_6_uop_ldst = slots_6_io_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2460 = issue_slots_6_grant ? issue_slots_6_uop_ldst : _GEN_2379; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_ldst_is_rs1 = slots_6_io_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2461 = issue_slots_6_grant ? issue_slots_6_uop_ldst_is_rs1 : _GEN_2380; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_flush_on_commit = slots_6_io_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2462 = issue_slots_6_grant ? issue_slots_6_uop_flush_on_commit : _GEN_2381; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_is_unique = slots_6_io_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2463 = issue_slots_6_grant ? issue_slots_6_uop_is_unique : _GEN_2382; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_is_sys_pc2epc = slots_6_io_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2464 = issue_slots_6_grant ? issue_slots_6_uop_is_sys_pc2epc : _GEN_2383; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_uses_stq = slots_6_io_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2465 = issue_slots_6_grant ? issue_slots_6_uop_uses_stq : _GEN_2384; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_uses_ldq = slots_6_io_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2466 = issue_slots_6_grant ? issue_slots_6_uop_uses_ldq : _GEN_2385; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_is_amo = slots_6_io_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2467 = issue_slots_6_grant ? issue_slots_6_uop_is_amo : _GEN_2386; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_is_fencei = slots_6_io_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2468 = issue_slots_6_grant ? issue_slots_6_uop_is_fencei : _GEN_2387; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_is_fence = slots_6_io_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2469 = issue_slots_6_grant ? issue_slots_6_uop_is_fence : _GEN_2388; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_mem_signed = slots_6_io_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2470 = issue_slots_6_grant ? issue_slots_6_uop_mem_signed : _GEN_2389; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_6_uop_mem_size = slots_6_io_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2471 = issue_slots_6_grant ? issue_slots_6_uop_mem_size : _GEN_2390; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_6_uop_mem_cmd = slots_6_io_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2472 = issue_slots_6_grant ? issue_slots_6_uop_mem_cmd : _GEN_2391; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_bypassable = slots_6_io_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2473 = issue_slots_6_grant ? issue_slots_6_uop_bypassable : _GEN_2392; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [63:0] issue_slots_6_uop_exc_cause = slots_6_io_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] _GEN_2474 = issue_slots_6_grant ? issue_slots_6_uop_exc_cause : _GEN_2393; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_exception = slots_6_io_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2475 = issue_slots_6_grant ? issue_slots_6_uop_exception : _GEN_2394; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_6_uop_stale_pdst = slots_6_io_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2476 = issue_slots_6_grant ? issue_slots_6_uop_stale_pdst : _GEN_2395; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_ppred_busy = slots_6_io_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2477 = issue_slots_6_grant ? issue_slots_6_uop_ppred_busy : _GEN_2396; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_prs3_busy = slots_6_io_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2478 = issue_slots_6_grant ? issue_slots_6_uop_prs3_busy : _GEN_2397; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_prs2_busy = slots_6_io_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2479 = issue_slots_6_grant ? issue_slots_6_uop_prs2_busy : _GEN_2398; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_prs1_busy = slots_6_io_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2480 = issue_slots_6_grant ? issue_slots_6_uop_prs1_busy : _GEN_2399; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_6_uop_ppred = slots_6_io_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2481 = issue_slots_6_grant ? issue_slots_6_uop_ppred : _GEN_2400; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_6_uop_prs3 = slots_6_io_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2482 = issue_slots_6_grant ? issue_slots_6_uop_prs3 : _GEN_2401; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_6_uop_prs2 = slots_6_io_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2483 = issue_slots_6_grant ? issue_slots_6_uop_prs2 : _GEN_2402; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_6_uop_prs1 = slots_6_io_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2484 = issue_slots_6_grant ? issue_slots_6_uop_prs1 : _GEN_2403; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_6_uop_pdst = slots_6_io_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2485 = issue_slots_6_grant ? issue_slots_6_uop_pdst : _GEN_2404; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_6_uop_rxq_idx = slots_6_io_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2486 = issue_slots_6_grant ? issue_slots_6_uop_rxq_idx : _GEN_2405; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_6_uop_stq_idx = slots_6_io_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2487 = issue_slots_6_grant ? issue_slots_6_uop_stq_idx : _GEN_2406; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_6_uop_ldq_idx = slots_6_io_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2488 = issue_slots_6_grant ? issue_slots_6_uop_ldq_idx : _GEN_2407; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_6_uop_rob_idx = slots_6_io_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2489 = issue_slots_6_grant ? issue_slots_6_uop_rob_idx : _GEN_2408; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [11:0] issue_slots_6_uop_csr_addr = slots_6_io_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2490 = issue_slots_6_grant ? issue_slots_6_uop_csr_addr : _GEN_2409; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [19:0] issue_slots_6_uop_imm_packed = slots_6_io_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] _GEN_2491 = issue_slots_6_grant ? issue_slots_6_uop_imm_packed : _GEN_2410; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_taken = slots_6_io_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2492 = issue_slots_6_grant ? issue_slots_6_uop_taken : _GEN_2411; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_6_uop_pc_lob = slots_6_io_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2493 = issue_slots_6_grant ? issue_slots_6_uop_pc_lob : _GEN_2412; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_edge_inst = slots_6_io_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2494 = issue_slots_6_grant ? issue_slots_6_uop_edge_inst : _GEN_2413; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_6_uop_ftq_idx = slots_6_io_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2495 = issue_slots_6_grant ? issue_slots_6_uop_ftq_idx : _GEN_2414; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_6_uop_br_tag = slots_6_io_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2496 = issue_slots_6_grant ? issue_slots_6_uop_br_tag : _GEN_2415; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [11:0] issue_slots_6_uop_br_mask = slots_6_io_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2497 = issue_slots_6_grant ? issue_slots_6_uop_br_mask : _GEN_2416; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_is_sfb = slots_6_io_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2498 = issue_slots_6_grant ? issue_slots_6_uop_is_sfb : _GEN_2417; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_is_jal = slots_6_io_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2499 = issue_slots_6_grant ? issue_slots_6_uop_is_jal : _GEN_2418; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_is_jalr = slots_6_io_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2500 = issue_slots_6_grant ? issue_slots_6_uop_is_jalr : _GEN_2419; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_is_br = slots_6_io_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2501 = issue_slots_6_grant ? issue_slots_6_uop_is_br : _GEN_2420; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_iw_p2_poisoned = slots_6_io_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2502 = issue_slots_6_grant ? issue_slots_6_uop_iw_p2_poisoned : _GEN_2421; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_iw_p1_poisoned = slots_6_io_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2503 = issue_slots_6_grant ? issue_slots_6_uop_iw_p1_poisoned : _GEN_2422; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_6_uop_iw_state = slots_6_io_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2504 = issue_slots_6_grant ? issue_slots_6_uop_iw_state : _GEN_2423; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_ctrl_is_std = slots_6_io_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2505 = issue_slots_6_grant ? issue_slots_6_uop_ctrl_is_std : _GEN_2424; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_ctrl_is_sta = slots_6_io_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2506 = issue_slots_6_grant ? issue_slots_6_uop_ctrl_is_sta : _GEN_2425; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_ctrl_is_load = slots_6_io_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2507 = issue_slots_6_grant ? issue_slots_6_uop_ctrl_is_load : _GEN_2426; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_6_uop_ctrl_csr_cmd = slots_6_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2508 = issue_slots_6_grant ? issue_slots_6_uop_ctrl_csr_cmd : _GEN_2427; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_ctrl_fcn_dw = slots_6_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2509 = issue_slots_6_grant ? issue_slots_6_uop_ctrl_fcn_dw : _GEN_2428; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_6_uop_ctrl_op_fcn = slots_6_io_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2510 = issue_slots_6_grant ? issue_slots_6_uop_ctrl_op_fcn : _GEN_2429; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_6_uop_ctrl_imm_sel = slots_6_io_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2511 = issue_slots_6_grant ? issue_slots_6_uop_ctrl_imm_sel : _GEN_2430; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_6_uop_ctrl_op2_sel = slots_6_io_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2512 = issue_slots_6_grant ? issue_slots_6_uop_ctrl_op2_sel : _GEN_2431; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_6_uop_ctrl_op1_sel = slots_6_io_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2513 = issue_slots_6_grant ? issue_slots_6_uop_ctrl_op1_sel : _GEN_2432; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_6_uop_ctrl_br_type = slots_6_io_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2514 = issue_slots_6_grant ? issue_slots_6_uop_ctrl_br_type : _GEN_2433; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [9:0] _GEN_2515 = issue_slots_6_grant ? issue_slots_6_uop_fu_code : _GEN_2434; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_6_uop_iq_type = slots_6_io_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2516 = issue_slots_6_grant ? issue_slots_6_uop_iq_type : _GEN_2435; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [39:0] issue_slots_6_uop_debug_pc = slots_6_io_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] _GEN_2517 = issue_slots_6_grant ? issue_slots_6_uop_debug_pc : _GEN_2436; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_6_uop_is_rvc = slots_6_io_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2518 = issue_slots_6_grant ? issue_slots_6_uop_is_rvc : _GEN_2437; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [31:0] issue_slots_6_uop_debug_inst = slots_6_io_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2519 = issue_slots_6_grant ? issue_slots_6_uop_debug_inst : _GEN_2438; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [31:0] issue_slots_6_uop_inst = slots_6_io_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2520 = issue_slots_6_grant ? issue_slots_6_uop_inst : _GEN_2439; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [6:0] issue_slots_6_uop_uopc = slots_6_io_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] _GEN_2521 = issue_slots_6_grant ? issue_slots_6_uop_uopc : _GEN_2440; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_7_uop_debug_tsrc = slots_7_io_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2524 = issue_slots_7_grant ? issue_slots_7_uop_debug_tsrc : _GEN_2443; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_7_uop_debug_fsrc = slots_7_io_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2525 = issue_slots_7_grant ? issue_slots_7_uop_debug_fsrc : _GEN_2444; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_bp_xcpt_if = slots_7_io_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2526 = issue_slots_7_grant ? issue_slots_7_uop_bp_xcpt_if : _GEN_2445; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_bp_debug_if = slots_7_io_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2527 = issue_slots_7_grant ? issue_slots_7_uop_bp_debug_if : _GEN_2446; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_xcpt_ma_if = slots_7_io_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2528 = issue_slots_7_grant ? issue_slots_7_uop_xcpt_ma_if : _GEN_2447; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_xcpt_ae_if = slots_7_io_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2529 = issue_slots_7_grant ? issue_slots_7_uop_xcpt_ae_if : _GEN_2448; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_xcpt_pf_if = slots_7_io_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2530 = issue_slots_7_grant ? issue_slots_7_uop_xcpt_pf_if : _GEN_2449; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_fp_single = slots_7_io_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2531 = issue_slots_7_grant ? issue_slots_7_uop_fp_single : _GEN_2450; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_fp_val = slots_7_io_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2532 = issue_slots_7_grant ? issue_slots_7_uop_fp_val : _GEN_2451; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_frs3_en = slots_7_io_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2533 = issue_slots_7_grant ? issue_slots_7_uop_frs3_en : _GEN_2452; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_7_uop_lrs2_rtype = slots_7_io_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2534 = issue_slots_7_grant ? issue_slots_7_uop_lrs2_rtype : _GEN_2453; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_7_uop_lrs1_rtype = slots_7_io_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2535 = issue_slots_7_grant ? issue_slots_7_uop_lrs1_rtype : _GEN_2454; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_7_uop_dst_rtype = slots_7_io_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2536 = issue_slots_7_grant ? issue_slots_7_uop_dst_rtype : _GEN_2455; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_ldst_val = slots_7_io_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2537 = issue_slots_7_grant ? issue_slots_7_uop_ldst_val : _GEN_2456; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_7_uop_lrs3 = slots_7_io_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2538 = issue_slots_7_grant ? issue_slots_7_uop_lrs3 : _GEN_2457; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_7_uop_lrs2 = slots_7_io_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2539 = issue_slots_7_grant ? issue_slots_7_uop_lrs2 : _GEN_2458; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_7_uop_lrs1 = slots_7_io_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2540 = issue_slots_7_grant ? issue_slots_7_uop_lrs1 : _GEN_2459; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_7_uop_ldst = slots_7_io_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2541 = issue_slots_7_grant ? issue_slots_7_uop_ldst : _GEN_2460; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_ldst_is_rs1 = slots_7_io_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2542 = issue_slots_7_grant ? issue_slots_7_uop_ldst_is_rs1 : _GEN_2461; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_flush_on_commit = slots_7_io_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2543 = issue_slots_7_grant ? issue_slots_7_uop_flush_on_commit : _GEN_2462; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_is_unique = slots_7_io_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2544 = issue_slots_7_grant ? issue_slots_7_uop_is_unique : _GEN_2463; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_is_sys_pc2epc = slots_7_io_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2545 = issue_slots_7_grant ? issue_slots_7_uop_is_sys_pc2epc : _GEN_2464; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_uses_stq = slots_7_io_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2546 = issue_slots_7_grant ? issue_slots_7_uop_uses_stq : _GEN_2465; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_uses_ldq = slots_7_io_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2547 = issue_slots_7_grant ? issue_slots_7_uop_uses_ldq : _GEN_2466; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_is_amo = slots_7_io_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2548 = issue_slots_7_grant ? issue_slots_7_uop_is_amo : _GEN_2467; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_is_fencei = slots_7_io_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2549 = issue_slots_7_grant ? issue_slots_7_uop_is_fencei : _GEN_2468; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_is_fence = slots_7_io_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2550 = issue_slots_7_grant ? issue_slots_7_uop_is_fence : _GEN_2469; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_mem_signed = slots_7_io_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2551 = issue_slots_7_grant ? issue_slots_7_uop_mem_signed : _GEN_2470; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_7_uop_mem_size = slots_7_io_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2552 = issue_slots_7_grant ? issue_slots_7_uop_mem_size : _GEN_2471; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_7_uop_mem_cmd = slots_7_io_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2553 = issue_slots_7_grant ? issue_slots_7_uop_mem_cmd : _GEN_2472; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_bypassable = slots_7_io_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2554 = issue_slots_7_grant ? issue_slots_7_uop_bypassable : _GEN_2473; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [63:0] issue_slots_7_uop_exc_cause = slots_7_io_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] _GEN_2555 = issue_slots_7_grant ? issue_slots_7_uop_exc_cause : _GEN_2474; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_exception = slots_7_io_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2556 = issue_slots_7_grant ? issue_slots_7_uop_exception : _GEN_2475; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_7_uop_stale_pdst = slots_7_io_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2557 = issue_slots_7_grant ? issue_slots_7_uop_stale_pdst : _GEN_2476; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_ppred_busy = slots_7_io_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2558 = issue_slots_7_grant ? issue_slots_7_uop_ppred_busy : _GEN_2477; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_prs3_busy = slots_7_io_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2559 = issue_slots_7_grant ? issue_slots_7_uop_prs3_busy : _GEN_2478; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_prs2_busy = slots_7_io_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2560 = issue_slots_7_grant ? issue_slots_7_uop_prs2_busy : _GEN_2479; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_prs1_busy = slots_7_io_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2561 = issue_slots_7_grant ? issue_slots_7_uop_prs1_busy : _GEN_2480; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_7_uop_ppred = slots_7_io_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2562 = issue_slots_7_grant ? issue_slots_7_uop_ppred : _GEN_2481; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_7_uop_prs3 = slots_7_io_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2563 = issue_slots_7_grant ? issue_slots_7_uop_prs3 : _GEN_2482; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_7_uop_prs2 = slots_7_io_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2564 = issue_slots_7_grant ? issue_slots_7_uop_prs2 : _GEN_2483; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_7_uop_prs1 = slots_7_io_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2565 = issue_slots_7_grant ? issue_slots_7_uop_prs1 : _GEN_2484; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_7_uop_pdst = slots_7_io_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2566 = issue_slots_7_grant ? issue_slots_7_uop_pdst : _GEN_2485; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_7_uop_rxq_idx = slots_7_io_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2567 = issue_slots_7_grant ? issue_slots_7_uop_rxq_idx : _GEN_2486; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_7_uop_stq_idx = slots_7_io_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2568 = issue_slots_7_grant ? issue_slots_7_uop_stq_idx : _GEN_2487; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_7_uop_ldq_idx = slots_7_io_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2569 = issue_slots_7_grant ? issue_slots_7_uop_ldq_idx : _GEN_2488; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_7_uop_rob_idx = slots_7_io_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2570 = issue_slots_7_grant ? issue_slots_7_uop_rob_idx : _GEN_2489; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [11:0] issue_slots_7_uop_csr_addr = slots_7_io_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2571 = issue_slots_7_grant ? issue_slots_7_uop_csr_addr : _GEN_2490; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [19:0] issue_slots_7_uop_imm_packed = slots_7_io_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] _GEN_2572 = issue_slots_7_grant ? issue_slots_7_uop_imm_packed : _GEN_2491; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_taken = slots_7_io_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2573 = issue_slots_7_grant ? issue_slots_7_uop_taken : _GEN_2492; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_7_uop_pc_lob = slots_7_io_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2574 = issue_slots_7_grant ? issue_slots_7_uop_pc_lob : _GEN_2493; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_edge_inst = slots_7_io_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2575 = issue_slots_7_grant ? issue_slots_7_uop_edge_inst : _GEN_2494; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_7_uop_ftq_idx = slots_7_io_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2576 = issue_slots_7_grant ? issue_slots_7_uop_ftq_idx : _GEN_2495; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_7_uop_br_tag = slots_7_io_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2577 = issue_slots_7_grant ? issue_slots_7_uop_br_tag : _GEN_2496; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [11:0] issue_slots_7_uop_br_mask = slots_7_io_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2578 = issue_slots_7_grant ? issue_slots_7_uop_br_mask : _GEN_2497; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_is_sfb = slots_7_io_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2579 = issue_slots_7_grant ? issue_slots_7_uop_is_sfb : _GEN_2498; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_is_jal = slots_7_io_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2580 = issue_slots_7_grant ? issue_slots_7_uop_is_jal : _GEN_2499; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_is_jalr = slots_7_io_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2581 = issue_slots_7_grant ? issue_slots_7_uop_is_jalr : _GEN_2500; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_is_br = slots_7_io_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2582 = issue_slots_7_grant ? issue_slots_7_uop_is_br : _GEN_2501; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_iw_p2_poisoned = slots_7_io_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2583 = issue_slots_7_grant ? issue_slots_7_uop_iw_p2_poisoned : _GEN_2502; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_iw_p1_poisoned = slots_7_io_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2584 = issue_slots_7_grant ? issue_slots_7_uop_iw_p1_poisoned : _GEN_2503; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_7_uop_iw_state = slots_7_io_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2585 = issue_slots_7_grant ? issue_slots_7_uop_iw_state : _GEN_2504; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_ctrl_is_std = slots_7_io_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2586 = issue_slots_7_grant ? issue_slots_7_uop_ctrl_is_std : _GEN_2505; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_ctrl_is_sta = slots_7_io_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2587 = issue_slots_7_grant ? issue_slots_7_uop_ctrl_is_sta : _GEN_2506; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_ctrl_is_load = slots_7_io_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2588 = issue_slots_7_grant ? issue_slots_7_uop_ctrl_is_load : _GEN_2507; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_7_uop_ctrl_csr_cmd = slots_7_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2589 = issue_slots_7_grant ? issue_slots_7_uop_ctrl_csr_cmd : _GEN_2508; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_ctrl_fcn_dw = slots_7_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2590 = issue_slots_7_grant ? issue_slots_7_uop_ctrl_fcn_dw : _GEN_2509; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_7_uop_ctrl_op_fcn = slots_7_io_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2591 = issue_slots_7_grant ? issue_slots_7_uop_ctrl_op_fcn : _GEN_2510; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_7_uop_ctrl_imm_sel = slots_7_io_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2592 = issue_slots_7_grant ? issue_slots_7_uop_ctrl_imm_sel : _GEN_2511; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_7_uop_ctrl_op2_sel = slots_7_io_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2593 = issue_slots_7_grant ? issue_slots_7_uop_ctrl_op2_sel : _GEN_2512; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_7_uop_ctrl_op1_sel = slots_7_io_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2594 = issue_slots_7_grant ? issue_slots_7_uop_ctrl_op1_sel : _GEN_2513; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_7_uop_ctrl_br_type = slots_7_io_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2595 = issue_slots_7_grant ? issue_slots_7_uop_ctrl_br_type : _GEN_2514; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [9:0] _GEN_2596 = issue_slots_7_grant ? issue_slots_7_uop_fu_code : _GEN_2515; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_7_uop_iq_type = slots_7_io_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2597 = issue_slots_7_grant ? issue_slots_7_uop_iq_type : _GEN_2516; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [39:0] issue_slots_7_uop_debug_pc = slots_7_io_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] _GEN_2598 = issue_slots_7_grant ? issue_slots_7_uop_debug_pc : _GEN_2517; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_7_uop_is_rvc = slots_7_io_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2599 = issue_slots_7_grant ? issue_slots_7_uop_is_rvc : _GEN_2518; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [31:0] issue_slots_7_uop_debug_inst = slots_7_io_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2600 = issue_slots_7_grant ? issue_slots_7_uop_debug_inst : _GEN_2519; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [31:0] issue_slots_7_uop_inst = slots_7_io_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2601 = issue_slots_7_grant ? issue_slots_7_uop_inst : _GEN_2520; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [6:0] issue_slots_7_uop_uopc = slots_7_io_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] _GEN_2602 = issue_slots_7_grant ? issue_slots_7_uop_uopc : _GEN_2521; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_8_uop_debug_tsrc = slots_8_io_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2605 = issue_slots_8_grant ? issue_slots_8_uop_debug_tsrc : _GEN_2524; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_8_uop_debug_fsrc = slots_8_io_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2606 = issue_slots_8_grant ? issue_slots_8_uop_debug_fsrc : _GEN_2525; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_bp_xcpt_if = slots_8_io_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2607 = issue_slots_8_grant ? issue_slots_8_uop_bp_xcpt_if : _GEN_2526; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_bp_debug_if = slots_8_io_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2608 = issue_slots_8_grant ? issue_slots_8_uop_bp_debug_if : _GEN_2527; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_xcpt_ma_if = slots_8_io_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2609 = issue_slots_8_grant ? issue_slots_8_uop_xcpt_ma_if : _GEN_2528; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_xcpt_ae_if = slots_8_io_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2610 = issue_slots_8_grant ? issue_slots_8_uop_xcpt_ae_if : _GEN_2529; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_xcpt_pf_if = slots_8_io_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2611 = issue_slots_8_grant ? issue_slots_8_uop_xcpt_pf_if : _GEN_2530; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_fp_single = slots_8_io_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2612 = issue_slots_8_grant ? issue_slots_8_uop_fp_single : _GEN_2531; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_fp_val = slots_8_io_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2613 = issue_slots_8_grant ? issue_slots_8_uop_fp_val : _GEN_2532; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_frs3_en = slots_8_io_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2614 = issue_slots_8_grant ? issue_slots_8_uop_frs3_en : _GEN_2533; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_8_uop_lrs2_rtype = slots_8_io_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2615 = issue_slots_8_grant ? issue_slots_8_uop_lrs2_rtype : _GEN_2534; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_8_uop_lrs1_rtype = slots_8_io_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2616 = issue_slots_8_grant ? issue_slots_8_uop_lrs1_rtype : _GEN_2535; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_8_uop_dst_rtype = slots_8_io_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2617 = issue_slots_8_grant ? issue_slots_8_uop_dst_rtype : _GEN_2536; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_ldst_val = slots_8_io_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2618 = issue_slots_8_grant ? issue_slots_8_uop_ldst_val : _GEN_2537; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_8_uop_lrs3 = slots_8_io_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2619 = issue_slots_8_grant ? issue_slots_8_uop_lrs3 : _GEN_2538; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_8_uop_lrs2 = slots_8_io_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2620 = issue_slots_8_grant ? issue_slots_8_uop_lrs2 : _GEN_2539; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_8_uop_lrs1 = slots_8_io_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2621 = issue_slots_8_grant ? issue_slots_8_uop_lrs1 : _GEN_2540; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_8_uop_ldst = slots_8_io_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2622 = issue_slots_8_grant ? issue_slots_8_uop_ldst : _GEN_2541; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_ldst_is_rs1 = slots_8_io_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2623 = issue_slots_8_grant ? issue_slots_8_uop_ldst_is_rs1 : _GEN_2542; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_flush_on_commit = slots_8_io_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2624 = issue_slots_8_grant ? issue_slots_8_uop_flush_on_commit : _GEN_2543; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_is_unique = slots_8_io_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2625 = issue_slots_8_grant ? issue_slots_8_uop_is_unique : _GEN_2544; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_is_sys_pc2epc = slots_8_io_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2626 = issue_slots_8_grant ? issue_slots_8_uop_is_sys_pc2epc : _GEN_2545; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_uses_stq = slots_8_io_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2627 = issue_slots_8_grant ? issue_slots_8_uop_uses_stq : _GEN_2546; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_uses_ldq = slots_8_io_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2628 = issue_slots_8_grant ? issue_slots_8_uop_uses_ldq : _GEN_2547; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_is_amo = slots_8_io_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2629 = issue_slots_8_grant ? issue_slots_8_uop_is_amo : _GEN_2548; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_is_fencei = slots_8_io_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2630 = issue_slots_8_grant ? issue_slots_8_uop_is_fencei : _GEN_2549; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_is_fence = slots_8_io_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2631 = issue_slots_8_grant ? issue_slots_8_uop_is_fence : _GEN_2550; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_mem_signed = slots_8_io_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2632 = issue_slots_8_grant ? issue_slots_8_uop_mem_signed : _GEN_2551; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_8_uop_mem_size = slots_8_io_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2633 = issue_slots_8_grant ? issue_slots_8_uop_mem_size : _GEN_2552; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_8_uop_mem_cmd = slots_8_io_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2634 = issue_slots_8_grant ? issue_slots_8_uop_mem_cmd : _GEN_2553; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_bypassable = slots_8_io_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2635 = issue_slots_8_grant ? issue_slots_8_uop_bypassable : _GEN_2554; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [63:0] issue_slots_8_uop_exc_cause = slots_8_io_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] _GEN_2636 = issue_slots_8_grant ? issue_slots_8_uop_exc_cause : _GEN_2555; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_exception = slots_8_io_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2637 = issue_slots_8_grant ? issue_slots_8_uop_exception : _GEN_2556; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_8_uop_stale_pdst = slots_8_io_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2638 = issue_slots_8_grant ? issue_slots_8_uop_stale_pdst : _GEN_2557; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_ppred_busy = slots_8_io_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2639 = issue_slots_8_grant ? issue_slots_8_uop_ppred_busy : _GEN_2558; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_prs3_busy = slots_8_io_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2640 = issue_slots_8_grant ? issue_slots_8_uop_prs3_busy : _GEN_2559; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_prs2_busy = slots_8_io_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2641 = issue_slots_8_grant ? issue_slots_8_uop_prs2_busy : _GEN_2560; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_prs1_busy = slots_8_io_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2642 = issue_slots_8_grant ? issue_slots_8_uop_prs1_busy : _GEN_2561; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_8_uop_ppred = slots_8_io_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2643 = issue_slots_8_grant ? issue_slots_8_uop_ppred : _GEN_2562; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_8_uop_prs3 = slots_8_io_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2644 = issue_slots_8_grant ? issue_slots_8_uop_prs3 : _GEN_2563; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_8_uop_prs2 = slots_8_io_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2645 = issue_slots_8_grant ? issue_slots_8_uop_prs2 : _GEN_2564; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_8_uop_prs1 = slots_8_io_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2646 = issue_slots_8_grant ? issue_slots_8_uop_prs1 : _GEN_2565; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_8_uop_pdst = slots_8_io_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2647 = issue_slots_8_grant ? issue_slots_8_uop_pdst : _GEN_2566; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_8_uop_rxq_idx = slots_8_io_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2648 = issue_slots_8_grant ? issue_slots_8_uop_rxq_idx : _GEN_2567; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_8_uop_stq_idx = slots_8_io_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2649 = issue_slots_8_grant ? issue_slots_8_uop_stq_idx : _GEN_2568; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_8_uop_ldq_idx = slots_8_io_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2650 = issue_slots_8_grant ? issue_slots_8_uop_ldq_idx : _GEN_2569; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_8_uop_rob_idx = slots_8_io_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2651 = issue_slots_8_grant ? issue_slots_8_uop_rob_idx : _GEN_2570; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [11:0] issue_slots_8_uop_csr_addr = slots_8_io_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2652 = issue_slots_8_grant ? issue_slots_8_uop_csr_addr : _GEN_2571; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [19:0] issue_slots_8_uop_imm_packed = slots_8_io_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] _GEN_2653 = issue_slots_8_grant ? issue_slots_8_uop_imm_packed : _GEN_2572; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_taken = slots_8_io_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2654 = issue_slots_8_grant ? issue_slots_8_uop_taken : _GEN_2573; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_8_uop_pc_lob = slots_8_io_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2655 = issue_slots_8_grant ? issue_slots_8_uop_pc_lob : _GEN_2574; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_edge_inst = slots_8_io_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2656 = issue_slots_8_grant ? issue_slots_8_uop_edge_inst : _GEN_2575; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_8_uop_ftq_idx = slots_8_io_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2657 = issue_slots_8_grant ? issue_slots_8_uop_ftq_idx : _GEN_2576; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_8_uop_br_tag = slots_8_io_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2658 = issue_slots_8_grant ? issue_slots_8_uop_br_tag : _GEN_2577; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [11:0] issue_slots_8_uop_br_mask = slots_8_io_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2659 = issue_slots_8_grant ? issue_slots_8_uop_br_mask : _GEN_2578; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_is_sfb = slots_8_io_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2660 = issue_slots_8_grant ? issue_slots_8_uop_is_sfb : _GEN_2579; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_is_jal = slots_8_io_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2661 = issue_slots_8_grant ? issue_slots_8_uop_is_jal : _GEN_2580; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_is_jalr = slots_8_io_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2662 = issue_slots_8_grant ? issue_slots_8_uop_is_jalr : _GEN_2581; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_is_br = slots_8_io_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2663 = issue_slots_8_grant ? issue_slots_8_uop_is_br : _GEN_2582; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_iw_p2_poisoned = slots_8_io_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2664 = issue_slots_8_grant ? issue_slots_8_uop_iw_p2_poisoned : _GEN_2583; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_iw_p1_poisoned = slots_8_io_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2665 = issue_slots_8_grant ? issue_slots_8_uop_iw_p1_poisoned : _GEN_2584; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_8_uop_iw_state = slots_8_io_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2666 = issue_slots_8_grant ? issue_slots_8_uop_iw_state : _GEN_2585; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_ctrl_is_std = slots_8_io_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2667 = issue_slots_8_grant ? issue_slots_8_uop_ctrl_is_std : _GEN_2586; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_ctrl_is_sta = slots_8_io_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2668 = issue_slots_8_grant ? issue_slots_8_uop_ctrl_is_sta : _GEN_2587; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_ctrl_is_load = slots_8_io_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2669 = issue_slots_8_grant ? issue_slots_8_uop_ctrl_is_load : _GEN_2588; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_8_uop_ctrl_csr_cmd = slots_8_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2670 = issue_slots_8_grant ? issue_slots_8_uop_ctrl_csr_cmd : _GEN_2589; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_ctrl_fcn_dw = slots_8_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2671 = issue_slots_8_grant ? issue_slots_8_uop_ctrl_fcn_dw : _GEN_2590; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_8_uop_ctrl_op_fcn = slots_8_io_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2672 = issue_slots_8_grant ? issue_slots_8_uop_ctrl_op_fcn : _GEN_2591; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_8_uop_ctrl_imm_sel = slots_8_io_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2673 = issue_slots_8_grant ? issue_slots_8_uop_ctrl_imm_sel : _GEN_2592; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_8_uop_ctrl_op2_sel = slots_8_io_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2674 = issue_slots_8_grant ? issue_slots_8_uop_ctrl_op2_sel : _GEN_2593; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_8_uop_ctrl_op1_sel = slots_8_io_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2675 = issue_slots_8_grant ? issue_slots_8_uop_ctrl_op1_sel : _GEN_2594; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_8_uop_ctrl_br_type = slots_8_io_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2676 = issue_slots_8_grant ? issue_slots_8_uop_ctrl_br_type : _GEN_2595; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [9:0] _GEN_2677 = issue_slots_8_grant ? issue_slots_8_uop_fu_code : _GEN_2596; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_8_uop_iq_type = slots_8_io_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2678 = issue_slots_8_grant ? issue_slots_8_uop_iq_type : _GEN_2597; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [39:0] issue_slots_8_uop_debug_pc = slots_8_io_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] _GEN_2679 = issue_slots_8_grant ? issue_slots_8_uop_debug_pc : _GEN_2598; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_8_uop_is_rvc = slots_8_io_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2680 = issue_slots_8_grant ? issue_slots_8_uop_is_rvc : _GEN_2599; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [31:0] issue_slots_8_uop_debug_inst = slots_8_io_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2681 = issue_slots_8_grant ? issue_slots_8_uop_debug_inst : _GEN_2600; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [31:0] issue_slots_8_uop_inst = slots_8_io_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2682 = issue_slots_8_grant ? issue_slots_8_uop_inst : _GEN_2601; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [6:0] issue_slots_8_uop_uopc = slots_8_io_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] _GEN_2683 = issue_slots_8_grant ? issue_slots_8_uop_uopc : _GEN_2602; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_9_uop_debug_tsrc = slots_9_io_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2686 = issue_slots_9_grant ? issue_slots_9_uop_debug_tsrc : _GEN_2605; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_9_uop_debug_fsrc = slots_9_io_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2687 = issue_slots_9_grant ? issue_slots_9_uop_debug_fsrc : _GEN_2606; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_bp_xcpt_if = slots_9_io_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2688 = issue_slots_9_grant ? issue_slots_9_uop_bp_xcpt_if : _GEN_2607; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_bp_debug_if = slots_9_io_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2689 = issue_slots_9_grant ? issue_slots_9_uop_bp_debug_if : _GEN_2608; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_xcpt_ma_if = slots_9_io_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2690 = issue_slots_9_grant ? issue_slots_9_uop_xcpt_ma_if : _GEN_2609; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_xcpt_ae_if = slots_9_io_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2691 = issue_slots_9_grant ? issue_slots_9_uop_xcpt_ae_if : _GEN_2610; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_xcpt_pf_if = slots_9_io_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2692 = issue_slots_9_grant ? issue_slots_9_uop_xcpt_pf_if : _GEN_2611; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_fp_single = slots_9_io_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2693 = issue_slots_9_grant ? issue_slots_9_uop_fp_single : _GEN_2612; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_fp_val = slots_9_io_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2694 = issue_slots_9_grant ? issue_slots_9_uop_fp_val : _GEN_2613; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_frs3_en = slots_9_io_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2695 = issue_slots_9_grant ? issue_slots_9_uop_frs3_en : _GEN_2614; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_9_uop_lrs2_rtype = slots_9_io_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2696 = issue_slots_9_grant ? issue_slots_9_uop_lrs2_rtype : _GEN_2615; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_9_uop_lrs1_rtype = slots_9_io_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2697 = issue_slots_9_grant ? issue_slots_9_uop_lrs1_rtype : _GEN_2616; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_9_uop_dst_rtype = slots_9_io_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2698 = issue_slots_9_grant ? issue_slots_9_uop_dst_rtype : _GEN_2617; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_ldst_val = slots_9_io_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2699 = issue_slots_9_grant ? issue_slots_9_uop_ldst_val : _GEN_2618; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_9_uop_lrs3 = slots_9_io_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2700 = issue_slots_9_grant ? issue_slots_9_uop_lrs3 : _GEN_2619; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_9_uop_lrs2 = slots_9_io_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2701 = issue_slots_9_grant ? issue_slots_9_uop_lrs2 : _GEN_2620; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_9_uop_lrs1 = slots_9_io_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2702 = issue_slots_9_grant ? issue_slots_9_uop_lrs1 : _GEN_2621; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_9_uop_ldst = slots_9_io_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2703 = issue_slots_9_grant ? issue_slots_9_uop_ldst : _GEN_2622; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_ldst_is_rs1 = slots_9_io_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2704 = issue_slots_9_grant ? issue_slots_9_uop_ldst_is_rs1 : _GEN_2623; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_flush_on_commit = slots_9_io_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2705 = issue_slots_9_grant ? issue_slots_9_uop_flush_on_commit : _GEN_2624; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_is_unique = slots_9_io_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2706 = issue_slots_9_grant ? issue_slots_9_uop_is_unique : _GEN_2625; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_is_sys_pc2epc = slots_9_io_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2707 = issue_slots_9_grant ? issue_slots_9_uop_is_sys_pc2epc : _GEN_2626; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_uses_stq = slots_9_io_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2708 = issue_slots_9_grant ? issue_slots_9_uop_uses_stq : _GEN_2627; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_uses_ldq = slots_9_io_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2709 = issue_slots_9_grant ? issue_slots_9_uop_uses_ldq : _GEN_2628; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_is_amo = slots_9_io_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2710 = issue_slots_9_grant ? issue_slots_9_uop_is_amo : _GEN_2629; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_is_fencei = slots_9_io_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2711 = issue_slots_9_grant ? issue_slots_9_uop_is_fencei : _GEN_2630; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_is_fence = slots_9_io_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2712 = issue_slots_9_grant ? issue_slots_9_uop_is_fence : _GEN_2631; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_mem_signed = slots_9_io_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2713 = issue_slots_9_grant ? issue_slots_9_uop_mem_signed : _GEN_2632; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_9_uop_mem_size = slots_9_io_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2714 = issue_slots_9_grant ? issue_slots_9_uop_mem_size : _GEN_2633; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_9_uop_mem_cmd = slots_9_io_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2715 = issue_slots_9_grant ? issue_slots_9_uop_mem_cmd : _GEN_2634; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_bypassable = slots_9_io_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2716 = issue_slots_9_grant ? issue_slots_9_uop_bypassable : _GEN_2635; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [63:0] issue_slots_9_uop_exc_cause = slots_9_io_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] _GEN_2717 = issue_slots_9_grant ? issue_slots_9_uop_exc_cause : _GEN_2636; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_exception = slots_9_io_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2718 = issue_slots_9_grant ? issue_slots_9_uop_exception : _GEN_2637; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_9_uop_stale_pdst = slots_9_io_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2719 = issue_slots_9_grant ? issue_slots_9_uop_stale_pdst : _GEN_2638; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_ppred_busy = slots_9_io_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2720 = issue_slots_9_grant ? issue_slots_9_uop_ppred_busy : _GEN_2639; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_prs3_busy = slots_9_io_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2721 = issue_slots_9_grant ? issue_slots_9_uop_prs3_busy : _GEN_2640; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_prs2_busy = slots_9_io_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2722 = issue_slots_9_grant ? issue_slots_9_uop_prs2_busy : _GEN_2641; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_prs1_busy = slots_9_io_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2723 = issue_slots_9_grant ? issue_slots_9_uop_prs1_busy : _GEN_2642; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_9_uop_ppred = slots_9_io_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2724 = issue_slots_9_grant ? issue_slots_9_uop_ppred : _GEN_2643; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_9_uop_prs3 = slots_9_io_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2725 = issue_slots_9_grant ? issue_slots_9_uop_prs3 : _GEN_2644; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_9_uop_prs2 = slots_9_io_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2726 = issue_slots_9_grant ? issue_slots_9_uop_prs2 : _GEN_2645; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_9_uop_prs1 = slots_9_io_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2727 = issue_slots_9_grant ? issue_slots_9_uop_prs1 : _GEN_2646; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_9_uop_pdst = slots_9_io_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2728 = issue_slots_9_grant ? issue_slots_9_uop_pdst : _GEN_2647; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_9_uop_rxq_idx = slots_9_io_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2729 = issue_slots_9_grant ? issue_slots_9_uop_rxq_idx : _GEN_2648; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_9_uop_stq_idx = slots_9_io_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2730 = issue_slots_9_grant ? issue_slots_9_uop_stq_idx : _GEN_2649; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_9_uop_ldq_idx = slots_9_io_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2731 = issue_slots_9_grant ? issue_slots_9_uop_ldq_idx : _GEN_2650; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_9_uop_rob_idx = slots_9_io_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2732 = issue_slots_9_grant ? issue_slots_9_uop_rob_idx : _GEN_2651; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [11:0] issue_slots_9_uop_csr_addr = slots_9_io_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2733 = issue_slots_9_grant ? issue_slots_9_uop_csr_addr : _GEN_2652; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [19:0] issue_slots_9_uop_imm_packed = slots_9_io_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] _GEN_2734 = issue_slots_9_grant ? issue_slots_9_uop_imm_packed : _GEN_2653; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_taken = slots_9_io_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2735 = issue_slots_9_grant ? issue_slots_9_uop_taken : _GEN_2654; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_9_uop_pc_lob = slots_9_io_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2736 = issue_slots_9_grant ? issue_slots_9_uop_pc_lob : _GEN_2655; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_edge_inst = slots_9_io_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2737 = issue_slots_9_grant ? issue_slots_9_uop_edge_inst : _GEN_2656; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_9_uop_ftq_idx = slots_9_io_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2738 = issue_slots_9_grant ? issue_slots_9_uop_ftq_idx : _GEN_2657; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_9_uop_br_tag = slots_9_io_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2739 = issue_slots_9_grant ? issue_slots_9_uop_br_tag : _GEN_2658; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [11:0] issue_slots_9_uop_br_mask = slots_9_io_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2740 = issue_slots_9_grant ? issue_slots_9_uop_br_mask : _GEN_2659; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_is_sfb = slots_9_io_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2741 = issue_slots_9_grant ? issue_slots_9_uop_is_sfb : _GEN_2660; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_is_jal = slots_9_io_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2742 = issue_slots_9_grant ? issue_slots_9_uop_is_jal : _GEN_2661; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_is_jalr = slots_9_io_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2743 = issue_slots_9_grant ? issue_slots_9_uop_is_jalr : _GEN_2662; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_is_br = slots_9_io_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2744 = issue_slots_9_grant ? issue_slots_9_uop_is_br : _GEN_2663; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_iw_p2_poisoned = slots_9_io_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2745 = issue_slots_9_grant ? issue_slots_9_uop_iw_p2_poisoned : _GEN_2664; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_iw_p1_poisoned = slots_9_io_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2746 = issue_slots_9_grant ? issue_slots_9_uop_iw_p1_poisoned : _GEN_2665; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_9_uop_iw_state = slots_9_io_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2747 = issue_slots_9_grant ? issue_slots_9_uop_iw_state : _GEN_2666; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_ctrl_is_std = slots_9_io_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2748 = issue_slots_9_grant ? issue_slots_9_uop_ctrl_is_std : _GEN_2667; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_ctrl_is_sta = slots_9_io_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2749 = issue_slots_9_grant ? issue_slots_9_uop_ctrl_is_sta : _GEN_2668; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_ctrl_is_load = slots_9_io_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2750 = issue_slots_9_grant ? issue_slots_9_uop_ctrl_is_load : _GEN_2669; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_9_uop_ctrl_csr_cmd = slots_9_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2751 = issue_slots_9_grant ? issue_slots_9_uop_ctrl_csr_cmd : _GEN_2670; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_ctrl_fcn_dw = slots_9_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2752 = issue_slots_9_grant ? issue_slots_9_uop_ctrl_fcn_dw : _GEN_2671; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_9_uop_ctrl_op_fcn = slots_9_io_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2753 = issue_slots_9_grant ? issue_slots_9_uop_ctrl_op_fcn : _GEN_2672; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_9_uop_ctrl_imm_sel = slots_9_io_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2754 = issue_slots_9_grant ? issue_slots_9_uop_ctrl_imm_sel : _GEN_2673; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_9_uop_ctrl_op2_sel = slots_9_io_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2755 = issue_slots_9_grant ? issue_slots_9_uop_ctrl_op2_sel : _GEN_2674; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_9_uop_ctrl_op1_sel = slots_9_io_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2756 = issue_slots_9_grant ? issue_slots_9_uop_ctrl_op1_sel : _GEN_2675; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_9_uop_ctrl_br_type = slots_9_io_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2757 = issue_slots_9_grant ? issue_slots_9_uop_ctrl_br_type : _GEN_2676; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [9:0] _GEN_2758 = issue_slots_9_grant ? issue_slots_9_uop_fu_code : _GEN_2677; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_9_uop_iq_type = slots_9_io_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2759 = issue_slots_9_grant ? issue_slots_9_uop_iq_type : _GEN_2678; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [39:0] issue_slots_9_uop_debug_pc = slots_9_io_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] _GEN_2760 = issue_slots_9_grant ? issue_slots_9_uop_debug_pc : _GEN_2679; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_9_uop_is_rvc = slots_9_io_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2761 = issue_slots_9_grant ? issue_slots_9_uop_is_rvc : _GEN_2680; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [31:0] issue_slots_9_uop_debug_inst = slots_9_io_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2762 = issue_slots_9_grant ? issue_slots_9_uop_debug_inst : _GEN_2681; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [31:0] issue_slots_9_uop_inst = slots_9_io_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2763 = issue_slots_9_grant ? issue_slots_9_uop_inst : _GEN_2682; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [6:0] issue_slots_9_uop_uopc = slots_9_io_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] _GEN_2764 = issue_slots_9_grant ? issue_slots_9_uop_uopc : _GEN_2683; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_10_uop_debug_tsrc = slots_10_io_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2767 = issue_slots_10_grant ? issue_slots_10_uop_debug_tsrc : _GEN_2686; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_10_uop_debug_fsrc = slots_10_io_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2768 = issue_slots_10_grant ? issue_slots_10_uop_debug_fsrc : _GEN_2687; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_bp_xcpt_if = slots_10_io_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2769 = issue_slots_10_grant ? issue_slots_10_uop_bp_xcpt_if : _GEN_2688; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_bp_debug_if = slots_10_io_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2770 = issue_slots_10_grant ? issue_slots_10_uop_bp_debug_if : _GEN_2689; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_xcpt_ma_if = slots_10_io_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2771 = issue_slots_10_grant ? issue_slots_10_uop_xcpt_ma_if : _GEN_2690; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_xcpt_ae_if = slots_10_io_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2772 = issue_slots_10_grant ? issue_slots_10_uop_xcpt_ae_if : _GEN_2691; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_xcpt_pf_if = slots_10_io_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2773 = issue_slots_10_grant ? issue_slots_10_uop_xcpt_pf_if : _GEN_2692; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_fp_single = slots_10_io_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2774 = issue_slots_10_grant ? issue_slots_10_uop_fp_single : _GEN_2693; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_fp_val = slots_10_io_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2775 = issue_slots_10_grant ? issue_slots_10_uop_fp_val : _GEN_2694; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_frs3_en = slots_10_io_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2776 = issue_slots_10_grant ? issue_slots_10_uop_frs3_en : _GEN_2695; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_10_uop_lrs2_rtype = slots_10_io_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2777 = issue_slots_10_grant ? issue_slots_10_uop_lrs2_rtype : _GEN_2696; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_10_uop_lrs1_rtype = slots_10_io_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2778 = issue_slots_10_grant ? issue_slots_10_uop_lrs1_rtype : _GEN_2697; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_10_uop_dst_rtype = slots_10_io_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2779 = issue_slots_10_grant ? issue_slots_10_uop_dst_rtype : _GEN_2698; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_ldst_val = slots_10_io_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2780 = issue_slots_10_grant ? issue_slots_10_uop_ldst_val : _GEN_2699; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_10_uop_lrs3 = slots_10_io_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2781 = issue_slots_10_grant ? issue_slots_10_uop_lrs3 : _GEN_2700; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_10_uop_lrs2 = slots_10_io_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2782 = issue_slots_10_grant ? issue_slots_10_uop_lrs2 : _GEN_2701; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_10_uop_lrs1 = slots_10_io_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2783 = issue_slots_10_grant ? issue_slots_10_uop_lrs1 : _GEN_2702; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_10_uop_ldst = slots_10_io_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2784 = issue_slots_10_grant ? issue_slots_10_uop_ldst : _GEN_2703; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_ldst_is_rs1 = slots_10_io_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2785 = issue_slots_10_grant ? issue_slots_10_uop_ldst_is_rs1 : _GEN_2704; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_flush_on_commit = slots_10_io_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2786 = issue_slots_10_grant ? issue_slots_10_uop_flush_on_commit : _GEN_2705; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_is_unique = slots_10_io_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2787 = issue_slots_10_grant ? issue_slots_10_uop_is_unique : _GEN_2706; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_is_sys_pc2epc = slots_10_io_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2788 = issue_slots_10_grant ? issue_slots_10_uop_is_sys_pc2epc : _GEN_2707; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_uses_stq = slots_10_io_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2789 = issue_slots_10_grant ? issue_slots_10_uop_uses_stq : _GEN_2708; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_uses_ldq = slots_10_io_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2790 = issue_slots_10_grant ? issue_slots_10_uop_uses_ldq : _GEN_2709; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_is_amo = slots_10_io_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2791 = issue_slots_10_grant ? issue_slots_10_uop_is_amo : _GEN_2710; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_is_fencei = slots_10_io_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2792 = issue_slots_10_grant ? issue_slots_10_uop_is_fencei : _GEN_2711; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_is_fence = slots_10_io_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2793 = issue_slots_10_grant ? issue_slots_10_uop_is_fence : _GEN_2712; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_mem_signed = slots_10_io_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2794 = issue_slots_10_grant ? issue_slots_10_uop_mem_signed : _GEN_2713; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_10_uop_mem_size = slots_10_io_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2795 = issue_slots_10_grant ? issue_slots_10_uop_mem_size : _GEN_2714; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_10_uop_mem_cmd = slots_10_io_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2796 = issue_slots_10_grant ? issue_slots_10_uop_mem_cmd : _GEN_2715; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_bypassable = slots_10_io_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2797 = issue_slots_10_grant ? issue_slots_10_uop_bypassable : _GEN_2716; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [63:0] issue_slots_10_uop_exc_cause = slots_10_io_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] _GEN_2798 = issue_slots_10_grant ? issue_slots_10_uop_exc_cause : _GEN_2717; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_exception = slots_10_io_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2799 = issue_slots_10_grant ? issue_slots_10_uop_exception : _GEN_2718; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_10_uop_stale_pdst = slots_10_io_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2800 = issue_slots_10_grant ? issue_slots_10_uop_stale_pdst : _GEN_2719; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_ppred_busy = slots_10_io_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2801 = issue_slots_10_grant ? issue_slots_10_uop_ppred_busy : _GEN_2720; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_prs3_busy = slots_10_io_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2802 = issue_slots_10_grant ? issue_slots_10_uop_prs3_busy : _GEN_2721; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_prs2_busy = slots_10_io_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2803 = issue_slots_10_grant ? issue_slots_10_uop_prs2_busy : _GEN_2722; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_prs1_busy = slots_10_io_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2804 = issue_slots_10_grant ? issue_slots_10_uop_prs1_busy : _GEN_2723; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_10_uop_ppred = slots_10_io_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2805 = issue_slots_10_grant ? issue_slots_10_uop_ppred : _GEN_2724; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_10_uop_prs3 = slots_10_io_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2806 = issue_slots_10_grant ? issue_slots_10_uop_prs3 : _GEN_2725; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_10_uop_prs2 = slots_10_io_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2807 = issue_slots_10_grant ? issue_slots_10_uop_prs2 : _GEN_2726; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_10_uop_prs1 = slots_10_io_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2808 = issue_slots_10_grant ? issue_slots_10_uop_prs1 : _GEN_2727; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_10_uop_pdst = slots_10_io_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2809 = issue_slots_10_grant ? issue_slots_10_uop_pdst : _GEN_2728; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_10_uop_rxq_idx = slots_10_io_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2810 = issue_slots_10_grant ? issue_slots_10_uop_rxq_idx : _GEN_2729; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_10_uop_stq_idx = slots_10_io_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2811 = issue_slots_10_grant ? issue_slots_10_uop_stq_idx : _GEN_2730; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_10_uop_ldq_idx = slots_10_io_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2812 = issue_slots_10_grant ? issue_slots_10_uop_ldq_idx : _GEN_2731; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_10_uop_rob_idx = slots_10_io_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2813 = issue_slots_10_grant ? issue_slots_10_uop_rob_idx : _GEN_2732; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [11:0] issue_slots_10_uop_csr_addr = slots_10_io_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2814 = issue_slots_10_grant ? issue_slots_10_uop_csr_addr : _GEN_2733; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [19:0] issue_slots_10_uop_imm_packed = slots_10_io_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] _GEN_2815 = issue_slots_10_grant ? issue_slots_10_uop_imm_packed : _GEN_2734; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_taken = slots_10_io_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2816 = issue_slots_10_grant ? issue_slots_10_uop_taken : _GEN_2735; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [5:0] issue_slots_10_uop_pc_lob = slots_10_io_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] _GEN_2817 = issue_slots_10_grant ? issue_slots_10_uop_pc_lob : _GEN_2736; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_edge_inst = slots_10_io_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2818 = issue_slots_10_grant ? issue_slots_10_uop_edge_inst : _GEN_2737; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [4:0] issue_slots_10_uop_ftq_idx = slots_10_io_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] _GEN_2819 = issue_slots_10_grant ? issue_slots_10_uop_ftq_idx : _GEN_2738; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_10_uop_br_tag = slots_10_io_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2820 = issue_slots_10_grant ? issue_slots_10_uop_br_tag : _GEN_2739; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [11:0] issue_slots_10_uop_br_mask = slots_10_io_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] _GEN_2821 = issue_slots_10_grant ? issue_slots_10_uop_br_mask : _GEN_2740; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_is_sfb = slots_10_io_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2822 = issue_slots_10_grant ? issue_slots_10_uop_is_sfb : _GEN_2741; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_is_jal = slots_10_io_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2823 = issue_slots_10_grant ? issue_slots_10_uop_is_jal : _GEN_2742; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_is_jalr = slots_10_io_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2824 = issue_slots_10_grant ? issue_slots_10_uop_is_jalr : _GEN_2743; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_is_br = slots_10_io_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2825 = issue_slots_10_grant ? issue_slots_10_uop_is_br : _GEN_2744; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_iw_p2_poisoned = slots_10_io_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2826 = issue_slots_10_grant ? issue_slots_10_uop_iw_p2_poisoned : _GEN_2745; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_iw_p1_poisoned = slots_10_io_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2827 = issue_slots_10_grant ? issue_slots_10_uop_iw_p1_poisoned : _GEN_2746; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_10_uop_iw_state = slots_10_io_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2828 = issue_slots_10_grant ? issue_slots_10_uop_iw_state : _GEN_2747; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_ctrl_is_std = slots_10_io_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2829 = issue_slots_10_grant ? issue_slots_10_uop_ctrl_is_std : _GEN_2748; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_ctrl_is_sta = slots_10_io_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2830 = issue_slots_10_grant ? issue_slots_10_uop_ctrl_is_sta : _GEN_2749; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_ctrl_is_load = slots_10_io_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2831 = issue_slots_10_grant ? issue_slots_10_uop_ctrl_is_load : _GEN_2750; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_10_uop_ctrl_csr_cmd = slots_10_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2832 = issue_slots_10_grant ? issue_slots_10_uop_ctrl_csr_cmd : _GEN_2751; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_ctrl_fcn_dw = slots_10_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2833 = issue_slots_10_grant ? issue_slots_10_uop_ctrl_fcn_dw : _GEN_2752; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_10_uop_ctrl_op_fcn = slots_10_io_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2834 = issue_slots_10_grant ? issue_slots_10_uop_ctrl_op_fcn : _GEN_2753; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_10_uop_ctrl_imm_sel = slots_10_io_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2835 = issue_slots_10_grant ? issue_slots_10_uop_ctrl_imm_sel : _GEN_2754; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_10_uop_ctrl_op2_sel = slots_10_io_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2836 = issue_slots_10_grant ? issue_slots_10_uop_ctrl_op2_sel : _GEN_2755; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_10_uop_ctrl_op1_sel = slots_10_io_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] _GEN_2837 = issue_slots_10_grant ? issue_slots_10_uop_ctrl_op1_sel : _GEN_2756; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [3:0] issue_slots_10_uop_ctrl_br_type = slots_10_io_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] _GEN_2838 = issue_slots_10_grant ? issue_slots_10_uop_ctrl_br_type : _GEN_2757; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [9:0] _GEN_2839 = issue_slots_10_grant ? issue_slots_10_uop_fu_code : _GEN_2758; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [2:0] issue_slots_10_uop_iq_type = slots_10_io_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] _GEN_2840 = issue_slots_10_grant ? issue_slots_10_uop_iq_type : _GEN_2759; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [39:0] issue_slots_10_uop_debug_pc = slots_10_io_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] _GEN_2841 = issue_slots_10_grant ? issue_slots_10_uop_debug_pc : _GEN_2760; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire  issue_slots_10_uop_is_rvc = slots_10_io_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  _GEN_2842 = issue_slots_10_grant ? issue_slots_10_uop_is_rvc : _GEN_2761; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [31:0] issue_slots_10_uop_debug_inst = slots_10_io_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2843 = issue_slots_10_grant ? issue_slots_10_uop_debug_inst : _GEN_2762; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [31:0] issue_slots_10_uop_inst = slots_10_io_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] _GEN_2844 = issue_slots_10_grant ? issue_slots_10_uop_inst : _GEN_2763; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [6:0] issue_slots_10_uop_uopc = slots_10_io_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] _GEN_2845 = issue_slots_10_grant ? issue_slots_10_uop_uopc : _GEN_2764; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  wire [1:0] issue_slots_11_uop_debug_tsrc = slots_11_io_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_11_uop_debug_fsrc = slots_11_io_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_bp_xcpt_if = slots_11_io_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_bp_debug_if = slots_11_io_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_xcpt_ma_if = slots_11_io_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_xcpt_ae_if = slots_11_io_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_xcpt_pf_if = slots_11_io_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_fp_single = slots_11_io_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_fp_val = slots_11_io_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_frs3_en = slots_11_io_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_11_uop_lrs2_rtype = slots_11_io_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_11_uop_lrs1_rtype = slots_11_io_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_11_uop_dst_rtype = slots_11_io_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_ldst_val = slots_11_io_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_uop_lrs3 = slots_11_io_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_uop_lrs2 = slots_11_io_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_uop_lrs1 = slots_11_io_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_uop_ldst = slots_11_io_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_ldst_is_rs1 = slots_11_io_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_flush_on_commit = slots_11_io_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_is_unique = slots_11_io_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_is_sys_pc2epc = slots_11_io_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_uses_stq = slots_11_io_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_uses_ldq = slots_11_io_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_is_amo = slots_11_io_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_is_fencei = slots_11_io_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_is_fence = slots_11_io_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_mem_signed = slots_11_io_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_11_uop_mem_size = slots_11_io_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_11_uop_mem_cmd = slots_11_io_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_bypassable = slots_11_io_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [63:0] issue_slots_11_uop_exc_cause = slots_11_io_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_exception = slots_11_io_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_uop_stale_pdst = slots_11_io_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_ppred_busy = slots_11_io_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_prs3_busy = slots_11_io_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_prs2_busy = slots_11_io_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_prs1_busy = slots_11_io_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_11_uop_ppred = slots_11_io_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_uop_prs3 = slots_11_io_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_uop_prs2 = slots_11_io_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_uop_prs1 = slots_11_io_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_uop_pdst = slots_11_io_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_11_uop_rxq_idx = slots_11_io_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_11_uop_stq_idx = slots_11_io_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_11_uop_ldq_idx = slots_11_io_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_uop_rob_idx = slots_11_io_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_11_uop_csr_addr = slots_11_io_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [19:0] issue_slots_11_uop_imm_packed = slots_11_io_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_taken = slots_11_io_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [5:0] issue_slots_11_uop_pc_lob = slots_11_io_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_edge_inst = slots_11_io_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [4:0] issue_slots_11_uop_ftq_idx = slots_11_io_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_11_uop_br_tag = slots_11_io_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [11:0] issue_slots_11_uop_br_mask = slots_11_io_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_is_sfb = slots_11_io_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_is_jal = slots_11_io_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_is_jalr = slots_11_io_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_is_br = slots_11_io_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_iw_p2_poisoned = slots_11_io_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_iw_p1_poisoned = slots_11_io_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_11_uop_iw_state = slots_11_io_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_ctrl_is_std = slots_11_io_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_ctrl_is_sta = slots_11_io_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_ctrl_is_load = slots_11_io_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_11_uop_ctrl_csr_cmd = slots_11_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_ctrl_fcn_dw = slots_11_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_11_uop_ctrl_op_fcn = slots_11_io_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_11_uop_ctrl_imm_sel = slots_11_io_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_11_uop_ctrl_op2_sel = slots_11_io_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [1:0] issue_slots_11_uop_ctrl_op1_sel = slots_11_io_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [3:0] issue_slots_11_uop_ctrl_br_type = slots_11_io_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [2:0] issue_slots_11_uop_iq_type = slots_11_io_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [39:0] issue_slots_11_uop_debug_pc = slots_11_io_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire  issue_slots_11_uop_is_rvc = slots_11_io_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_11_uop_debug_inst = slots_11_io_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [31:0] issue_slots_11_uop_inst = slots_11_io_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  wire [6:0] issue_slots_11_uop_uopc = slots_11_io_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 154:28]
  IssueSlot_16 slots_0 ( // @[issue-unit.scala 153:73]
    .clock(slots_0_clock),
    .reset(slots_0_reset),
    .io_valid(slots_0_io_valid),
    .io_will_be_valid(slots_0_io_will_be_valid),
    .io_request(slots_0_io_request),
    .io_request_hp(slots_0_io_request_hp),
    .io_grant(slots_0_io_grant),
    .io_brupdate_b1_resolve_mask(slots_0_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_0_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_uopc(slots_0_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_0_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_0_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_0_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_0_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_0_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_0_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_0_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_0_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_0_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_0_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_0_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_0_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_0_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_0_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_0_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_0_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_iw_state(slots_0_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_0_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_0_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_0_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_0_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_0_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_0_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_0_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_0_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_0_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_0_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_0_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_0_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_0_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_0_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_0_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_0_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_0_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_0_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_0_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_0_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_0_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_0_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_0_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_0_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_0_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_0_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_0_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_0_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_0_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_0_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_0_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_0_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_0_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_0_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_0_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_0_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_0_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_0_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_0_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_0_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_0_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_0_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_0_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_0_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_0_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_0_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_0_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_0_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_0_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_0_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_0_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_0_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_0_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_0_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_0_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_0_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_0_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_0_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_0_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_0_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_0_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_0_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_0_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_0_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_0_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_0_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_0_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_0_io_brupdate_b2_target_offset),
    .io_kill(slots_0_io_kill),
    .io_clear(slots_0_io_clear),
    .io_ldspec_miss(slots_0_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_0_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_0_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_0_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_1_valid(slots_0_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_0_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_0_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_2_valid(slots_0_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_0_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_0_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_3_valid(slots_0_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_0_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_0_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_4_valid(slots_0_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_0_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_0_io_wakeup_ports_4_bits_poisoned),
    .io_pred_wakeup_port_valid(slots_0_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_0_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_0_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_0_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_0_io_in_uop_valid),
    .io_in_uop_bits_uopc(slots_0_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_0_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_0_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_0_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_0_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_0_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_0_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_0_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_0_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_0_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_0_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_0_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_0_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_0_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_0_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_0_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_0_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_iw_state(slots_0_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_0_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_0_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_0_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_0_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_0_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_0_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_0_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_0_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_0_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_0_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_0_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_0_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_0_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_0_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_0_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_0_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_0_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_0_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_0_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_0_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_0_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_0_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_0_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_0_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_0_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_0_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_0_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_0_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_0_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_0_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_0_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_0_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_0_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_0_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_0_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_0_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_0_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_0_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_0_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_0_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_0_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_0_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_0_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_0_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_0_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_0_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_0_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_0_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_0_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_0_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_0_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_0_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_0_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_0_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_0_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_0_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_0_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_0_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_0_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_0_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_0_io_in_uop_bits_debug_tsrc),
    .io_out_uop_uopc(slots_0_io_out_uop_uopc),
    .io_out_uop_inst(slots_0_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_0_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_0_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_0_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_0_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_0_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_0_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_0_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_0_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_0_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_0_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_0_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_0_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_0_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_0_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_0_io_out_uop_ctrl_is_std),
    .io_out_uop_iw_state(slots_0_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_0_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_0_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_0_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_0_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_0_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_0_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_0_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_0_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_0_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_0_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_0_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_0_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_0_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_0_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_0_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_0_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_0_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_0_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_0_io_out_uop_pdst),
    .io_out_uop_prs1(slots_0_io_out_uop_prs1),
    .io_out_uop_prs2(slots_0_io_out_uop_prs2),
    .io_out_uop_prs3(slots_0_io_out_uop_prs3),
    .io_out_uop_ppred(slots_0_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_0_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_0_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_0_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_0_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_0_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_0_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_0_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_0_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_0_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_0_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_0_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_0_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_0_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_0_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_0_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_0_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_0_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_0_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_0_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_0_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_0_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_0_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_0_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_0_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_0_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_0_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_0_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_0_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_0_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_0_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_0_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_0_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_0_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_0_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_0_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_0_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_0_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_0_io_out_uop_debug_tsrc),
    .io_uop_uopc(slots_0_io_uop_uopc),
    .io_uop_inst(slots_0_io_uop_inst),
    .io_uop_debug_inst(slots_0_io_uop_debug_inst),
    .io_uop_is_rvc(slots_0_io_uop_is_rvc),
    .io_uop_debug_pc(slots_0_io_uop_debug_pc),
    .io_uop_iq_type(slots_0_io_uop_iq_type),
    .io_uop_fu_code(slots_0_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_0_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_0_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_0_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_0_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_0_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_0_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_0_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_0_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_0_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_0_io_uop_ctrl_is_std),
    .io_uop_iw_state(slots_0_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_0_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_0_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_0_io_uop_is_br),
    .io_uop_is_jalr(slots_0_io_uop_is_jalr),
    .io_uop_is_jal(slots_0_io_uop_is_jal),
    .io_uop_is_sfb(slots_0_io_uop_is_sfb),
    .io_uop_br_mask(slots_0_io_uop_br_mask),
    .io_uop_br_tag(slots_0_io_uop_br_tag),
    .io_uop_ftq_idx(slots_0_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_0_io_uop_edge_inst),
    .io_uop_pc_lob(slots_0_io_uop_pc_lob),
    .io_uop_taken(slots_0_io_uop_taken),
    .io_uop_imm_packed(slots_0_io_uop_imm_packed),
    .io_uop_csr_addr(slots_0_io_uop_csr_addr),
    .io_uop_rob_idx(slots_0_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_0_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_0_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_0_io_uop_rxq_idx),
    .io_uop_pdst(slots_0_io_uop_pdst),
    .io_uop_prs1(slots_0_io_uop_prs1),
    .io_uop_prs2(slots_0_io_uop_prs2),
    .io_uop_prs3(slots_0_io_uop_prs3),
    .io_uop_ppred(slots_0_io_uop_ppred),
    .io_uop_prs1_busy(slots_0_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_0_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_0_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_0_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_0_io_uop_stale_pdst),
    .io_uop_exception(slots_0_io_uop_exception),
    .io_uop_exc_cause(slots_0_io_uop_exc_cause),
    .io_uop_bypassable(slots_0_io_uop_bypassable),
    .io_uop_mem_cmd(slots_0_io_uop_mem_cmd),
    .io_uop_mem_size(slots_0_io_uop_mem_size),
    .io_uop_mem_signed(slots_0_io_uop_mem_signed),
    .io_uop_is_fence(slots_0_io_uop_is_fence),
    .io_uop_is_fencei(slots_0_io_uop_is_fencei),
    .io_uop_is_amo(slots_0_io_uop_is_amo),
    .io_uop_uses_ldq(slots_0_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_0_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_0_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_0_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_0_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_0_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_0_io_uop_ldst),
    .io_uop_lrs1(slots_0_io_uop_lrs1),
    .io_uop_lrs2(slots_0_io_uop_lrs2),
    .io_uop_lrs3(slots_0_io_uop_lrs3),
    .io_uop_ldst_val(slots_0_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_0_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_0_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_0_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_0_io_uop_frs3_en),
    .io_uop_fp_val(slots_0_io_uop_fp_val),
    .io_uop_fp_single(slots_0_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_0_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_0_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_0_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_0_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_0_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_0_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_0_io_uop_debug_tsrc),
    .io_debug_p1(slots_0_io_debug_p1),
    .io_debug_p2(slots_0_io_debug_p2),
    .io_debug_p3(slots_0_io_debug_p3),
    .io_debug_ppred(slots_0_io_debug_ppred),
    .io_debug_state(slots_0_io_debug_state)
  );
  IssueSlot_16 slots_1 ( // @[issue-unit.scala 153:73]
    .clock(slots_1_clock),
    .reset(slots_1_reset),
    .io_valid(slots_1_io_valid),
    .io_will_be_valid(slots_1_io_will_be_valid),
    .io_request(slots_1_io_request),
    .io_request_hp(slots_1_io_request_hp),
    .io_grant(slots_1_io_grant),
    .io_brupdate_b1_resolve_mask(slots_1_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_1_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_uopc(slots_1_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_1_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_1_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_1_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_1_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_1_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_1_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_1_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_1_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_1_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_1_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_1_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_1_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_1_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_1_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_1_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_1_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_iw_state(slots_1_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_1_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_1_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_1_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_1_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_1_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_1_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_1_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_1_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_1_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_1_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_1_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_1_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_1_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_1_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_1_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_1_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_1_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_1_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_1_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_1_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_1_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_1_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_1_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_1_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_1_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_1_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_1_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_1_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_1_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_1_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_1_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_1_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_1_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_1_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_1_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_1_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_1_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_1_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_1_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_1_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_1_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_1_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_1_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_1_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_1_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_1_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_1_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_1_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_1_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_1_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_1_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_1_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_1_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_1_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_1_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_1_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_1_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_1_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_1_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_1_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_1_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_1_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_1_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_1_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_1_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_1_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_1_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_1_io_brupdate_b2_target_offset),
    .io_kill(slots_1_io_kill),
    .io_clear(slots_1_io_clear),
    .io_ldspec_miss(slots_1_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_1_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_1_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_1_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_1_valid(slots_1_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_1_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_1_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_2_valid(slots_1_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_1_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_1_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_3_valid(slots_1_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_1_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_1_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_4_valid(slots_1_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_1_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_1_io_wakeup_ports_4_bits_poisoned),
    .io_pred_wakeup_port_valid(slots_1_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_1_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_1_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_1_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_1_io_in_uop_valid),
    .io_in_uop_bits_uopc(slots_1_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_1_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_1_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_1_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_1_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_1_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_1_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_1_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_1_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_1_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_1_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_1_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_1_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_1_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_1_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_1_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_1_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_iw_state(slots_1_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_1_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_1_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_1_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_1_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_1_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_1_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_1_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_1_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_1_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_1_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_1_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_1_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_1_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_1_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_1_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_1_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_1_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_1_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_1_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_1_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_1_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_1_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_1_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_1_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_1_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_1_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_1_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_1_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_1_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_1_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_1_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_1_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_1_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_1_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_1_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_1_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_1_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_1_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_1_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_1_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_1_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_1_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_1_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_1_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_1_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_1_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_1_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_1_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_1_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_1_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_1_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_1_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_1_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_1_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_1_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_1_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_1_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_1_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_1_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_1_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_1_io_in_uop_bits_debug_tsrc),
    .io_out_uop_uopc(slots_1_io_out_uop_uopc),
    .io_out_uop_inst(slots_1_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_1_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_1_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_1_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_1_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_1_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_1_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_1_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_1_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_1_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_1_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_1_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_1_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_1_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_1_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_1_io_out_uop_ctrl_is_std),
    .io_out_uop_iw_state(slots_1_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_1_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_1_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_1_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_1_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_1_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_1_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_1_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_1_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_1_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_1_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_1_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_1_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_1_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_1_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_1_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_1_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_1_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_1_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_1_io_out_uop_pdst),
    .io_out_uop_prs1(slots_1_io_out_uop_prs1),
    .io_out_uop_prs2(slots_1_io_out_uop_prs2),
    .io_out_uop_prs3(slots_1_io_out_uop_prs3),
    .io_out_uop_ppred(slots_1_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_1_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_1_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_1_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_1_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_1_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_1_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_1_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_1_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_1_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_1_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_1_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_1_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_1_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_1_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_1_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_1_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_1_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_1_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_1_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_1_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_1_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_1_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_1_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_1_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_1_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_1_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_1_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_1_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_1_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_1_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_1_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_1_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_1_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_1_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_1_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_1_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_1_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_1_io_out_uop_debug_tsrc),
    .io_uop_uopc(slots_1_io_uop_uopc),
    .io_uop_inst(slots_1_io_uop_inst),
    .io_uop_debug_inst(slots_1_io_uop_debug_inst),
    .io_uop_is_rvc(slots_1_io_uop_is_rvc),
    .io_uop_debug_pc(slots_1_io_uop_debug_pc),
    .io_uop_iq_type(slots_1_io_uop_iq_type),
    .io_uop_fu_code(slots_1_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_1_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_1_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_1_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_1_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_1_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_1_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_1_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_1_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_1_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_1_io_uop_ctrl_is_std),
    .io_uop_iw_state(slots_1_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_1_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_1_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_1_io_uop_is_br),
    .io_uop_is_jalr(slots_1_io_uop_is_jalr),
    .io_uop_is_jal(slots_1_io_uop_is_jal),
    .io_uop_is_sfb(slots_1_io_uop_is_sfb),
    .io_uop_br_mask(slots_1_io_uop_br_mask),
    .io_uop_br_tag(slots_1_io_uop_br_tag),
    .io_uop_ftq_idx(slots_1_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_1_io_uop_edge_inst),
    .io_uop_pc_lob(slots_1_io_uop_pc_lob),
    .io_uop_taken(slots_1_io_uop_taken),
    .io_uop_imm_packed(slots_1_io_uop_imm_packed),
    .io_uop_csr_addr(slots_1_io_uop_csr_addr),
    .io_uop_rob_idx(slots_1_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_1_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_1_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_1_io_uop_rxq_idx),
    .io_uop_pdst(slots_1_io_uop_pdst),
    .io_uop_prs1(slots_1_io_uop_prs1),
    .io_uop_prs2(slots_1_io_uop_prs2),
    .io_uop_prs3(slots_1_io_uop_prs3),
    .io_uop_ppred(slots_1_io_uop_ppred),
    .io_uop_prs1_busy(slots_1_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_1_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_1_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_1_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_1_io_uop_stale_pdst),
    .io_uop_exception(slots_1_io_uop_exception),
    .io_uop_exc_cause(slots_1_io_uop_exc_cause),
    .io_uop_bypassable(slots_1_io_uop_bypassable),
    .io_uop_mem_cmd(slots_1_io_uop_mem_cmd),
    .io_uop_mem_size(slots_1_io_uop_mem_size),
    .io_uop_mem_signed(slots_1_io_uop_mem_signed),
    .io_uop_is_fence(slots_1_io_uop_is_fence),
    .io_uop_is_fencei(slots_1_io_uop_is_fencei),
    .io_uop_is_amo(slots_1_io_uop_is_amo),
    .io_uop_uses_ldq(slots_1_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_1_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_1_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_1_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_1_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_1_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_1_io_uop_ldst),
    .io_uop_lrs1(slots_1_io_uop_lrs1),
    .io_uop_lrs2(slots_1_io_uop_lrs2),
    .io_uop_lrs3(slots_1_io_uop_lrs3),
    .io_uop_ldst_val(slots_1_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_1_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_1_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_1_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_1_io_uop_frs3_en),
    .io_uop_fp_val(slots_1_io_uop_fp_val),
    .io_uop_fp_single(slots_1_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_1_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_1_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_1_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_1_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_1_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_1_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_1_io_uop_debug_tsrc),
    .io_debug_p1(slots_1_io_debug_p1),
    .io_debug_p2(slots_1_io_debug_p2),
    .io_debug_p3(slots_1_io_debug_p3),
    .io_debug_ppred(slots_1_io_debug_ppred),
    .io_debug_state(slots_1_io_debug_state)
  );
  IssueSlot_16 slots_2 ( // @[issue-unit.scala 153:73]
    .clock(slots_2_clock),
    .reset(slots_2_reset),
    .io_valid(slots_2_io_valid),
    .io_will_be_valid(slots_2_io_will_be_valid),
    .io_request(slots_2_io_request),
    .io_request_hp(slots_2_io_request_hp),
    .io_grant(slots_2_io_grant),
    .io_brupdate_b1_resolve_mask(slots_2_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_2_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_uopc(slots_2_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_2_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_2_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_2_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_2_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_2_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_2_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_2_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_2_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_2_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_2_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_2_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_2_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_2_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_2_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_2_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_2_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_iw_state(slots_2_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_2_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_2_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_2_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_2_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_2_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_2_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_2_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_2_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_2_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_2_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_2_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_2_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_2_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_2_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_2_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_2_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_2_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_2_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_2_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_2_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_2_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_2_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_2_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_2_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_2_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_2_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_2_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_2_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_2_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_2_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_2_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_2_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_2_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_2_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_2_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_2_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_2_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_2_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_2_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_2_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_2_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_2_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_2_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_2_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_2_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_2_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_2_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_2_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_2_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_2_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_2_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_2_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_2_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_2_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_2_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_2_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_2_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_2_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_2_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_2_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_2_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_2_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_2_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_2_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_2_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_2_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_2_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_2_io_brupdate_b2_target_offset),
    .io_kill(slots_2_io_kill),
    .io_clear(slots_2_io_clear),
    .io_ldspec_miss(slots_2_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_2_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_2_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_2_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_1_valid(slots_2_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_2_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_2_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_2_valid(slots_2_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_2_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_2_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_3_valid(slots_2_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_2_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_2_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_4_valid(slots_2_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_2_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_2_io_wakeup_ports_4_bits_poisoned),
    .io_pred_wakeup_port_valid(slots_2_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_2_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_2_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_2_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_2_io_in_uop_valid),
    .io_in_uop_bits_uopc(slots_2_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_2_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_2_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_2_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_2_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_2_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_2_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_2_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_2_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_2_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_2_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_2_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_2_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_2_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_2_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_2_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_2_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_iw_state(slots_2_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_2_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_2_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_2_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_2_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_2_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_2_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_2_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_2_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_2_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_2_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_2_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_2_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_2_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_2_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_2_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_2_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_2_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_2_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_2_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_2_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_2_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_2_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_2_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_2_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_2_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_2_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_2_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_2_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_2_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_2_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_2_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_2_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_2_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_2_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_2_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_2_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_2_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_2_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_2_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_2_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_2_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_2_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_2_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_2_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_2_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_2_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_2_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_2_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_2_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_2_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_2_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_2_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_2_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_2_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_2_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_2_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_2_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_2_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_2_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_2_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_2_io_in_uop_bits_debug_tsrc),
    .io_out_uop_uopc(slots_2_io_out_uop_uopc),
    .io_out_uop_inst(slots_2_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_2_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_2_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_2_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_2_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_2_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_2_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_2_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_2_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_2_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_2_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_2_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_2_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_2_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_2_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_2_io_out_uop_ctrl_is_std),
    .io_out_uop_iw_state(slots_2_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_2_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_2_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_2_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_2_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_2_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_2_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_2_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_2_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_2_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_2_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_2_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_2_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_2_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_2_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_2_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_2_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_2_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_2_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_2_io_out_uop_pdst),
    .io_out_uop_prs1(slots_2_io_out_uop_prs1),
    .io_out_uop_prs2(slots_2_io_out_uop_prs2),
    .io_out_uop_prs3(slots_2_io_out_uop_prs3),
    .io_out_uop_ppred(slots_2_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_2_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_2_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_2_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_2_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_2_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_2_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_2_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_2_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_2_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_2_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_2_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_2_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_2_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_2_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_2_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_2_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_2_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_2_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_2_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_2_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_2_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_2_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_2_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_2_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_2_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_2_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_2_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_2_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_2_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_2_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_2_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_2_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_2_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_2_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_2_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_2_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_2_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_2_io_out_uop_debug_tsrc),
    .io_uop_uopc(slots_2_io_uop_uopc),
    .io_uop_inst(slots_2_io_uop_inst),
    .io_uop_debug_inst(slots_2_io_uop_debug_inst),
    .io_uop_is_rvc(slots_2_io_uop_is_rvc),
    .io_uop_debug_pc(slots_2_io_uop_debug_pc),
    .io_uop_iq_type(slots_2_io_uop_iq_type),
    .io_uop_fu_code(slots_2_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_2_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_2_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_2_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_2_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_2_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_2_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_2_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_2_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_2_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_2_io_uop_ctrl_is_std),
    .io_uop_iw_state(slots_2_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_2_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_2_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_2_io_uop_is_br),
    .io_uop_is_jalr(slots_2_io_uop_is_jalr),
    .io_uop_is_jal(slots_2_io_uop_is_jal),
    .io_uop_is_sfb(slots_2_io_uop_is_sfb),
    .io_uop_br_mask(slots_2_io_uop_br_mask),
    .io_uop_br_tag(slots_2_io_uop_br_tag),
    .io_uop_ftq_idx(slots_2_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_2_io_uop_edge_inst),
    .io_uop_pc_lob(slots_2_io_uop_pc_lob),
    .io_uop_taken(slots_2_io_uop_taken),
    .io_uop_imm_packed(slots_2_io_uop_imm_packed),
    .io_uop_csr_addr(slots_2_io_uop_csr_addr),
    .io_uop_rob_idx(slots_2_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_2_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_2_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_2_io_uop_rxq_idx),
    .io_uop_pdst(slots_2_io_uop_pdst),
    .io_uop_prs1(slots_2_io_uop_prs1),
    .io_uop_prs2(slots_2_io_uop_prs2),
    .io_uop_prs3(slots_2_io_uop_prs3),
    .io_uop_ppred(slots_2_io_uop_ppred),
    .io_uop_prs1_busy(slots_2_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_2_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_2_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_2_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_2_io_uop_stale_pdst),
    .io_uop_exception(slots_2_io_uop_exception),
    .io_uop_exc_cause(slots_2_io_uop_exc_cause),
    .io_uop_bypassable(slots_2_io_uop_bypassable),
    .io_uop_mem_cmd(slots_2_io_uop_mem_cmd),
    .io_uop_mem_size(slots_2_io_uop_mem_size),
    .io_uop_mem_signed(slots_2_io_uop_mem_signed),
    .io_uop_is_fence(slots_2_io_uop_is_fence),
    .io_uop_is_fencei(slots_2_io_uop_is_fencei),
    .io_uop_is_amo(slots_2_io_uop_is_amo),
    .io_uop_uses_ldq(slots_2_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_2_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_2_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_2_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_2_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_2_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_2_io_uop_ldst),
    .io_uop_lrs1(slots_2_io_uop_lrs1),
    .io_uop_lrs2(slots_2_io_uop_lrs2),
    .io_uop_lrs3(slots_2_io_uop_lrs3),
    .io_uop_ldst_val(slots_2_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_2_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_2_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_2_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_2_io_uop_frs3_en),
    .io_uop_fp_val(slots_2_io_uop_fp_val),
    .io_uop_fp_single(slots_2_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_2_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_2_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_2_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_2_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_2_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_2_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_2_io_uop_debug_tsrc),
    .io_debug_p1(slots_2_io_debug_p1),
    .io_debug_p2(slots_2_io_debug_p2),
    .io_debug_p3(slots_2_io_debug_p3),
    .io_debug_ppred(slots_2_io_debug_ppred),
    .io_debug_state(slots_2_io_debug_state)
  );
  IssueSlot_16 slots_3 ( // @[issue-unit.scala 153:73]
    .clock(slots_3_clock),
    .reset(slots_3_reset),
    .io_valid(slots_3_io_valid),
    .io_will_be_valid(slots_3_io_will_be_valid),
    .io_request(slots_3_io_request),
    .io_request_hp(slots_3_io_request_hp),
    .io_grant(slots_3_io_grant),
    .io_brupdate_b1_resolve_mask(slots_3_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_3_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_uopc(slots_3_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_3_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_3_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_3_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_3_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_3_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_3_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_3_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_3_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_3_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_3_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_3_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_3_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_3_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_3_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_3_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_3_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_iw_state(slots_3_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_3_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_3_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_3_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_3_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_3_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_3_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_3_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_3_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_3_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_3_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_3_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_3_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_3_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_3_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_3_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_3_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_3_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_3_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_3_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_3_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_3_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_3_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_3_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_3_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_3_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_3_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_3_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_3_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_3_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_3_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_3_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_3_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_3_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_3_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_3_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_3_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_3_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_3_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_3_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_3_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_3_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_3_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_3_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_3_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_3_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_3_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_3_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_3_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_3_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_3_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_3_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_3_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_3_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_3_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_3_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_3_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_3_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_3_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_3_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_3_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_3_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_3_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_3_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_3_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_3_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_3_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_3_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_3_io_brupdate_b2_target_offset),
    .io_kill(slots_3_io_kill),
    .io_clear(slots_3_io_clear),
    .io_ldspec_miss(slots_3_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_3_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_3_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_3_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_1_valid(slots_3_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_3_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_3_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_2_valid(slots_3_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_3_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_3_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_3_valid(slots_3_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_3_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_3_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_4_valid(slots_3_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_3_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_3_io_wakeup_ports_4_bits_poisoned),
    .io_pred_wakeup_port_valid(slots_3_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_3_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_3_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_3_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_3_io_in_uop_valid),
    .io_in_uop_bits_uopc(slots_3_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_3_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_3_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_3_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_3_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_3_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_3_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_3_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_3_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_3_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_3_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_3_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_3_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_3_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_3_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_3_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_3_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_iw_state(slots_3_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_3_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_3_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_3_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_3_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_3_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_3_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_3_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_3_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_3_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_3_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_3_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_3_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_3_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_3_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_3_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_3_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_3_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_3_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_3_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_3_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_3_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_3_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_3_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_3_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_3_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_3_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_3_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_3_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_3_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_3_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_3_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_3_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_3_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_3_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_3_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_3_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_3_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_3_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_3_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_3_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_3_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_3_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_3_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_3_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_3_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_3_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_3_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_3_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_3_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_3_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_3_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_3_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_3_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_3_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_3_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_3_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_3_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_3_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_3_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_3_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_3_io_in_uop_bits_debug_tsrc),
    .io_out_uop_uopc(slots_3_io_out_uop_uopc),
    .io_out_uop_inst(slots_3_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_3_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_3_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_3_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_3_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_3_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_3_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_3_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_3_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_3_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_3_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_3_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_3_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_3_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_3_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_3_io_out_uop_ctrl_is_std),
    .io_out_uop_iw_state(slots_3_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_3_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_3_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_3_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_3_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_3_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_3_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_3_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_3_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_3_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_3_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_3_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_3_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_3_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_3_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_3_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_3_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_3_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_3_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_3_io_out_uop_pdst),
    .io_out_uop_prs1(slots_3_io_out_uop_prs1),
    .io_out_uop_prs2(slots_3_io_out_uop_prs2),
    .io_out_uop_prs3(slots_3_io_out_uop_prs3),
    .io_out_uop_ppred(slots_3_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_3_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_3_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_3_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_3_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_3_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_3_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_3_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_3_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_3_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_3_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_3_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_3_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_3_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_3_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_3_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_3_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_3_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_3_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_3_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_3_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_3_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_3_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_3_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_3_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_3_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_3_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_3_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_3_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_3_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_3_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_3_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_3_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_3_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_3_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_3_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_3_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_3_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_3_io_out_uop_debug_tsrc),
    .io_uop_uopc(slots_3_io_uop_uopc),
    .io_uop_inst(slots_3_io_uop_inst),
    .io_uop_debug_inst(slots_3_io_uop_debug_inst),
    .io_uop_is_rvc(slots_3_io_uop_is_rvc),
    .io_uop_debug_pc(slots_3_io_uop_debug_pc),
    .io_uop_iq_type(slots_3_io_uop_iq_type),
    .io_uop_fu_code(slots_3_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_3_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_3_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_3_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_3_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_3_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_3_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_3_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_3_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_3_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_3_io_uop_ctrl_is_std),
    .io_uop_iw_state(slots_3_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_3_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_3_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_3_io_uop_is_br),
    .io_uop_is_jalr(slots_3_io_uop_is_jalr),
    .io_uop_is_jal(slots_3_io_uop_is_jal),
    .io_uop_is_sfb(slots_3_io_uop_is_sfb),
    .io_uop_br_mask(slots_3_io_uop_br_mask),
    .io_uop_br_tag(slots_3_io_uop_br_tag),
    .io_uop_ftq_idx(slots_3_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_3_io_uop_edge_inst),
    .io_uop_pc_lob(slots_3_io_uop_pc_lob),
    .io_uop_taken(slots_3_io_uop_taken),
    .io_uop_imm_packed(slots_3_io_uop_imm_packed),
    .io_uop_csr_addr(slots_3_io_uop_csr_addr),
    .io_uop_rob_idx(slots_3_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_3_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_3_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_3_io_uop_rxq_idx),
    .io_uop_pdst(slots_3_io_uop_pdst),
    .io_uop_prs1(slots_3_io_uop_prs1),
    .io_uop_prs2(slots_3_io_uop_prs2),
    .io_uop_prs3(slots_3_io_uop_prs3),
    .io_uop_ppred(slots_3_io_uop_ppred),
    .io_uop_prs1_busy(slots_3_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_3_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_3_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_3_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_3_io_uop_stale_pdst),
    .io_uop_exception(slots_3_io_uop_exception),
    .io_uop_exc_cause(slots_3_io_uop_exc_cause),
    .io_uop_bypassable(slots_3_io_uop_bypassable),
    .io_uop_mem_cmd(slots_3_io_uop_mem_cmd),
    .io_uop_mem_size(slots_3_io_uop_mem_size),
    .io_uop_mem_signed(slots_3_io_uop_mem_signed),
    .io_uop_is_fence(slots_3_io_uop_is_fence),
    .io_uop_is_fencei(slots_3_io_uop_is_fencei),
    .io_uop_is_amo(slots_3_io_uop_is_amo),
    .io_uop_uses_ldq(slots_3_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_3_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_3_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_3_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_3_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_3_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_3_io_uop_ldst),
    .io_uop_lrs1(slots_3_io_uop_lrs1),
    .io_uop_lrs2(slots_3_io_uop_lrs2),
    .io_uop_lrs3(slots_3_io_uop_lrs3),
    .io_uop_ldst_val(slots_3_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_3_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_3_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_3_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_3_io_uop_frs3_en),
    .io_uop_fp_val(slots_3_io_uop_fp_val),
    .io_uop_fp_single(slots_3_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_3_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_3_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_3_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_3_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_3_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_3_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_3_io_uop_debug_tsrc),
    .io_debug_p1(slots_3_io_debug_p1),
    .io_debug_p2(slots_3_io_debug_p2),
    .io_debug_p3(slots_3_io_debug_p3),
    .io_debug_ppred(slots_3_io_debug_ppred),
    .io_debug_state(slots_3_io_debug_state)
  );
  IssueSlot_16 slots_4 ( // @[issue-unit.scala 153:73]
    .clock(slots_4_clock),
    .reset(slots_4_reset),
    .io_valid(slots_4_io_valid),
    .io_will_be_valid(slots_4_io_will_be_valid),
    .io_request(slots_4_io_request),
    .io_request_hp(slots_4_io_request_hp),
    .io_grant(slots_4_io_grant),
    .io_brupdate_b1_resolve_mask(slots_4_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_4_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_uopc(slots_4_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_4_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_4_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_4_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_4_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_4_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_4_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_4_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_4_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_4_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_4_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_4_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_4_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_4_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_4_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_4_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_4_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_iw_state(slots_4_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_4_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_4_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_4_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_4_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_4_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_4_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_4_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_4_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_4_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_4_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_4_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_4_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_4_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_4_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_4_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_4_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_4_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_4_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_4_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_4_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_4_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_4_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_4_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_4_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_4_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_4_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_4_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_4_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_4_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_4_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_4_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_4_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_4_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_4_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_4_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_4_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_4_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_4_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_4_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_4_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_4_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_4_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_4_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_4_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_4_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_4_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_4_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_4_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_4_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_4_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_4_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_4_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_4_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_4_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_4_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_4_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_4_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_4_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_4_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_4_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_4_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_4_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_4_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_4_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_4_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_4_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_4_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_4_io_brupdate_b2_target_offset),
    .io_kill(slots_4_io_kill),
    .io_clear(slots_4_io_clear),
    .io_ldspec_miss(slots_4_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_4_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_4_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_4_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_1_valid(slots_4_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_4_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_4_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_2_valid(slots_4_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_4_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_4_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_3_valid(slots_4_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_4_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_4_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_4_valid(slots_4_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_4_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_4_io_wakeup_ports_4_bits_poisoned),
    .io_pred_wakeup_port_valid(slots_4_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_4_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_4_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_4_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_4_io_in_uop_valid),
    .io_in_uop_bits_uopc(slots_4_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_4_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_4_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_4_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_4_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_4_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_4_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_4_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_4_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_4_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_4_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_4_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_4_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_4_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_4_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_4_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_4_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_iw_state(slots_4_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_4_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_4_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_4_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_4_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_4_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_4_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_4_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_4_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_4_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_4_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_4_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_4_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_4_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_4_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_4_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_4_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_4_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_4_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_4_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_4_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_4_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_4_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_4_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_4_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_4_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_4_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_4_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_4_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_4_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_4_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_4_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_4_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_4_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_4_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_4_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_4_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_4_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_4_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_4_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_4_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_4_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_4_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_4_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_4_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_4_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_4_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_4_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_4_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_4_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_4_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_4_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_4_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_4_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_4_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_4_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_4_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_4_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_4_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_4_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_4_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_4_io_in_uop_bits_debug_tsrc),
    .io_out_uop_uopc(slots_4_io_out_uop_uopc),
    .io_out_uop_inst(slots_4_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_4_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_4_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_4_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_4_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_4_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_4_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_4_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_4_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_4_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_4_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_4_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_4_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_4_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_4_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_4_io_out_uop_ctrl_is_std),
    .io_out_uop_iw_state(slots_4_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_4_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_4_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_4_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_4_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_4_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_4_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_4_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_4_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_4_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_4_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_4_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_4_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_4_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_4_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_4_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_4_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_4_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_4_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_4_io_out_uop_pdst),
    .io_out_uop_prs1(slots_4_io_out_uop_prs1),
    .io_out_uop_prs2(slots_4_io_out_uop_prs2),
    .io_out_uop_prs3(slots_4_io_out_uop_prs3),
    .io_out_uop_ppred(slots_4_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_4_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_4_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_4_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_4_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_4_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_4_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_4_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_4_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_4_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_4_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_4_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_4_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_4_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_4_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_4_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_4_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_4_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_4_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_4_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_4_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_4_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_4_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_4_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_4_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_4_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_4_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_4_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_4_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_4_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_4_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_4_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_4_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_4_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_4_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_4_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_4_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_4_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_4_io_out_uop_debug_tsrc),
    .io_uop_uopc(slots_4_io_uop_uopc),
    .io_uop_inst(slots_4_io_uop_inst),
    .io_uop_debug_inst(slots_4_io_uop_debug_inst),
    .io_uop_is_rvc(slots_4_io_uop_is_rvc),
    .io_uop_debug_pc(slots_4_io_uop_debug_pc),
    .io_uop_iq_type(slots_4_io_uop_iq_type),
    .io_uop_fu_code(slots_4_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_4_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_4_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_4_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_4_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_4_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_4_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_4_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_4_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_4_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_4_io_uop_ctrl_is_std),
    .io_uop_iw_state(slots_4_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_4_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_4_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_4_io_uop_is_br),
    .io_uop_is_jalr(slots_4_io_uop_is_jalr),
    .io_uop_is_jal(slots_4_io_uop_is_jal),
    .io_uop_is_sfb(slots_4_io_uop_is_sfb),
    .io_uop_br_mask(slots_4_io_uop_br_mask),
    .io_uop_br_tag(slots_4_io_uop_br_tag),
    .io_uop_ftq_idx(slots_4_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_4_io_uop_edge_inst),
    .io_uop_pc_lob(slots_4_io_uop_pc_lob),
    .io_uop_taken(slots_4_io_uop_taken),
    .io_uop_imm_packed(slots_4_io_uop_imm_packed),
    .io_uop_csr_addr(slots_4_io_uop_csr_addr),
    .io_uop_rob_idx(slots_4_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_4_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_4_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_4_io_uop_rxq_idx),
    .io_uop_pdst(slots_4_io_uop_pdst),
    .io_uop_prs1(slots_4_io_uop_prs1),
    .io_uop_prs2(slots_4_io_uop_prs2),
    .io_uop_prs3(slots_4_io_uop_prs3),
    .io_uop_ppred(slots_4_io_uop_ppred),
    .io_uop_prs1_busy(slots_4_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_4_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_4_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_4_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_4_io_uop_stale_pdst),
    .io_uop_exception(slots_4_io_uop_exception),
    .io_uop_exc_cause(slots_4_io_uop_exc_cause),
    .io_uop_bypassable(slots_4_io_uop_bypassable),
    .io_uop_mem_cmd(slots_4_io_uop_mem_cmd),
    .io_uop_mem_size(slots_4_io_uop_mem_size),
    .io_uop_mem_signed(slots_4_io_uop_mem_signed),
    .io_uop_is_fence(slots_4_io_uop_is_fence),
    .io_uop_is_fencei(slots_4_io_uop_is_fencei),
    .io_uop_is_amo(slots_4_io_uop_is_amo),
    .io_uop_uses_ldq(slots_4_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_4_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_4_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_4_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_4_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_4_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_4_io_uop_ldst),
    .io_uop_lrs1(slots_4_io_uop_lrs1),
    .io_uop_lrs2(slots_4_io_uop_lrs2),
    .io_uop_lrs3(slots_4_io_uop_lrs3),
    .io_uop_ldst_val(slots_4_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_4_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_4_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_4_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_4_io_uop_frs3_en),
    .io_uop_fp_val(slots_4_io_uop_fp_val),
    .io_uop_fp_single(slots_4_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_4_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_4_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_4_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_4_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_4_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_4_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_4_io_uop_debug_tsrc),
    .io_debug_p1(slots_4_io_debug_p1),
    .io_debug_p2(slots_4_io_debug_p2),
    .io_debug_p3(slots_4_io_debug_p3),
    .io_debug_ppred(slots_4_io_debug_ppred),
    .io_debug_state(slots_4_io_debug_state)
  );
  IssueSlot_16 slots_5 ( // @[issue-unit.scala 153:73]
    .clock(slots_5_clock),
    .reset(slots_5_reset),
    .io_valid(slots_5_io_valid),
    .io_will_be_valid(slots_5_io_will_be_valid),
    .io_request(slots_5_io_request),
    .io_request_hp(slots_5_io_request_hp),
    .io_grant(slots_5_io_grant),
    .io_brupdate_b1_resolve_mask(slots_5_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_5_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_uopc(slots_5_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_5_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_5_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_5_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_5_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_5_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_5_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_5_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_5_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_5_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_5_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_5_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_5_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_5_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_5_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_5_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_5_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_iw_state(slots_5_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_5_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_5_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_5_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_5_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_5_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_5_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_5_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_5_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_5_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_5_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_5_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_5_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_5_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_5_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_5_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_5_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_5_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_5_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_5_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_5_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_5_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_5_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_5_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_5_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_5_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_5_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_5_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_5_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_5_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_5_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_5_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_5_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_5_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_5_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_5_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_5_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_5_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_5_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_5_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_5_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_5_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_5_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_5_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_5_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_5_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_5_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_5_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_5_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_5_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_5_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_5_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_5_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_5_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_5_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_5_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_5_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_5_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_5_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_5_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_5_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_5_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_5_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_5_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_5_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_5_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_5_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_5_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_5_io_brupdate_b2_target_offset),
    .io_kill(slots_5_io_kill),
    .io_clear(slots_5_io_clear),
    .io_ldspec_miss(slots_5_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_5_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_5_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_5_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_1_valid(slots_5_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_5_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_5_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_2_valid(slots_5_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_5_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_5_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_3_valid(slots_5_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_5_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_5_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_4_valid(slots_5_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_5_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_5_io_wakeup_ports_4_bits_poisoned),
    .io_pred_wakeup_port_valid(slots_5_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_5_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_5_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_5_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_5_io_in_uop_valid),
    .io_in_uop_bits_uopc(slots_5_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_5_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_5_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_5_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_5_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_5_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_5_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_5_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_5_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_5_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_5_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_5_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_5_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_5_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_5_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_5_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_5_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_iw_state(slots_5_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_5_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_5_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_5_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_5_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_5_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_5_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_5_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_5_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_5_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_5_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_5_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_5_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_5_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_5_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_5_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_5_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_5_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_5_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_5_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_5_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_5_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_5_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_5_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_5_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_5_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_5_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_5_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_5_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_5_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_5_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_5_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_5_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_5_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_5_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_5_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_5_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_5_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_5_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_5_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_5_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_5_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_5_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_5_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_5_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_5_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_5_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_5_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_5_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_5_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_5_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_5_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_5_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_5_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_5_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_5_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_5_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_5_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_5_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_5_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_5_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_5_io_in_uop_bits_debug_tsrc),
    .io_out_uop_uopc(slots_5_io_out_uop_uopc),
    .io_out_uop_inst(slots_5_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_5_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_5_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_5_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_5_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_5_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_5_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_5_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_5_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_5_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_5_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_5_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_5_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_5_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_5_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_5_io_out_uop_ctrl_is_std),
    .io_out_uop_iw_state(slots_5_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_5_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_5_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_5_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_5_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_5_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_5_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_5_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_5_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_5_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_5_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_5_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_5_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_5_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_5_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_5_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_5_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_5_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_5_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_5_io_out_uop_pdst),
    .io_out_uop_prs1(slots_5_io_out_uop_prs1),
    .io_out_uop_prs2(slots_5_io_out_uop_prs2),
    .io_out_uop_prs3(slots_5_io_out_uop_prs3),
    .io_out_uop_ppred(slots_5_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_5_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_5_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_5_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_5_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_5_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_5_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_5_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_5_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_5_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_5_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_5_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_5_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_5_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_5_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_5_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_5_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_5_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_5_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_5_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_5_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_5_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_5_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_5_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_5_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_5_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_5_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_5_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_5_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_5_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_5_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_5_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_5_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_5_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_5_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_5_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_5_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_5_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_5_io_out_uop_debug_tsrc),
    .io_uop_uopc(slots_5_io_uop_uopc),
    .io_uop_inst(slots_5_io_uop_inst),
    .io_uop_debug_inst(slots_5_io_uop_debug_inst),
    .io_uop_is_rvc(slots_5_io_uop_is_rvc),
    .io_uop_debug_pc(slots_5_io_uop_debug_pc),
    .io_uop_iq_type(slots_5_io_uop_iq_type),
    .io_uop_fu_code(slots_5_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_5_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_5_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_5_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_5_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_5_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_5_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_5_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_5_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_5_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_5_io_uop_ctrl_is_std),
    .io_uop_iw_state(slots_5_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_5_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_5_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_5_io_uop_is_br),
    .io_uop_is_jalr(slots_5_io_uop_is_jalr),
    .io_uop_is_jal(slots_5_io_uop_is_jal),
    .io_uop_is_sfb(slots_5_io_uop_is_sfb),
    .io_uop_br_mask(slots_5_io_uop_br_mask),
    .io_uop_br_tag(slots_5_io_uop_br_tag),
    .io_uop_ftq_idx(slots_5_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_5_io_uop_edge_inst),
    .io_uop_pc_lob(slots_5_io_uop_pc_lob),
    .io_uop_taken(slots_5_io_uop_taken),
    .io_uop_imm_packed(slots_5_io_uop_imm_packed),
    .io_uop_csr_addr(slots_5_io_uop_csr_addr),
    .io_uop_rob_idx(slots_5_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_5_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_5_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_5_io_uop_rxq_idx),
    .io_uop_pdst(slots_5_io_uop_pdst),
    .io_uop_prs1(slots_5_io_uop_prs1),
    .io_uop_prs2(slots_5_io_uop_prs2),
    .io_uop_prs3(slots_5_io_uop_prs3),
    .io_uop_ppred(slots_5_io_uop_ppred),
    .io_uop_prs1_busy(slots_5_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_5_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_5_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_5_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_5_io_uop_stale_pdst),
    .io_uop_exception(slots_5_io_uop_exception),
    .io_uop_exc_cause(slots_5_io_uop_exc_cause),
    .io_uop_bypassable(slots_5_io_uop_bypassable),
    .io_uop_mem_cmd(slots_5_io_uop_mem_cmd),
    .io_uop_mem_size(slots_5_io_uop_mem_size),
    .io_uop_mem_signed(slots_5_io_uop_mem_signed),
    .io_uop_is_fence(slots_5_io_uop_is_fence),
    .io_uop_is_fencei(slots_5_io_uop_is_fencei),
    .io_uop_is_amo(slots_5_io_uop_is_amo),
    .io_uop_uses_ldq(slots_5_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_5_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_5_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_5_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_5_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_5_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_5_io_uop_ldst),
    .io_uop_lrs1(slots_5_io_uop_lrs1),
    .io_uop_lrs2(slots_5_io_uop_lrs2),
    .io_uop_lrs3(slots_5_io_uop_lrs3),
    .io_uop_ldst_val(slots_5_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_5_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_5_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_5_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_5_io_uop_frs3_en),
    .io_uop_fp_val(slots_5_io_uop_fp_val),
    .io_uop_fp_single(slots_5_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_5_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_5_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_5_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_5_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_5_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_5_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_5_io_uop_debug_tsrc),
    .io_debug_p1(slots_5_io_debug_p1),
    .io_debug_p2(slots_5_io_debug_p2),
    .io_debug_p3(slots_5_io_debug_p3),
    .io_debug_ppred(slots_5_io_debug_ppred),
    .io_debug_state(slots_5_io_debug_state)
  );
  IssueSlot_16 slots_6 ( // @[issue-unit.scala 153:73]
    .clock(slots_6_clock),
    .reset(slots_6_reset),
    .io_valid(slots_6_io_valid),
    .io_will_be_valid(slots_6_io_will_be_valid),
    .io_request(slots_6_io_request),
    .io_request_hp(slots_6_io_request_hp),
    .io_grant(slots_6_io_grant),
    .io_brupdate_b1_resolve_mask(slots_6_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_6_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_uopc(slots_6_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_6_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_6_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_6_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_6_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_6_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_6_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_6_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_6_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_6_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_6_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_6_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_6_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_6_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_6_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_6_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_6_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_iw_state(slots_6_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_6_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_6_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_6_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_6_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_6_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_6_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_6_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_6_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_6_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_6_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_6_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_6_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_6_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_6_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_6_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_6_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_6_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_6_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_6_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_6_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_6_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_6_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_6_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_6_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_6_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_6_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_6_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_6_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_6_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_6_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_6_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_6_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_6_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_6_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_6_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_6_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_6_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_6_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_6_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_6_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_6_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_6_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_6_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_6_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_6_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_6_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_6_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_6_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_6_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_6_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_6_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_6_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_6_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_6_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_6_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_6_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_6_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_6_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_6_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_6_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_6_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_6_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_6_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_6_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_6_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_6_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_6_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_6_io_brupdate_b2_target_offset),
    .io_kill(slots_6_io_kill),
    .io_clear(slots_6_io_clear),
    .io_ldspec_miss(slots_6_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_6_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_6_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_6_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_1_valid(slots_6_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_6_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_6_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_2_valid(slots_6_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_6_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_6_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_3_valid(slots_6_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_6_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_6_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_4_valid(slots_6_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_6_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_6_io_wakeup_ports_4_bits_poisoned),
    .io_pred_wakeup_port_valid(slots_6_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_6_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_6_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_6_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_6_io_in_uop_valid),
    .io_in_uop_bits_uopc(slots_6_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_6_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_6_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_6_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_6_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_6_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_6_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_6_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_6_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_6_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_6_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_6_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_6_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_6_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_6_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_6_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_6_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_iw_state(slots_6_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_6_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_6_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_6_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_6_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_6_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_6_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_6_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_6_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_6_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_6_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_6_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_6_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_6_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_6_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_6_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_6_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_6_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_6_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_6_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_6_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_6_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_6_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_6_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_6_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_6_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_6_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_6_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_6_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_6_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_6_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_6_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_6_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_6_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_6_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_6_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_6_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_6_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_6_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_6_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_6_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_6_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_6_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_6_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_6_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_6_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_6_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_6_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_6_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_6_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_6_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_6_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_6_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_6_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_6_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_6_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_6_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_6_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_6_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_6_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_6_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_6_io_in_uop_bits_debug_tsrc),
    .io_out_uop_uopc(slots_6_io_out_uop_uopc),
    .io_out_uop_inst(slots_6_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_6_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_6_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_6_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_6_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_6_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_6_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_6_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_6_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_6_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_6_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_6_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_6_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_6_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_6_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_6_io_out_uop_ctrl_is_std),
    .io_out_uop_iw_state(slots_6_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_6_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_6_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_6_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_6_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_6_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_6_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_6_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_6_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_6_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_6_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_6_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_6_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_6_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_6_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_6_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_6_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_6_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_6_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_6_io_out_uop_pdst),
    .io_out_uop_prs1(slots_6_io_out_uop_prs1),
    .io_out_uop_prs2(slots_6_io_out_uop_prs2),
    .io_out_uop_prs3(slots_6_io_out_uop_prs3),
    .io_out_uop_ppred(slots_6_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_6_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_6_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_6_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_6_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_6_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_6_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_6_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_6_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_6_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_6_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_6_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_6_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_6_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_6_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_6_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_6_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_6_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_6_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_6_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_6_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_6_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_6_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_6_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_6_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_6_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_6_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_6_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_6_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_6_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_6_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_6_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_6_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_6_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_6_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_6_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_6_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_6_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_6_io_out_uop_debug_tsrc),
    .io_uop_uopc(slots_6_io_uop_uopc),
    .io_uop_inst(slots_6_io_uop_inst),
    .io_uop_debug_inst(slots_6_io_uop_debug_inst),
    .io_uop_is_rvc(slots_6_io_uop_is_rvc),
    .io_uop_debug_pc(slots_6_io_uop_debug_pc),
    .io_uop_iq_type(slots_6_io_uop_iq_type),
    .io_uop_fu_code(slots_6_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_6_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_6_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_6_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_6_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_6_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_6_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_6_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_6_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_6_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_6_io_uop_ctrl_is_std),
    .io_uop_iw_state(slots_6_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_6_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_6_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_6_io_uop_is_br),
    .io_uop_is_jalr(slots_6_io_uop_is_jalr),
    .io_uop_is_jal(slots_6_io_uop_is_jal),
    .io_uop_is_sfb(slots_6_io_uop_is_sfb),
    .io_uop_br_mask(slots_6_io_uop_br_mask),
    .io_uop_br_tag(slots_6_io_uop_br_tag),
    .io_uop_ftq_idx(slots_6_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_6_io_uop_edge_inst),
    .io_uop_pc_lob(slots_6_io_uop_pc_lob),
    .io_uop_taken(slots_6_io_uop_taken),
    .io_uop_imm_packed(slots_6_io_uop_imm_packed),
    .io_uop_csr_addr(slots_6_io_uop_csr_addr),
    .io_uop_rob_idx(slots_6_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_6_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_6_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_6_io_uop_rxq_idx),
    .io_uop_pdst(slots_6_io_uop_pdst),
    .io_uop_prs1(slots_6_io_uop_prs1),
    .io_uop_prs2(slots_6_io_uop_prs2),
    .io_uop_prs3(slots_6_io_uop_prs3),
    .io_uop_ppred(slots_6_io_uop_ppred),
    .io_uop_prs1_busy(slots_6_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_6_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_6_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_6_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_6_io_uop_stale_pdst),
    .io_uop_exception(slots_6_io_uop_exception),
    .io_uop_exc_cause(slots_6_io_uop_exc_cause),
    .io_uop_bypassable(slots_6_io_uop_bypassable),
    .io_uop_mem_cmd(slots_6_io_uop_mem_cmd),
    .io_uop_mem_size(slots_6_io_uop_mem_size),
    .io_uop_mem_signed(slots_6_io_uop_mem_signed),
    .io_uop_is_fence(slots_6_io_uop_is_fence),
    .io_uop_is_fencei(slots_6_io_uop_is_fencei),
    .io_uop_is_amo(slots_6_io_uop_is_amo),
    .io_uop_uses_ldq(slots_6_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_6_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_6_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_6_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_6_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_6_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_6_io_uop_ldst),
    .io_uop_lrs1(slots_6_io_uop_lrs1),
    .io_uop_lrs2(slots_6_io_uop_lrs2),
    .io_uop_lrs3(slots_6_io_uop_lrs3),
    .io_uop_ldst_val(slots_6_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_6_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_6_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_6_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_6_io_uop_frs3_en),
    .io_uop_fp_val(slots_6_io_uop_fp_val),
    .io_uop_fp_single(slots_6_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_6_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_6_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_6_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_6_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_6_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_6_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_6_io_uop_debug_tsrc),
    .io_debug_p1(slots_6_io_debug_p1),
    .io_debug_p2(slots_6_io_debug_p2),
    .io_debug_p3(slots_6_io_debug_p3),
    .io_debug_ppred(slots_6_io_debug_ppred),
    .io_debug_state(slots_6_io_debug_state)
  );
  IssueSlot_16 slots_7 ( // @[issue-unit.scala 153:73]
    .clock(slots_7_clock),
    .reset(slots_7_reset),
    .io_valid(slots_7_io_valid),
    .io_will_be_valid(slots_7_io_will_be_valid),
    .io_request(slots_7_io_request),
    .io_request_hp(slots_7_io_request_hp),
    .io_grant(slots_7_io_grant),
    .io_brupdate_b1_resolve_mask(slots_7_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_7_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_uopc(slots_7_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_7_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_7_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_7_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_7_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_7_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_7_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_7_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_7_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_7_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_7_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_7_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_7_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_7_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_7_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_7_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_7_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_iw_state(slots_7_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_7_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_7_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_7_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_7_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_7_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_7_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_7_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_7_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_7_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_7_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_7_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_7_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_7_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_7_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_7_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_7_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_7_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_7_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_7_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_7_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_7_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_7_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_7_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_7_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_7_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_7_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_7_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_7_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_7_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_7_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_7_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_7_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_7_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_7_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_7_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_7_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_7_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_7_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_7_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_7_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_7_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_7_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_7_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_7_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_7_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_7_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_7_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_7_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_7_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_7_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_7_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_7_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_7_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_7_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_7_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_7_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_7_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_7_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_7_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_7_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_7_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_7_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_7_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_7_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_7_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_7_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_7_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_7_io_brupdate_b2_target_offset),
    .io_kill(slots_7_io_kill),
    .io_clear(slots_7_io_clear),
    .io_ldspec_miss(slots_7_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_7_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_7_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_7_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_1_valid(slots_7_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_7_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_7_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_2_valid(slots_7_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_7_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_7_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_3_valid(slots_7_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_7_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_7_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_4_valid(slots_7_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_7_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_7_io_wakeup_ports_4_bits_poisoned),
    .io_pred_wakeup_port_valid(slots_7_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_7_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_7_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_7_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_7_io_in_uop_valid),
    .io_in_uop_bits_uopc(slots_7_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_7_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_7_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_7_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_7_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_7_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_7_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_7_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_7_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_7_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_7_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_7_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_7_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_7_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_7_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_7_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_7_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_iw_state(slots_7_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_7_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_7_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_7_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_7_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_7_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_7_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_7_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_7_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_7_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_7_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_7_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_7_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_7_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_7_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_7_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_7_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_7_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_7_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_7_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_7_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_7_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_7_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_7_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_7_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_7_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_7_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_7_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_7_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_7_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_7_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_7_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_7_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_7_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_7_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_7_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_7_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_7_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_7_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_7_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_7_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_7_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_7_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_7_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_7_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_7_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_7_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_7_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_7_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_7_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_7_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_7_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_7_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_7_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_7_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_7_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_7_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_7_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_7_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_7_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_7_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_7_io_in_uop_bits_debug_tsrc),
    .io_out_uop_uopc(slots_7_io_out_uop_uopc),
    .io_out_uop_inst(slots_7_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_7_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_7_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_7_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_7_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_7_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_7_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_7_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_7_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_7_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_7_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_7_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_7_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_7_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_7_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_7_io_out_uop_ctrl_is_std),
    .io_out_uop_iw_state(slots_7_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_7_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_7_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_7_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_7_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_7_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_7_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_7_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_7_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_7_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_7_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_7_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_7_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_7_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_7_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_7_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_7_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_7_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_7_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_7_io_out_uop_pdst),
    .io_out_uop_prs1(slots_7_io_out_uop_prs1),
    .io_out_uop_prs2(slots_7_io_out_uop_prs2),
    .io_out_uop_prs3(slots_7_io_out_uop_prs3),
    .io_out_uop_ppred(slots_7_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_7_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_7_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_7_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_7_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_7_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_7_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_7_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_7_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_7_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_7_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_7_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_7_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_7_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_7_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_7_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_7_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_7_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_7_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_7_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_7_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_7_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_7_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_7_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_7_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_7_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_7_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_7_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_7_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_7_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_7_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_7_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_7_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_7_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_7_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_7_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_7_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_7_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_7_io_out_uop_debug_tsrc),
    .io_uop_uopc(slots_7_io_uop_uopc),
    .io_uop_inst(slots_7_io_uop_inst),
    .io_uop_debug_inst(slots_7_io_uop_debug_inst),
    .io_uop_is_rvc(slots_7_io_uop_is_rvc),
    .io_uop_debug_pc(slots_7_io_uop_debug_pc),
    .io_uop_iq_type(slots_7_io_uop_iq_type),
    .io_uop_fu_code(slots_7_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_7_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_7_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_7_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_7_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_7_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_7_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_7_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_7_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_7_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_7_io_uop_ctrl_is_std),
    .io_uop_iw_state(slots_7_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_7_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_7_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_7_io_uop_is_br),
    .io_uop_is_jalr(slots_7_io_uop_is_jalr),
    .io_uop_is_jal(slots_7_io_uop_is_jal),
    .io_uop_is_sfb(slots_7_io_uop_is_sfb),
    .io_uop_br_mask(slots_7_io_uop_br_mask),
    .io_uop_br_tag(slots_7_io_uop_br_tag),
    .io_uop_ftq_idx(slots_7_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_7_io_uop_edge_inst),
    .io_uop_pc_lob(slots_7_io_uop_pc_lob),
    .io_uop_taken(slots_7_io_uop_taken),
    .io_uop_imm_packed(slots_7_io_uop_imm_packed),
    .io_uop_csr_addr(slots_7_io_uop_csr_addr),
    .io_uop_rob_idx(slots_7_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_7_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_7_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_7_io_uop_rxq_idx),
    .io_uop_pdst(slots_7_io_uop_pdst),
    .io_uop_prs1(slots_7_io_uop_prs1),
    .io_uop_prs2(slots_7_io_uop_prs2),
    .io_uop_prs3(slots_7_io_uop_prs3),
    .io_uop_ppred(slots_7_io_uop_ppred),
    .io_uop_prs1_busy(slots_7_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_7_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_7_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_7_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_7_io_uop_stale_pdst),
    .io_uop_exception(slots_7_io_uop_exception),
    .io_uop_exc_cause(slots_7_io_uop_exc_cause),
    .io_uop_bypassable(slots_7_io_uop_bypassable),
    .io_uop_mem_cmd(slots_7_io_uop_mem_cmd),
    .io_uop_mem_size(slots_7_io_uop_mem_size),
    .io_uop_mem_signed(slots_7_io_uop_mem_signed),
    .io_uop_is_fence(slots_7_io_uop_is_fence),
    .io_uop_is_fencei(slots_7_io_uop_is_fencei),
    .io_uop_is_amo(slots_7_io_uop_is_amo),
    .io_uop_uses_ldq(slots_7_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_7_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_7_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_7_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_7_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_7_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_7_io_uop_ldst),
    .io_uop_lrs1(slots_7_io_uop_lrs1),
    .io_uop_lrs2(slots_7_io_uop_lrs2),
    .io_uop_lrs3(slots_7_io_uop_lrs3),
    .io_uop_ldst_val(slots_7_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_7_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_7_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_7_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_7_io_uop_frs3_en),
    .io_uop_fp_val(slots_7_io_uop_fp_val),
    .io_uop_fp_single(slots_7_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_7_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_7_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_7_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_7_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_7_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_7_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_7_io_uop_debug_tsrc),
    .io_debug_p1(slots_7_io_debug_p1),
    .io_debug_p2(slots_7_io_debug_p2),
    .io_debug_p3(slots_7_io_debug_p3),
    .io_debug_ppred(slots_7_io_debug_ppred),
    .io_debug_state(slots_7_io_debug_state)
  );
  IssueSlot_16 slots_8 ( // @[issue-unit.scala 153:73]
    .clock(slots_8_clock),
    .reset(slots_8_reset),
    .io_valid(slots_8_io_valid),
    .io_will_be_valid(slots_8_io_will_be_valid),
    .io_request(slots_8_io_request),
    .io_request_hp(slots_8_io_request_hp),
    .io_grant(slots_8_io_grant),
    .io_brupdate_b1_resolve_mask(slots_8_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_8_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_uopc(slots_8_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_8_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_8_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_8_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_8_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_8_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_8_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_8_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_8_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_8_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_8_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_8_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_8_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_8_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_8_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_8_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_8_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_iw_state(slots_8_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_8_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_8_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_8_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_8_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_8_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_8_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_8_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_8_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_8_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_8_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_8_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_8_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_8_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_8_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_8_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_8_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_8_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_8_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_8_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_8_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_8_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_8_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_8_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_8_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_8_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_8_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_8_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_8_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_8_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_8_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_8_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_8_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_8_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_8_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_8_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_8_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_8_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_8_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_8_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_8_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_8_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_8_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_8_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_8_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_8_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_8_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_8_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_8_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_8_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_8_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_8_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_8_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_8_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_8_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_8_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_8_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_8_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_8_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_8_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_8_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_8_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_8_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_8_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_8_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_8_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_8_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_8_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_8_io_brupdate_b2_target_offset),
    .io_kill(slots_8_io_kill),
    .io_clear(slots_8_io_clear),
    .io_ldspec_miss(slots_8_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_8_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_8_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_8_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_1_valid(slots_8_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_8_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_8_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_2_valid(slots_8_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_8_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_8_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_3_valid(slots_8_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_8_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_8_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_4_valid(slots_8_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_8_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_8_io_wakeup_ports_4_bits_poisoned),
    .io_pred_wakeup_port_valid(slots_8_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_8_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_8_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_8_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_8_io_in_uop_valid),
    .io_in_uop_bits_uopc(slots_8_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_8_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_8_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_8_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_8_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_8_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_8_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_8_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_8_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_8_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_8_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_8_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_8_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_8_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_8_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_8_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_8_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_iw_state(slots_8_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_8_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_8_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_8_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_8_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_8_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_8_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_8_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_8_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_8_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_8_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_8_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_8_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_8_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_8_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_8_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_8_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_8_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_8_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_8_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_8_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_8_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_8_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_8_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_8_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_8_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_8_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_8_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_8_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_8_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_8_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_8_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_8_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_8_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_8_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_8_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_8_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_8_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_8_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_8_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_8_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_8_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_8_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_8_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_8_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_8_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_8_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_8_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_8_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_8_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_8_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_8_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_8_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_8_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_8_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_8_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_8_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_8_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_8_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_8_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_8_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_8_io_in_uop_bits_debug_tsrc),
    .io_out_uop_uopc(slots_8_io_out_uop_uopc),
    .io_out_uop_inst(slots_8_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_8_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_8_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_8_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_8_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_8_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_8_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_8_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_8_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_8_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_8_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_8_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_8_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_8_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_8_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_8_io_out_uop_ctrl_is_std),
    .io_out_uop_iw_state(slots_8_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_8_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_8_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_8_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_8_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_8_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_8_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_8_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_8_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_8_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_8_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_8_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_8_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_8_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_8_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_8_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_8_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_8_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_8_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_8_io_out_uop_pdst),
    .io_out_uop_prs1(slots_8_io_out_uop_prs1),
    .io_out_uop_prs2(slots_8_io_out_uop_prs2),
    .io_out_uop_prs3(slots_8_io_out_uop_prs3),
    .io_out_uop_ppred(slots_8_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_8_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_8_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_8_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_8_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_8_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_8_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_8_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_8_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_8_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_8_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_8_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_8_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_8_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_8_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_8_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_8_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_8_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_8_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_8_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_8_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_8_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_8_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_8_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_8_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_8_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_8_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_8_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_8_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_8_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_8_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_8_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_8_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_8_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_8_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_8_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_8_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_8_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_8_io_out_uop_debug_tsrc),
    .io_uop_uopc(slots_8_io_uop_uopc),
    .io_uop_inst(slots_8_io_uop_inst),
    .io_uop_debug_inst(slots_8_io_uop_debug_inst),
    .io_uop_is_rvc(slots_8_io_uop_is_rvc),
    .io_uop_debug_pc(slots_8_io_uop_debug_pc),
    .io_uop_iq_type(slots_8_io_uop_iq_type),
    .io_uop_fu_code(slots_8_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_8_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_8_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_8_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_8_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_8_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_8_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_8_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_8_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_8_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_8_io_uop_ctrl_is_std),
    .io_uop_iw_state(slots_8_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_8_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_8_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_8_io_uop_is_br),
    .io_uop_is_jalr(slots_8_io_uop_is_jalr),
    .io_uop_is_jal(slots_8_io_uop_is_jal),
    .io_uop_is_sfb(slots_8_io_uop_is_sfb),
    .io_uop_br_mask(slots_8_io_uop_br_mask),
    .io_uop_br_tag(slots_8_io_uop_br_tag),
    .io_uop_ftq_idx(slots_8_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_8_io_uop_edge_inst),
    .io_uop_pc_lob(slots_8_io_uop_pc_lob),
    .io_uop_taken(slots_8_io_uop_taken),
    .io_uop_imm_packed(slots_8_io_uop_imm_packed),
    .io_uop_csr_addr(slots_8_io_uop_csr_addr),
    .io_uop_rob_idx(slots_8_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_8_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_8_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_8_io_uop_rxq_idx),
    .io_uop_pdst(slots_8_io_uop_pdst),
    .io_uop_prs1(slots_8_io_uop_prs1),
    .io_uop_prs2(slots_8_io_uop_prs2),
    .io_uop_prs3(slots_8_io_uop_prs3),
    .io_uop_ppred(slots_8_io_uop_ppred),
    .io_uop_prs1_busy(slots_8_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_8_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_8_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_8_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_8_io_uop_stale_pdst),
    .io_uop_exception(slots_8_io_uop_exception),
    .io_uop_exc_cause(slots_8_io_uop_exc_cause),
    .io_uop_bypassable(slots_8_io_uop_bypassable),
    .io_uop_mem_cmd(slots_8_io_uop_mem_cmd),
    .io_uop_mem_size(slots_8_io_uop_mem_size),
    .io_uop_mem_signed(slots_8_io_uop_mem_signed),
    .io_uop_is_fence(slots_8_io_uop_is_fence),
    .io_uop_is_fencei(slots_8_io_uop_is_fencei),
    .io_uop_is_amo(slots_8_io_uop_is_amo),
    .io_uop_uses_ldq(slots_8_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_8_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_8_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_8_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_8_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_8_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_8_io_uop_ldst),
    .io_uop_lrs1(slots_8_io_uop_lrs1),
    .io_uop_lrs2(slots_8_io_uop_lrs2),
    .io_uop_lrs3(slots_8_io_uop_lrs3),
    .io_uop_ldst_val(slots_8_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_8_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_8_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_8_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_8_io_uop_frs3_en),
    .io_uop_fp_val(slots_8_io_uop_fp_val),
    .io_uop_fp_single(slots_8_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_8_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_8_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_8_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_8_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_8_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_8_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_8_io_uop_debug_tsrc),
    .io_debug_p1(slots_8_io_debug_p1),
    .io_debug_p2(slots_8_io_debug_p2),
    .io_debug_p3(slots_8_io_debug_p3),
    .io_debug_ppred(slots_8_io_debug_ppred),
    .io_debug_state(slots_8_io_debug_state)
  );
  IssueSlot_16 slots_9 ( // @[issue-unit.scala 153:73]
    .clock(slots_9_clock),
    .reset(slots_9_reset),
    .io_valid(slots_9_io_valid),
    .io_will_be_valid(slots_9_io_will_be_valid),
    .io_request(slots_9_io_request),
    .io_request_hp(slots_9_io_request_hp),
    .io_grant(slots_9_io_grant),
    .io_brupdate_b1_resolve_mask(slots_9_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_9_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_uopc(slots_9_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_9_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_9_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_9_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_9_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_9_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_9_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_9_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_9_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_9_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_9_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_9_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_9_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_9_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_9_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_9_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_9_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_iw_state(slots_9_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_9_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_9_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_9_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_9_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_9_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_9_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_9_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_9_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_9_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_9_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_9_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_9_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_9_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_9_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_9_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_9_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_9_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_9_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_9_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_9_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_9_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_9_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_9_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_9_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_9_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_9_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_9_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_9_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_9_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_9_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_9_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_9_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_9_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_9_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_9_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_9_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_9_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_9_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_9_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_9_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_9_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_9_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_9_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_9_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_9_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_9_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_9_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_9_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_9_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_9_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_9_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_9_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_9_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_9_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_9_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_9_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_9_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_9_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_9_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_9_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_9_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_9_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_9_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_9_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_9_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_9_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_9_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_9_io_brupdate_b2_target_offset),
    .io_kill(slots_9_io_kill),
    .io_clear(slots_9_io_clear),
    .io_ldspec_miss(slots_9_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_9_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_9_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_9_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_1_valid(slots_9_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_9_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_9_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_2_valid(slots_9_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_9_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_9_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_3_valid(slots_9_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_9_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_9_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_4_valid(slots_9_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_9_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_9_io_wakeup_ports_4_bits_poisoned),
    .io_pred_wakeup_port_valid(slots_9_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_9_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_9_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_9_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_9_io_in_uop_valid),
    .io_in_uop_bits_uopc(slots_9_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_9_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_9_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_9_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_9_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_9_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_9_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_9_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_9_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_9_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_9_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_9_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_9_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_9_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_9_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_9_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_9_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_iw_state(slots_9_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_9_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_9_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_9_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_9_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_9_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_9_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_9_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_9_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_9_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_9_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_9_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_9_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_9_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_9_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_9_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_9_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_9_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_9_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_9_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_9_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_9_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_9_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_9_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_9_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_9_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_9_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_9_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_9_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_9_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_9_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_9_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_9_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_9_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_9_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_9_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_9_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_9_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_9_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_9_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_9_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_9_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_9_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_9_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_9_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_9_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_9_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_9_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_9_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_9_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_9_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_9_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_9_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_9_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_9_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_9_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_9_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_9_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_9_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_9_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_9_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_9_io_in_uop_bits_debug_tsrc),
    .io_out_uop_uopc(slots_9_io_out_uop_uopc),
    .io_out_uop_inst(slots_9_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_9_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_9_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_9_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_9_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_9_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_9_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_9_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_9_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_9_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_9_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_9_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_9_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_9_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_9_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_9_io_out_uop_ctrl_is_std),
    .io_out_uop_iw_state(slots_9_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_9_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_9_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_9_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_9_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_9_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_9_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_9_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_9_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_9_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_9_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_9_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_9_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_9_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_9_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_9_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_9_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_9_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_9_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_9_io_out_uop_pdst),
    .io_out_uop_prs1(slots_9_io_out_uop_prs1),
    .io_out_uop_prs2(slots_9_io_out_uop_prs2),
    .io_out_uop_prs3(slots_9_io_out_uop_prs3),
    .io_out_uop_ppred(slots_9_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_9_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_9_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_9_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_9_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_9_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_9_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_9_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_9_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_9_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_9_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_9_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_9_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_9_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_9_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_9_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_9_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_9_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_9_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_9_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_9_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_9_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_9_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_9_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_9_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_9_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_9_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_9_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_9_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_9_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_9_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_9_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_9_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_9_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_9_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_9_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_9_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_9_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_9_io_out_uop_debug_tsrc),
    .io_uop_uopc(slots_9_io_uop_uopc),
    .io_uop_inst(slots_9_io_uop_inst),
    .io_uop_debug_inst(slots_9_io_uop_debug_inst),
    .io_uop_is_rvc(slots_9_io_uop_is_rvc),
    .io_uop_debug_pc(slots_9_io_uop_debug_pc),
    .io_uop_iq_type(slots_9_io_uop_iq_type),
    .io_uop_fu_code(slots_9_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_9_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_9_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_9_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_9_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_9_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_9_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_9_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_9_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_9_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_9_io_uop_ctrl_is_std),
    .io_uop_iw_state(slots_9_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_9_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_9_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_9_io_uop_is_br),
    .io_uop_is_jalr(slots_9_io_uop_is_jalr),
    .io_uop_is_jal(slots_9_io_uop_is_jal),
    .io_uop_is_sfb(slots_9_io_uop_is_sfb),
    .io_uop_br_mask(slots_9_io_uop_br_mask),
    .io_uop_br_tag(slots_9_io_uop_br_tag),
    .io_uop_ftq_idx(slots_9_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_9_io_uop_edge_inst),
    .io_uop_pc_lob(slots_9_io_uop_pc_lob),
    .io_uop_taken(slots_9_io_uop_taken),
    .io_uop_imm_packed(slots_9_io_uop_imm_packed),
    .io_uop_csr_addr(slots_9_io_uop_csr_addr),
    .io_uop_rob_idx(slots_9_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_9_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_9_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_9_io_uop_rxq_idx),
    .io_uop_pdst(slots_9_io_uop_pdst),
    .io_uop_prs1(slots_9_io_uop_prs1),
    .io_uop_prs2(slots_9_io_uop_prs2),
    .io_uop_prs3(slots_9_io_uop_prs3),
    .io_uop_ppred(slots_9_io_uop_ppred),
    .io_uop_prs1_busy(slots_9_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_9_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_9_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_9_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_9_io_uop_stale_pdst),
    .io_uop_exception(slots_9_io_uop_exception),
    .io_uop_exc_cause(slots_9_io_uop_exc_cause),
    .io_uop_bypassable(slots_9_io_uop_bypassable),
    .io_uop_mem_cmd(slots_9_io_uop_mem_cmd),
    .io_uop_mem_size(slots_9_io_uop_mem_size),
    .io_uop_mem_signed(slots_9_io_uop_mem_signed),
    .io_uop_is_fence(slots_9_io_uop_is_fence),
    .io_uop_is_fencei(slots_9_io_uop_is_fencei),
    .io_uop_is_amo(slots_9_io_uop_is_amo),
    .io_uop_uses_ldq(slots_9_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_9_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_9_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_9_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_9_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_9_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_9_io_uop_ldst),
    .io_uop_lrs1(slots_9_io_uop_lrs1),
    .io_uop_lrs2(slots_9_io_uop_lrs2),
    .io_uop_lrs3(slots_9_io_uop_lrs3),
    .io_uop_ldst_val(slots_9_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_9_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_9_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_9_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_9_io_uop_frs3_en),
    .io_uop_fp_val(slots_9_io_uop_fp_val),
    .io_uop_fp_single(slots_9_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_9_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_9_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_9_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_9_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_9_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_9_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_9_io_uop_debug_tsrc),
    .io_debug_p1(slots_9_io_debug_p1),
    .io_debug_p2(slots_9_io_debug_p2),
    .io_debug_p3(slots_9_io_debug_p3),
    .io_debug_ppred(slots_9_io_debug_ppred),
    .io_debug_state(slots_9_io_debug_state)
  );
  IssueSlot_16 slots_10 ( // @[issue-unit.scala 153:73]
    .clock(slots_10_clock),
    .reset(slots_10_reset),
    .io_valid(slots_10_io_valid),
    .io_will_be_valid(slots_10_io_will_be_valid),
    .io_request(slots_10_io_request),
    .io_request_hp(slots_10_io_request_hp),
    .io_grant(slots_10_io_grant),
    .io_brupdate_b1_resolve_mask(slots_10_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_10_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_uopc(slots_10_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_10_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_10_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_10_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_10_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_10_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_10_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_10_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_10_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_10_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_10_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_10_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_10_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_10_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_10_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_10_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_10_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_iw_state(slots_10_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_10_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_10_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_10_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_10_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_10_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_10_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_10_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_10_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_10_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_10_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_10_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_10_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_10_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_10_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_10_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_10_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_10_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_10_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_10_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_10_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_10_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_10_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_10_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_10_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_10_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_10_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_10_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_10_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_10_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_10_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_10_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_10_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_10_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_10_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_10_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_10_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_10_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_10_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_10_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_10_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_10_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_10_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_10_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_10_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_10_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_10_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_10_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_10_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_10_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_10_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_10_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_10_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_10_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_10_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_10_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_10_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_10_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_10_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_10_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_10_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_10_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_10_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_10_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_10_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_10_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_10_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_10_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_10_io_brupdate_b2_target_offset),
    .io_kill(slots_10_io_kill),
    .io_clear(slots_10_io_clear),
    .io_ldspec_miss(slots_10_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_10_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_10_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_10_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_1_valid(slots_10_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_10_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_10_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_2_valid(slots_10_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_10_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_10_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_3_valid(slots_10_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_10_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_10_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_4_valid(slots_10_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_10_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_10_io_wakeup_ports_4_bits_poisoned),
    .io_pred_wakeup_port_valid(slots_10_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_10_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_10_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_10_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_10_io_in_uop_valid),
    .io_in_uop_bits_uopc(slots_10_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_10_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_10_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_10_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_10_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_10_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_10_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_10_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_10_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_10_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_10_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_10_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_10_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_10_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_10_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_10_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_10_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_iw_state(slots_10_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_10_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_10_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_10_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_10_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_10_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_10_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_10_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_10_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_10_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_10_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_10_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_10_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_10_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_10_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_10_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_10_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_10_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_10_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_10_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_10_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_10_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_10_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_10_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_10_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_10_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_10_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_10_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_10_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_10_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_10_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_10_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_10_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_10_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_10_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_10_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_10_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_10_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_10_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_10_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_10_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_10_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_10_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_10_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_10_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_10_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_10_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_10_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_10_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_10_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_10_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_10_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_10_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_10_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_10_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_10_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_10_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_10_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_10_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_10_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_10_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_10_io_in_uop_bits_debug_tsrc),
    .io_out_uop_uopc(slots_10_io_out_uop_uopc),
    .io_out_uop_inst(slots_10_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_10_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_10_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_10_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_10_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_10_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_10_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_10_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_10_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_10_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_10_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_10_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_10_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_10_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_10_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_10_io_out_uop_ctrl_is_std),
    .io_out_uop_iw_state(slots_10_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_10_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_10_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_10_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_10_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_10_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_10_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_10_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_10_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_10_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_10_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_10_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_10_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_10_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_10_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_10_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_10_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_10_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_10_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_10_io_out_uop_pdst),
    .io_out_uop_prs1(slots_10_io_out_uop_prs1),
    .io_out_uop_prs2(slots_10_io_out_uop_prs2),
    .io_out_uop_prs3(slots_10_io_out_uop_prs3),
    .io_out_uop_ppred(slots_10_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_10_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_10_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_10_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_10_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_10_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_10_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_10_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_10_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_10_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_10_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_10_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_10_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_10_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_10_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_10_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_10_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_10_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_10_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_10_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_10_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_10_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_10_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_10_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_10_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_10_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_10_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_10_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_10_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_10_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_10_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_10_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_10_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_10_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_10_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_10_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_10_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_10_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_10_io_out_uop_debug_tsrc),
    .io_uop_uopc(slots_10_io_uop_uopc),
    .io_uop_inst(slots_10_io_uop_inst),
    .io_uop_debug_inst(slots_10_io_uop_debug_inst),
    .io_uop_is_rvc(slots_10_io_uop_is_rvc),
    .io_uop_debug_pc(slots_10_io_uop_debug_pc),
    .io_uop_iq_type(slots_10_io_uop_iq_type),
    .io_uop_fu_code(slots_10_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_10_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_10_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_10_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_10_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_10_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_10_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_10_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_10_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_10_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_10_io_uop_ctrl_is_std),
    .io_uop_iw_state(slots_10_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_10_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_10_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_10_io_uop_is_br),
    .io_uop_is_jalr(slots_10_io_uop_is_jalr),
    .io_uop_is_jal(slots_10_io_uop_is_jal),
    .io_uop_is_sfb(slots_10_io_uop_is_sfb),
    .io_uop_br_mask(slots_10_io_uop_br_mask),
    .io_uop_br_tag(slots_10_io_uop_br_tag),
    .io_uop_ftq_idx(slots_10_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_10_io_uop_edge_inst),
    .io_uop_pc_lob(slots_10_io_uop_pc_lob),
    .io_uop_taken(slots_10_io_uop_taken),
    .io_uop_imm_packed(slots_10_io_uop_imm_packed),
    .io_uop_csr_addr(slots_10_io_uop_csr_addr),
    .io_uop_rob_idx(slots_10_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_10_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_10_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_10_io_uop_rxq_idx),
    .io_uop_pdst(slots_10_io_uop_pdst),
    .io_uop_prs1(slots_10_io_uop_prs1),
    .io_uop_prs2(slots_10_io_uop_prs2),
    .io_uop_prs3(slots_10_io_uop_prs3),
    .io_uop_ppred(slots_10_io_uop_ppred),
    .io_uop_prs1_busy(slots_10_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_10_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_10_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_10_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_10_io_uop_stale_pdst),
    .io_uop_exception(slots_10_io_uop_exception),
    .io_uop_exc_cause(slots_10_io_uop_exc_cause),
    .io_uop_bypassable(slots_10_io_uop_bypassable),
    .io_uop_mem_cmd(slots_10_io_uop_mem_cmd),
    .io_uop_mem_size(slots_10_io_uop_mem_size),
    .io_uop_mem_signed(slots_10_io_uop_mem_signed),
    .io_uop_is_fence(slots_10_io_uop_is_fence),
    .io_uop_is_fencei(slots_10_io_uop_is_fencei),
    .io_uop_is_amo(slots_10_io_uop_is_amo),
    .io_uop_uses_ldq(slots_10_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_10_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_10_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_10_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_10_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_10_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_10_io_uop_ldst),
    .io_uop_lrs1(slots_10_io_uop_lrs1),
    .io_uop_lrs2(slots_10_io_uop_lrs2),
    .io_uop_lrs3(slots_10_io_uop_lrs3),
    .io_uop_ldst_val(slots_10_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_10_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_10_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_10_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_10_io_uop_frs3_en),
    .io_uop_fp_val(slots_10_io_uop_fp_val),
    .io_uop_fp_single(slots_10_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_10_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_10_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_10_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_10_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_10_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_10_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_10_io_uop_debug_tsrc),
    .io_debug_p1(slots_10_io_debug_p1),
    .io_debug_p2(slots_10_io_debug_p2),
    .io_debug_p3(slots_10_io_debug_p3),
    .io_debug_ppred(slots_10_io_debug_ppred),
    .io_debug_state(slots_10_io_debug_state)
  );
  IssueSlot_16 slots_11 ( // @[issue-unit.scala 153:73]
    .clock(slots_11_clock),
    .reset(slots_11_reset),
    .io_valid(slots_11_io_valid),
    .io_will_be_valid(slots_11_io_will_be_valid),
    .io_request(slots_11_io_request),
    .io_request_hp(slots_11_io_request_hp),
    .io_grant(slots_11_io_grant),
    .io_brupdate_b1_resolve_mask(slots_11_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_11_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_uopc(slots_11_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_11_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_11_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_11_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_11_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_11_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_11_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_11_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_11_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_11_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_11_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_11_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_11_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_11_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_11_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_11_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_11_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_iw_state(slots_11_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_11_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_11_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_11_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_11_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_11_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_11_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_11_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_11_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_11_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_11_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_11_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_11_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_11_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_11_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_11_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_11_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_11_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_11_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_11_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_11_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_11_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_11_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_11_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_11_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_11_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_11_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_11_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_11_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_11_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_11_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_11_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_11_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_11_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_11_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_11_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_11_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_11_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_11_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_11_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_11_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_11_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_11_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_11_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_11_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_11_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_11_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_11_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_11_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_11_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_11_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_11_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_11_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_11_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_11_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_11_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_11_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_11_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_11_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_11_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_11_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_11_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_11_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_11_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_11_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_11_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_11_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_11_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_11_io_brupdate_b2_target_offset),
    .io_kill(slots_11_io_kill),
    .io_clear(slots_11_io_clear),
    .io_ldspec_miss(slots_11_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_11_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_11_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_11_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_1_valid(slots_11_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_11_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_11_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_2_valid(slots_11_io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst(slots_11_io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_2_bits_poisoned(slots_11_io_wakeup_ports_2_bits_poisoned),
    .io_wakeup_ports_3_valid(slots_11_io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst(slots_11_io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_3_bits_poisoned(slots_11_io_wakeup_ports_3_bits_poisoned),
    .io_wakeup_ports_4_valid(slots_11_io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst(slots_11_io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_4_bits_poisoned(slots_11_io_wakeup_ports_4_bits_poisoned),
    .io_pred_wakeup_port_valid(slots_11_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_11_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_11_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_11_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_11_io_in_uop_valid),
    .io_in_uop_bits_uopc(slots_11_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_11_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_11_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_11_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_11_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_11_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_11_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_11_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_11_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_11_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_11_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_11_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_11_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_11_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_11_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_11_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_11_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_iw_state(slots_11_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_11_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_11_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_11_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_11_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_11_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_11_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_11_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_11_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_11_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_11_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_11_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_11_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_11_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_11_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_11_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_11_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_11_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_11_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_11_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_11_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_11_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_11_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_11_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_11_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_11_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_11_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_11_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_11_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_11_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_11_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_11_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_11_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_11_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_11_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_11_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_11_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_11_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_11_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_11_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_11_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_11_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_11_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_11_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_11_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_11_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_11_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_11_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_11_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_11_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_11_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_11_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_11_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_11_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_11_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_11_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_11_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_11_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_11_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_11_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_11_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_11_io_in_uop_bits_debug_tsrc),
    .io_out_uop_uopc(slots_11_io_out_uop_uopc),
    .io_out_uop_inst(slots_11_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_11_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_11_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_11_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_11_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_11_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_11_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_11_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_11_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_11_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_11_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_11_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_11_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_11_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_11_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_11_io_out_uop_ctrl_is_std),
    .io_out_uop_iw_state(slots_11_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_11_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_11_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_11_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_11_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_11_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_11_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_11_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_11_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_11_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_11_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_11_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_11_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_11_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_11_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_11_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_11_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_11_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_11_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_11_io_out_uop_pdst),
    .io_out_uop_prs1(slots_11_io_out_uop_prs1),
    .io_out_uop_prs2(slots_11_io_out_uop_prs2),
    .io_out_uop_prs3(slots_11_io_out_uop_prs3),
    .io_out_uop_ppred(slots_11_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_11_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_11_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_11_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_11_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_11_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_11_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_11_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_11_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_11_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_11_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_11_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_11_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_11_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_11_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_11_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_11_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_11_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_11_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_11_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_11_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_11_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_11_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_11_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_11_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_11_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_11_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_11_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_11_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_11_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_11_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_11_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_11_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_11_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_11_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_11_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_11_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_11_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_11_io_out_uop_debug_tsrc),
    .io_uop_uopc(slots_11_io_uop_uopc),
    .io_uop_inst(slots_11_io_uop_inst),
    .io_uop_debug_inst(slots_11_io_uop_debug_inst),
    .io_uop_is_rvc(slots_11_io_uop_is_rvc),
    .io_uop_debug_pc(slots_11_io_uop_debug_pc),
    .io_uop_iq_type(slots_11_io_uop_iq_type),
    .io_uop_fu_code(slots_11_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_11_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_11_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_11_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_11_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_11_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_11_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_11_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_11_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_11_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_11_io_uop_ctrl_is_std),
    .io_uop_iw_state(slots_11_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_11_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_11_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_11_io_uop_is_br),
    .io_uop_is_jalr(slots_11_io_uop_is_jalr),
    .io_uop_is_jal(slots_11_io_uop_is_jal),
    .io_uop_is_sfb(slots_11_io_uop_is_sfb),
    .io_uop_br_mask(slots_11_io_uop_br_mask),
    .io_uop_br_tag(slots_11_io_uop_br_tag),
    .io_uop_ftq_idx(slots_11_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_11_io_uop_edge_inst),
    .io_uop_pc_lob(slots_11_io_uop_pc_lob),
    .io_uop_taken(slots_11_io_uop_taken),
    .io_uop_imm_packed(slots_11_io_uop_imm_packed),
    .io_uop_csr_addr(slots_11_io_uop_csr_addr),
    .io_uop_rob_idx(slots_11_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_11_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_11_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_11_io_uop_rxq_idx),
    .io_uop_pdst(slots_11_io_uop_pdst),
    .io_uop_prs1(slots_11_io_uop_prs1),
    .io_uop_prs2(slots_11_io_uop_prs2),
    .io_uop_prs3(slots_11_io_uop_prs3),
    .io_uop_ppred(slots_11_io_uop_ppred),
    .io_uop_prs1_busy(slots_11_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_11_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_11_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_11_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_11_io_uop_stale_pdst),
    .io_uop_exception(slots_11_io_uop_exception),
    .io_uop_exc_cause(slots_11_io_uop_exc_cause),
    .io_uop_bypassable(slots_11_io_uop_bypassable),
    .io_uop_mem_cmd(slots_11_io_uop_mem_cmd),
    .io_uop_mem_size(slots_11_io_uop_mem_size),
    .io_uop_mem_signed(slots_11_io_uop_mem_signed),
    .io_uop_is_fence(slots_11_io_uop_is_fence),
    .io_uop_is_fencei(slots_11_io_uop_is_fencei),
    .io_uop_is_amo(slots_11_io_uop_is_amo),
    .io_uop_uses_ldq(slots_11_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_11_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_11_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_11_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_11_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_11_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_11_io_uop_ldst),
    .io_uop_lrs1(slots_11_io_uop_lrs1),
    .io_uop_lrs2(slots_11_io_uop_lrs2),
    .io_uop_lrs3(slots_11_io_uop_lrs3),
    .io_uop_ldst_val(slots_11_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_11_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_11_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_11_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_11_io_uop_frs3_en),
    .io_uop_fp_val(slots_11_io_uop_fp_val),
    .io_uop_fp_single(slots_11_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_11_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_11_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_11_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_11_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_11_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_11_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_11_io_uop_debug_tsrc),
    .io_debug_p1(slots_11_io_debug_p1),
    .io_debug_p2(slots_11_io_debug_p2),
    .io_debug_p3(slots_11_io_debug_p3),
    .io_debug_ppred(slots_11_io_debug_ppred),
    .io_debug_state(slots_11_io_debug_state)
  );
  assign io_dis_uops_0_ready = REG; // @[issue-unit-age-ordered.scala 87:26]
  assign io_dis_uops_1_ready = REG_1; // @[issue-unit-age-ordered.scala 87:26]
  assign io_iss_valids_0 = issue_slots_11_grant | (issue_slots_10_grant | (issue_slots_9_grant | (issue_slots_8_grant |
    (issue_slots_7_grant | (issue_slots_6_grant | (issue_slots_5_grant | (issue_slots_4_grant | (issue_slots_3_grant | (
    issue_slots_2_grant | (issue_slots_1_grant | _T_279)))))))))); // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 120:26]
  assign io_iss_uops_0_uopc = issue_slots_11_grant ? issue_slots_11_uop_uopc : _GEN_2845; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_inst = issue_slots_11_grant ? issue_slots_11_uop_inst : _GEN_2844; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_debug_inst = issue_slots_11_grant ? issue_slots_11_uop_debug_inst : _GEN_2843; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_is_rvc = issue_slots_11_grant ? issue_slots_11_uop_is_rvc : _GEN_2842; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_debug_pc = issue_slots_11_grant ? issue_slots_11_uop_debug_pc : _GEN_2841; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_iq_type = issue_slots_11_grant ? issue_slots_11_uop_iq_type : _GEN_2840; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_fu_code = issue_slots_11_grant ? issue_slots_11_uop_fu_code : _GEN_2839; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_ctrl_br_type = issue_slots_11_grant ? issue_slots_11_uop_ctrl_br_type : _GEN_2838; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_ctrl_op1_sel = issue_slots_11_grant ? issue_slots_11_uop_ctrl_op1_sel : _GEN_2837; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_ctrl_op2_sel = issue_slots_11_grant ? issue_slots_11_uop_ctrl_op2_sel : _GEN_2836; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_ctrl_imm_sel = issue_slots_11_grant ? issue_slots_11_uop_ctrl_imm_sel : _GEN_2835; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_ctrl_op_fcn = issue_slots_11_grant ? issue_slots_11_uop_ctrl_op_fcn : _GEN_2834; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_ctrl_fcn_dw = issue_slots_11_grant ? issue_slots_11_uop_ctrl_fcn_dw : _GEN_2833; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_ctrl_csr_cmd = issue_slots_11_grant ? issue_slots_11_uop_ctrl_csr_cmd : _GEN_2832; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_ctrl_is_load = issue_slots_11_grant ? issue_slots_11_uop_ctrl_is_load : _GEN_2831; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_ctrl_is_sta = issue_slots_11_grant ? issue_slots_11_uop_ctrl_is_sta : _GEN_2830; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_ctrl_is_std = issue_slots_11_grant ? issue_slots_11_uop_ctrl_is_std : _GEN_2829; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_iw_state = issue_slots_11_grant ? issue_slots_11_uop_iw_state : _GEN_2828; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_iw_p1_poisoned = issue_slots_11_grant ? issue_slots_11_uop_iw_p1_poisoned : _GEN_2827; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_iw_p2_poisoned = issue_slots_11_grant ? issue_slots_11_uop_iw_p2_poisoned : _GEN_2826; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_is_br = issue_slots_11_grant ? issue_slots_11_uop_is_br : _GEN_2825; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_is_jalr = issue_slots_11_grant ? issue_slots_11_uop_is_jalr : _GEN_2824; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_is_jal = issue_slots_11_grant ? issue_slots_11_uop_is_jal : _GEN_2823; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_is_sfb = issue_slots_11_grant ? issue_slots_11_uop_is_sfb : _GEN_2822; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_br_mask = issue_slots_11_grant ? issue_slots_11_uop_br_mask : _GEN_2821; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_br_tag = issue_slots_11_grant ? issue_slots_11_uop_br_tag : _GEN_2820; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_ftq_idx = issue_slots_11_grant ? issue_slots_11_uop_ftq_idx : _GEN_2819; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_edge_inst = issue_slots_11_grant ? issue_slots_11_uop_edge_inst : _GEN_2818; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_pc_lob = issue_slots_11_grant ? issue_slots_11_uop_pc_lob : _GEN_2817; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_taken = issue_slots_11_grant ? issue_slots_11_uop_taken : _GEN_2816; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_imm_packed = issue_slots_11_grant ? issue_slots_11_uop_imm_packed : _GEN_2815; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_csr_addr = issue_slots_11_grant ? issue_slots_11_uop_csr_addr : _GEN_2814; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_rob_idx = issue_slots_11_grant ? issue_slots_11_uop_rob_idx : _GEN_2813; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_ldq_idx = issue_slots_11_grant ? issue_slots_11_uop_ldq_idx : _GEN_2812; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_stq_idx = issue_slots_11_grant ? issue_slots_11_uop_stq_idx : _GEN_2811; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_rxq_idx = issue_slots_11_grant ? issue_slots_11_uop_rxq_idx : _GEN_2810; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_pdst = issue_slots_11_grant ? issue_slots_11_uop_pdst : _GEN_2809; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_prs1 = issue_slots_11_grant ? issue_slots_11_uop_prs1 : _GEN_2808; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_prs2 = issue_slots_11_grant ? issue_slots_11_uop_prs2 : _GEN_2807; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_prs3 = issue_slots_11_grant ? issue_slots_11_uop_prs3 : _GEN_2806; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_ppred = issue_slots_11_grant ? issue_slots_11_uop_ppred : _GEN_2805; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_prs1_busy = issue_slots_11_grant ? issue_slots_11_uop_prs1_busy : _GEN_2804; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_prs2_busy = issue_slots_11_grant ? issue_slots_11_uop_prs2_busy : _GEN_2803; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_prs3_busy = issue_slots_11_grant ? issue_slots_11_uop_prs3_busy : _GEN_2802; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_ppred_busy = issue_slots_11_grant ? issue_slots_11_uop_ppred_busy : _GEN_2801; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_stale_pdst = issue_slots_11_grant ? issue_slots_11_uop_stale_pdst : _GEN_2800; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_exception = issue_slots_11_grant ? issue_slots_11_uop_exception : _GEN_2799; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_exc_cause = issue_slots_11_grant ? issue_slots_11_uop_exc_cause : _GEN_2798; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_bypassable = issue_slots_11_grant ? issue_slots_11_uop_bypassable : _GEN_2797; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_mem_cmd = issue_slots_11_grant ? issue_slots_11_uop_mem_cmd : _GEN_2796; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_mem_size = issue_slots_11_grant ? issue_slots_11_uop_mem_size : _GEN_2795; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_mem_signed = issue_slots_11_grant ? issue_slots_11_uop_mem_signed : _GEN_2794; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_is_fence = issue_slots_11_grant ? issue_slots_11_uop_is_fence : _GEN_2793; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_is_fencei = issue_slots_11_grant ? issue_slots_11_uop_is_fencei : _GEN_2792; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_is_amo = issue_slots_11_grant ? issue_slots_11_uop_is_amo : _GEN_2791; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_uses_ldq = issue_slots_11_grant ? issue_slots_11_uop_uses_ldq : _GEN_2790; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_uses_stq = issue_slots_11_grant ? issue_slots_11_uop_uses_stq : _GEN_2789; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_is_sys_pc2epc = issue_slots_11_grant ? issue_slots_11_uop_is_sys_pc2epc : _GEN_2788; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_is_unique = issue_slots_11_grant ? issue_slots_11_uop_is_unique : _GEN_2787; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_flush_on_commit = issue_slots_11_grant ? issue_slots_11_uop_flush_on_commit : _GEN_2786; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_ldst_is_rs1 = issue_slots_11_grant ? issue_slots_11_uop_ldst_is_rs1 : _GEN_2785; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_ldst = issue_slots_11_grant ? issue_slots_11_uop_ldst : _GEN_2784; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_lrs1 = issue_slots_11_grant ? issue_slots_11_uop_lrs1 : _GEN_2783; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_lrs2 = issue_slots_11_grant ? issue_slots_11_uop_lrs2 : _GEN_2782; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_lrs3 = issue_slots_11_grant ? issue_slots_11_uop_lrs3 : _GEN_2781; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_ldst_val = issue_slots_11_grant ? issue_slots_11_uop_ldst_val : _GEN_2780; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_dst_rtype = issue_slots_11_grant ? issue_slots_11_uop_dst_rtype : _GEN_2779; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_lrs1_rtype = issue_slots_11_grant ? issue_slots_11_uop_lrs1_rtype : _GEN_2778; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_lrs2_rtype = issue_slots_11_grant ? issue_slots_11_uop_lrs2_rtype : _GEN_2777; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_frs3_en = issue_slots_11_grant ? issue_slots_11_uop_frs3_en : _GEN_2776; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_fp_val = issue_slots_11_grant ? issue_slots_11_uop_fp_val : _GEN_2775; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_fp_single = issue_slots_11_grant ? issue_slots_11_uop_fp_single : _GEN_2774; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_xcpt_pf_if = issue_slots_11_grant ? issue_slots_11_uop_xcpt_pf_if : _GEN_2773; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_xcpt_ae_if = issue_slots_11_grant ? issue_slots_11_uop_xcpt_ae_if : _GEN_2772; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_xcpt_ma_if = issue_slots_11_grant ? issue_slots_11_uop_xcpt_ma_if : _GEN_2771; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_bp_debug_if = issue_slots_11_grant ? issue_slots_11_uop_bp_debug_if : _GEN_2770; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_bp_xcpt_if = issue_slots_11_grant ? issue_slots_11_uop_bp_xcpt_if : _GEN_2769; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_debug_fsrc = issue_slots_11_grant ? issue_slots_11_uop_debug_fsrc : _GEN_2768; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_iss_uops_0_debug_tsrc = issue_slots_11_grant ? issue_slots_11_uop_debug_tsrc : _GEN_2767; // @[issue-unit-age-ordered.scala 118:76 issue-unit-age-ordered.scala 121:24]
  assign io_event_empty = ~(issue_slots_0_valid | issue_slots_1_valid | issue_slots_2_valid | issue_slots_3_valid |
    issue_slots_4_valid | issue_slots_5_valid | issue_slots_6_valid | issue_slots_7_valid | issue_slots_8_valid |
    issue_slots_9_valid | issue_slots_10_valid | issue_slots_11_valid); // @[issue-unit.scala 165:21]
  assign slots_0_clock = clock;
  assign slots_0_reset = reset;
  assign slots_0_io_grant = issue_slots_0_request & _T_271; // @[issue-unit-age-ordered.scala 118:40]
  assign slots_0_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_0_io_kill = io_flush_pipeline; // @[issue-unit.scala 154:28 issue-unit.scala 162:37]
  assign slots_0_io_clear = 1'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_0_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 154:28 issue-unit.scala 160:37]
  assign slots_0_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_0_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_0_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_0_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_0_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_0_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_0_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_0_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_0_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_0_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_0_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_0_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_0_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_0_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_0_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_0_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_0_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_0_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_0_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_0_io_in_uop_valid = _GEN_13[1:0] == 2'h2 ? issue_slots_2_will_be_valid : _GEN_36; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_0_io_in_uop_bits_uopc = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_uopc : issue_slots_1_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_inst = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_inst : issue_slots_1_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_debug_inst = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_debug_inst :
    issue_slots_1_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_rvc = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_is_rvc :
    issue_slots_1_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_debug_pc = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_debug_pc :
    issue_slots_1_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_iq_type = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_iq_type :
    issue_slots_1_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_fu_code = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_fu_code :
    issue_slots_1_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_br_type = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_br_type :
    issue_slots_1_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_op1_sel = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_op1_sel :
    issue_slots_1_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_op2_sel = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_op2_sel :
    issue_slots_1_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_imm_sel = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_imm_sel :
    issue_slots_1_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_op_fcn = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_op_fcn :
    issue_slots_1_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_fcn_dw = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_fcn_dw :
    issue_slots_1_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_csr_cmd = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_csr_cmd :
    issue_slots_1_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_is_load = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_is_load :
    issue_slots_1_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_is_sta = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_is_sta :
    issue_slots_1_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_is_std = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_is_std :
    issue_slots_1_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_iw_state = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_iw_state :
    issue_slots_1_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_iw_p1_poisoned = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_iw_p1_poisoned :
    issue_slots_1_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_iw_p2_poisoned = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_iw_p2_poisoned :
    issue_slots_1_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_br = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_is_br : issue_slots_1_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_jalr = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_is_jalr :
    issue_slots_1_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_jal = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_is_jal :
    issue_slots_1_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_sfb = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_is_sfb :
    issue_slots_1_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_br_mask = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_br_mask :
    issue_slots_1_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_br_tag = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_br_tag :
    issue_slots_1_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ftq_idx = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ftq_idx :
    issue_slots_1_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_edge_inst = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_edge_inst :
    issue_slots_1_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_pc_lob = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_pc_lob :
    issue_slots_1_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_taken = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_taken : issue_slots_1_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_imm_packed = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_imm_packed :
    issue_slots_1_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_csr_addr = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_csr_addr :
    issue_slots_1_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_rob_idx = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_rob_idx :
    issue_slots_1_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ldq_idx = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ldq_idx :
    issue_slots_1_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_stq_idx = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_stq_idx :
    issue_slots_1_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_rxq_idx = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_rxq_idx :
    issue_slots_1_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_pdst = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_pdst : issue_slots_1_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_prs1 = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_prs1 : issue_slots_1_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_prs2 = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_prs2 : issue_slots_1_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_prs3 = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_prs3 : issue_slots_1_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ppred = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ppred : issue_slots_1_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_prs1_busy = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_prs1_busy :
    issue_slots_1_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_prs2_busy = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_prs2_busy :
    issue_slots_1_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_prs3_busy = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_prs3_busy :
    issue_slots_1_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ppred_busy = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ppred_busy :
    issue_slots_1_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_stale_pdst = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_stale_pdst :
    issue_slots_1_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_exception = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_exception :
    issue_slots_1_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_exc_cause = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_exc_cause :
    issue_slots_1_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_bypassable = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_bypassable :
    issue_slots_1_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_mem_cmd = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_mem_cmd :
    issue_slots_1_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_mem_size = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_mem_size :
    issue_slots_1_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_mem_signed = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_mem_signed :
    issue_slots_1_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_fence = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_is_fence :
    issue_slots_1_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_fencei = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_is_fencei :
    issue_slots_1_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_amo = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_is_amo :
    issue_slots_1_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_uses_ldq = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_uses_ldq :
    issue_slots_1_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_uses_stq = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_uses_stq :
    issue_slots_1_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_sys_pc2epc = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_is_sys_pc2epc :
    issue_slots_1_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_unique = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_is_unique :
    issue_slots_1_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_flush_on_commit = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_flush_on_commit :
    issue_slots_1_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ldst_is_rs1 = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ldst_is_rs1 :
    issue_slots_1_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ldst = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ldst : issue_slots_1_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_lrs1 = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_lrs1 : issue_slots_1_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_lrs2 = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_lrs2 : issue_slots_1_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_lrs3 = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_lrs3 : issue_slots_1_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ldst_val = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_ldst_val :
    issue_slots_1_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_dst_rtype = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_dst_rtype :
    issue_slots_1_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_lrs1_rtype = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_lrs1_rtype :
    issue_slots_1_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_lrs2_rtype = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_lrs2_rtype :
    issue_slots_1_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_frs3_en = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_frs3_en :
    issue_slots_1_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_fp_val = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_fp_val :
    issue_slots_1_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_fp_single = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_fp_single :
    issue_slots_1_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_xcpt_pf_if = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_xcpt_pf_if :
    issue_slots_1_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_xcpt_ae_if = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_xcpt_ae_if :
    issue_slots_1_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_xcpt_ma_if = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_xcpt_ma_if :
    issue_slots_1_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_bp_debug_if = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_bp_debug_if :
    issue_slots_1_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_bp_xcpt_if = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_bp_xcpt_if :
    issue_slots_1_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_debug_fsrc = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_debug_fsrc :
    issue_slots_1_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_debug_tsrc = _GEN_13[1:0] == 2'h2 ? issue_slots_2_out_uop_debug_tsrc :
    issue_slots_1_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_clock = clock;
  assign slots_1_reset = reset;
  assign slots_1_io_grant = issue_slots_1_request & _T_286 & ~_T_279; // @[issue-unit-age-ordered.scala 118:56]
  assign slots_1_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_1_io_kill = io_flush_pipeline; // @[issue-unit.scala 154:28 issue-unit.scala 162:37]
  assign slots_1_io_clear = _GEN_11[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_1_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 154:28 issue-unit.scala 160:37]
  assign slots_1_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_1_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_1_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_1_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_1_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_1_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_1_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_1_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_1_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_1_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_1_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_1_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_1_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_1_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_1_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_1_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_1_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_1_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_1_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_1_io_in_uop_valid = _GEN_15[1:0] == 2'h2 ? issue_slots_3_will_be_valid : _GEN_196; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_1_io_in_uop_bits_uopc = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_uopc : issue_slots_2_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_inst = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_inst : issue_slots_2_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_debug_inst = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_debug_inst :
    issue_slots_2_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_rvc = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_is_rvc :
    issue_slots_2_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_debug_pc = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_debug_pc :
    issue_slots_2_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_iq_type = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_iq_type :
    issue_slots_2_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_fu_code = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_fu_code :
    issue_slots_2_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_br_type = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_br_type :
    issue_slots_2_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_op1_sel = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_op1_sel :
    issue_slots_2_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_op2_sel = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_op2_sel :
    issue_slots_2_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_imm_sel = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_imm_sel :
    issue_slots_2_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_op_fcn = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_op_fcn :
    issue_slots_2_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_fcn_dw = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_fcn_dw :
    issue_slots_2_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_csr_cmd = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_csr_cmd :
    issue_slots_2_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_is_load = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_is_load :
    issue_slots_2_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_is_sta = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_is_sta :
    issue_slots_2_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_is_std = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_is_std :
    issue_slots_2_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_iw_state = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_iw_state :
    issue_slots_2_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_iw_p1_poisoned = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_iw_p1_poisoned :
    issue_slots_2_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_iw_p2_poisoned = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_iw_p2_poisoned :
    issue_slots_2_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_br = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_is_br : issue_slots_2_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_jalr = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_is_jalr :
    issue_slots_2_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_jal = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_is_jal :
    issue_slots_2_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_sfb = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_is_sfb :
    issue_slots_2_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_br_mask = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_br_mask :
    issue_slots_2_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_br_tag = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_br_tag :
    issue_slots_2_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ftq_idx = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ftq_idx :
    issue_slots_2_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_edge_inst = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_edge_inst :
    issue_slots_2_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_pc_lob = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_pc_lob :
    issue_slots_2_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_taken = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_taken : issue_slots_2_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_imm_packed = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_imm_packed :
    issue_slots_2_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_csr_addr = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_csr_addr :
    issue_slots_2_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_rob_idx = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_rob_idx :
    issue_slots_2_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ldq_idx = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ldq_idx :
    issue_slots_2_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_stq_idx = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_stq_idx :
    issue_slots_2_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_rxq_idx = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_rxq_idx :
    issue_slots_2_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_pdst = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_pdst : issue_slots_2_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_prs1 = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_prs1 : issue_slots_2_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_prs2 = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_prs2 : issue_slots_2_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_prs3 = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_prs3 : issue_slots_2_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ppred = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ppred : issue_slots_2_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_prs1_busy = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_prs1_busy :
    issue_slots_2_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_prs2_busy = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_prs2_busy :
    issue_slots_2_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_prs3_busy = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_prs3_busy :
    issue_slots_2_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ppred_busy = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ppred_busy :
    issue_slots_2_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_stale_pdst = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_stale_pdst :
    issue_slots_2_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_exception = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_exception :
    issue_slots_2_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_exc_cause = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_exc_cause :
    issue_slots_2_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_bypassable = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_bypassable :
    issue_slots_2_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_mem_cmd = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_mem_cmd :
    issue_slots_2_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_mem_size = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_mem_size :
    issue_slots_2_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_mem_signed = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_mem_signed :
    issue_slots_2_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_fence = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_is_fence :
    issue_slots_2_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_fencei = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_is_fencei :
    issue_slots_2_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_amo = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_is_amo :
    issue_slots_2_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_uses_ldq = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_uses_ldq :
    issue_slots_2_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_uses_stq = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_uses_stq :
    issue_slots_2_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_sys_pc2epc = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_is_sys_pc2epc :
    issue_slots_2_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_unique = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_is_unique :
    issue_slots_2_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_flush_on_commit = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_flush_on_commit :
    issue_slots_2_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ldst_is_rs1 = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ldst_is_rs1 :
    issue_slots_2_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ldst = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ldst : issue_slots_2_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_lrs1 = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_lrs1 : issue_slots_2_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_lrs2 = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_lrs2 : issue_slots_2_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_lrs3 = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_lrs3 : issue_slots_2_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ldst_val = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_ldst_val :
    issue_slots_2_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_dst_rtype = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_dst_rtype :
    issue_slots_2_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_lrs1_rtype = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_lrs1_rtype :
    issue_slots_2_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_lrs2_rtype = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_lrs2_rtype :
    issue_slots_2_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_frs3_en = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_frs3_en :
    issue_slots_2_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_fp_val = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_fp_val :
    issue_slots_2_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_fp_single = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_fp_single :
    issue_slots_2_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_xcpt_pf_if = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_xcpt_pf_if :
    issue_slots_2_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_xcpt_ae_if = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_xcpt_ae_if :
    issue_slots_2_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_xcpt_ma_if = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_xcpt_ma_if :
    issue_slots_2_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_bp_debug_if = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_bp_debug_if :
    issue_slots_2_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_bp_xcpt_if = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_bp_xcpt_if :
    issue_slots_2_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_debug_fsrc = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_debug_fsrc :
    issue_slots_2_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_debug_tsrc = _GEN_15[1:0] == 2'h2 ? issue_slots_3_out_uop_debug_tsrc :
    issue_slots_2_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_clock = clock;
  assign slots_2_reset = reset;
  assign slots_2_io_grant = issue_slots_2_request & _T_301 & ~_T_295; // @[issue-unit-age-ordered.scala 118:56]
  assign slots_2_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_2_io_kill = io_flush_pipeline; // @[issue-unit.scala 154:28 issue-unit.scala 162:37]
  assign slots_2_io_clear = _GEN_13[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_2_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 154:28 issue-unit.scala 160:37]
  assign slots_2_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_2_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_2_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_2_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_2_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_2_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_2_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_2_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_2_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_2_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_2_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_2_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_2_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_2_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_2_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_2_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_2_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_2_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_2_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_2_io_in_uop_valid = _GEN_17[1:0] == 2'h2 ? issue_slots_4_will_be_valid : _GEN_356; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_2_io_in_uop_bits_uopc = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_uopc : issue_slots_3_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_inst = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_inst : issue_slots_3_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_debug_inst = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_debug_inst :
    issue_slots_3_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_rvc = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_is_rvc :
    issue_slots_3_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_debug_pc = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_debug_pc :
    issue_slots_3_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_iq_type = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_iq_type :
    issue_slots_3_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_fu_code = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_fu_code :
    issue_slots_3_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_br_type = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_br_type :
    issue_slots_3_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_op1_sel = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_op1_sel :
    issue_slots_3_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_op2_sel = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_op2_sel :
    issue_slots_3_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_imm_sel = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_imm_sel :
    issue_slots_3_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_op_fcn = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_op_fcn :
    issue_slots_3_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_fcn_dw = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_fcn_dw :
    issue_slots_3_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_csr_cmd = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_csr_cmd :
    issue_slots_3_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_is_load = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_is_load :
    issue_slots_3_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_is_sta = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_is_sta :
    issue_slots_3_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_is_std = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_is_std :
    issue_slots_3_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_iw_state = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_iw_state :
    issue_slots_3_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_iw_p1_poisoned = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_iw_p1_poisoned :
    issue_slots_3_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_iw_p2_poisoned = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_iw_p2_poisoned :
    issue_slots_3_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_br = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_is_br : issue_slots_3_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_jalr = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_is_jalr :
    issue_slots_3_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_jal = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_is_jal :
    issue_slots_3_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_sfb = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_is_sfb :
    issue_slots_3_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_br_mask = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_br_mask :
    issue_slots_3_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_br_tag = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_br_tag :
    issue_slots_3_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ftq_idx = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ftq_idx :
    issue_slots_3_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_edge_inst = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_edge_inst :
    issue_slots_3_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_pc_lob = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_pc_lob :
    issue_slots_3_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_taken = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_taken : issue_slots_3_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_imm_packed = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_imm_packed :
    issue_slots_3_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_csr_addr = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_csr_addr :
    issue_slots_3_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_rob_idx = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_rob_idx :
    issue_slots_3_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ldq_idx = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ldq_idx :
    issue_slots_3_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_stq_idx = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_stq_idx :
    issue_slots_3_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_rxq_idx = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_rxq_idx :
    issue_slots_3_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_pdst = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_pdst : issue_slots_3_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_prs1 = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_prs1 : issue_slots_3_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_prs2 = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_prs2 : issue_slots_3_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_prs3 = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_prs3 : issue_slots_3_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ppred = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ppred : issue_slots_3_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_prs1_busy = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_prs1_busy :
    issue_slots_3_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_prs2_busy = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_prs2_busy :
    issue_slots_3_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_prs3_busy = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_prs3_busy :
    issue_slots_3_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ppred_busy = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ppred_busy :
    issue_slots_3_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_stale_pdst = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_stale_pdst :
    issue_slots_3_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_exception = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_exception :
    issue_slots_3_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_exc_cause = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_exc_cause :
    issue_slots_3_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_bypassable = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_bypassable :
    issue_slots_3_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_mem_cmd = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_mem_cmd :
    issue_slots_3_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_mem_size = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_mem_size :
    issue_slots_3_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_mem_signed = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_mem_signed :
    issue_slots_3_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_fence = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_is_fence :
    issue_slots_3_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_fencei = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_is_fencei :
    issue_slots_3_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_amo = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_is_amo :
    issue_slots_3_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_uses_ldq = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_uses_ldq :
    issue_slots_3_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_uses_stq = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_uses_stq :
    issue_slots_3_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_sys_pc2epc = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_is_sys_pc2epc :
    issue_slots_3_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_unique = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_is_unique :
    issue_slots_3_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_flush_on_commit = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_flush_on_commit :
    issue_slots_3_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ldst_is_rs1 = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ldst_is_rs1 :
    issue_slots_3_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ldst = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ldst : issue_slots_3_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_lrs1 = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_lrs1 : issue_slots_3_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_lrs2 = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_lrs2 : issue_slots_3_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_lrs3 = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_lrs3 : issue_slots_3_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ldst_val = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_ldst_val :
    issue_slots_3_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_dst_rtype = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_dst_rtype :
    issue_slots_3_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_lrs1_rtype = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_lrs1_rtype :
    issue_slots_3_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_lrs2_rtype = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_lrs2_rtype :
    issue_slots_3_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_frs3_en = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_frs3_en :
    issue_slots_3_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_fp_val = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_fp_val :
    issue_slots_3_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_fp_single = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_fp_single :
    issue_slots_3_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_xcpt_pf_if = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_xcpt_pf_if :
    issue_slots_3_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_xcpt_ae_if = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_xcpt_ae_if :
    issue_slots_3_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_xcpt_ma_if = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_xcpt_ma_if :
    issue_slots_3_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_bp_debug_if = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_bp_debug_if :
    issue_slots_3_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_bp_xcpt_if = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_bp_xcpt_if :
    issue_slots_3_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_debug_fsrc = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_debug_fsrc :
    issue_slots_3_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_debug_tsrc = _GEN_17[1:0] == 2'h2 ? issue_slots_4_out_uop_debug_tsrc :
    issue_slots_3_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_clock = clock;
  assign slots_3_reset = reset;
  assign slots_3_io_grant = _T_324 & ~_T_310; // @[issue-unit-age-ordered.scala 118:56]
  assign slots_3_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_3_io_kill = io_flush_pipeline; // @[issue-unit.scala 154:28 issue-unit.scala 162:37]
  assign slots_3_io_clear = _GEN_15[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_3_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 154:28 issue-unit.scala 160:37]
  assign slots_3_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_3_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_3_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_3_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_3_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_3_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_3_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_3_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_3_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_3_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_3_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_3_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_3_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_3_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_3_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_3_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_3_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_3_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_3_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_3_io_in_uop_valid = _GEN_19[1:0] == 2'h2 ? issue_slots_5_will_be_valid : _GEN_516; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_3_io_in_uop_bits_uopc = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_uopc : issue_slots_4_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_inst = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_inst : issue_slots_4_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_debug_inst = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_debug_inst :
    issue_slots_4_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_rvc = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_is_rvc :
    issue_slots_4_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_debug_pc = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_debug_pc :
    issue_slots_4_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_iq_type = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_iq_type :
    issue_slots_4_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_fu_code = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_fu_code :
    issue_slots_4_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_br_type = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_br_type :
    issue_slots_4_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_op1_sel = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_op1_sel :
    issue_slots_4_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_op2_sel = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_op2_sel :
    issue_slots_4_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_imm_sel = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_imm_sel :
    issue_slots_4_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_op_fcn = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_op_fcn :
    issue_slots_4_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_fcn_dw = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_fcn_dw :
    issue_slots_4_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_csr_cmd = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_csr_cmd :
    issue_slots_4_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_is_load = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_is_load :
    issue_slots_4_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_is_sta = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_is_sta :
    issue_slots_4_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_is_std = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_is_std :
    issue_slots_4_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_iw_state = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_iw_state :
    issue_slots_4_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_iw_p1_poisoned = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_iw_p1_poisoned :
    issue_slots_4_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_iw_p2_poisoned = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_iw_p2_poisoned :
    issue_slots_4_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_br = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_is_br : issue_slots_4_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_jalr = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_is_jalr :
    issue_slots_4_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_jal = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_is_jal :
    issue_slots_4_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_sfb = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_is_sfb :
    issue_slots_4_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_br_mask = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_br_mask :
    issue_slots_4_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_br_tag = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_br_tag :
    issue_slots_4_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ftq_idx = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ftq_idx :
    issue_slots_4_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_edge_inst = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_edge_inst :
    issue_slots_4_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_pc_lob = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_pc_lob :
    issue_slots_4_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_taken = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_taken : issue_slots_4_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_imm_packed = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_imm_packed :
    issue_slots_4_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_csr_addr = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_csr_addr :
    issue_slots_4_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_rob_idx = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_rob_idx :
    issue_slots_4_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ldq_idx = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ldq_idx :
    issue_slots_4_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_stq_idx = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_stq_idx :
    issue_slots_4_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_rxq_idx = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_rxq_idx :
    issue_slots_4_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_pdst = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_pdst : issue_slots_4_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_prs1 = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_prs1 : issue_slots_4_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_prs2 = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_prs2 : issue_slots_4_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_prs3 = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_prs3 : issue_slots_4_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ppred = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ppred : issue_slots_4_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_prs1_busy = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_prs1_busy :
    issue_slots_4_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_prs2_busy = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_prs2_busy :
    issue_slots_4_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_prs3_busy = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_prs3_busy :
    issue_slots_4_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ppred_busy = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ppred_busy :
    issue_slots_4_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_stale_pdst = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_stale_pdst :
    issue_slots_4_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_exception = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_exception :
    issue_slots_4_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_exc_cause = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_exc_cause :
    issue_slots_4_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_bypassable = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_bypassable :
    issue_slots_4_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_mem_cmd = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_mem_cmd :
    issue_slots_4_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_mem_size = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_mem_size :
    issue_slots_4_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_mem_signed = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_mem_signed :
    issue_slots_4_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_fence = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_is_fence :
    issue_slots_4_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_fencei = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_is_fencei :
    issue_slots_4_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_amo = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_is_amo :
    issue_slots_4_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_uses_ldq = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_uses_ldq :
    issue_slots_4_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_uses_stq = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_uses_stq :
    issue_slots_4_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_sys_pc2epc = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_is_sys_pc2epc :
    issue_slots_4_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_unique = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_is_unique :
    issue_slots_4_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_flush_on_commit = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_flush_on_commit :
    issue_slots_4_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ldst_is_rs1 = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ldst_is_rs1 :
    issue_slots_4_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ldst = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ldst : issue_slots_4_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_lrs1 = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_lrs1 : issue_slots_4_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_lrs2 = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_lrs2 : issue_slots_4_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_lrs3 = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_lrs3 : issue_slots_4_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ldst_val = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_ldst_val :
    issue_slots_4_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_dst_rtype = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_dst_rtype :
    issue_slots_4_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_lrs1_rtype = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_lrs1_rtype :
    issue_slots_4_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_lrs2_rtype = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_lrs2_rtype :
    issue_slots_4_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_frs3_en = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_frs3_en :
    issue_slots_4_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_fp_val = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_fp_val :
    issue_slots_4_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_fp_single = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_fp_single :
    issue_slots_4_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_xcpt_pf_if = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_xcpt_pf_if :
    issue_slots_4_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_xcpt_ae_if = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_xcpt_ae_if :
    issue_slots_4_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_xcpt_ma_if = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_xcpt_ma_if :
    issue_slots_4_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_bp_debug_if = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_bp_debug_if :
    issue_slots_4_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_bp_xcpt_if = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_bp_xcpt_if :
    issue_slots_4_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_debug_fsrc = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_debug_fsrc :
    issue_slots_4_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_debug_tsrc = _GEN_19[1:0] == 2'h2 ? issue_slots_5_out_uop_debug_tsrc :
    issue_slots_4_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_clock = clock;
  assign slots_4_reset = reset;
  assign slots_4_io_grant = issue_slots_4_request & _T_331 & ~_T_325; // @[issue-unit-age-ordered.scala 118:56]
  assign slots_4_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_4_io_kill = io_flush_pipeline; // @[issue-unit.scala 154:28 issue-unit.scala 162:37]
  assign slots_4_io_clear = _GEN_17[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_4_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 154:28 issue-unit.scala 160:37]
  assign slots_4_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_4_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_4_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_4_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_4_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_4_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_4_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_4_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_4_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_4_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_4_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_4_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_4_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_4_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_4_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_4_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_4_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_4_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_4_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_4_io_in_uop_valid = _GEN_21[1:0] == 2'h2 ? issue_slots_6_will_be_valid : _GEN_676; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_4_io_in_uop_bits_uopc = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_uopc : issue_slots_5_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_inst = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_inst : issue_slots_5_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_debug_inst = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_debug_inst :
    issue_slots_5_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_rvc = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_is_rvc :
    issue_slots_5_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_debug_pc = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_debug_pc :
    issue_slots_5_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_iq_type = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_iq_type :
    issue_slots_5_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_fu_code = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_fu_code :
    issue_slots_5_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_br_type = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_br_type :
    issue_slots_5_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_op1_sel = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_op1_sel :
    issue_slots_5_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_op2_sel = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_op2_sel :
    issue_slots_5_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_imm_sel = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_imm_sel :
    issue_slots_5_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_op_fcn = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_op_fcn :
    issue_slots_5_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_fcn_dw = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_fcn_dw :
    issue_slots_5_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_csr_cmd = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_csr_cmd :
    issue_slots_5_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_is_load = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_is_load :
    issue_slots_5_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_is_sta = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_is_sta :
    issue_slots_5_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_is_std = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_is_std :
    issue_slots_5_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_iw_state = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_iw_state :
    issue_slots_5_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_iw_p1_poisoned = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_iw_p1_poisoned :
    issue_slots_5_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_iw_p2_poisoned = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_iw_p2_poisoned :
    issue_slots_5_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_br = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_is_br : issue_slots_5_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_jalr = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_is_jalr :
    issue_slots_5_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_jal = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_is_jal :
    issue_slots_5_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_sfb = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_is_sfb :
    issue_slots_5_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_br_mask = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_br_mask :
    issue_slots_5_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_br_tag = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_br_tag :
    issue_slots_5_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ftq_idx = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ftq_idx :
    issue_slots_5_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_edge_inst = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_edge_inst :
    issue_slots_5_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_pc_lob = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_pc_lob :
    issue_slots_5_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_taken = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_taken : issue_slots_5_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_imm_packed = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_imm_packed :
    issue_slots_5_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_csr_addr = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_csr_addr :
    issue_slots_5_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_rob_idx = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_rob_idx :
    issue_slots_5_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ldq_idx = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ldq_idx :
    issue_slots_5_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_stq_idx = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_stq_idx :
    issue_slots_5_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_rxq_idx = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_rxq_idx :
    issue_slots_5_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_pdst = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_pdst : issue_slots_5_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_prs1 = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_prs1 : issue_slots_5_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_prs2 = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_prs2 : issue_slots_5_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_prs3 = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_prs3 : issue_slots_5_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ppred = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ppred : issue_slots_5_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_prs1_busy = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_prs1_busy :
    issue_slots_5_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_prs2_busy = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_prs2_busy :
    issue_slots_5_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_prs3_busy = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_prs3_busy :
    issue_slots_5_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ppred_busy = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ppred_busy :
    issue_slots_5_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_stale_pdst = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_stale_pdst :
    issue_slots_5_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_exception = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_exception :
    issue_slots_5_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_exc_cause = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_exc_cause :
    issue_slots_5_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_bypassable = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_bypassable :
    issue_slots_5_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_mem_cmd = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_mem_cmd :
    issue_slots_5_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_mem_size = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_mem_size :
    issue_slots_5_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_mem_signed = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_mem_signed :
    issue_slots_5_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_fence = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_is_fence :
    issue_slots_5_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_fencei = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_is_fencei :
    issue_slots_5_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_amo = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_is_amo :
    issue_slots_5_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_uses_ldq = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_uses_ldq :
    issue_slots_5_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_uses_stq = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_uses_stq :
    issue_slots_5_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_sys_pc2epc = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_is_sys_pc2epc :
    issue_slots_5_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_unique = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_is_unique :
    issue_slots_5_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_flush_on_commit = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_flush_on_commit :
    issue_slots_5_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ldst_is_rs1 = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ldst_is_rs1 :
    issue_slots_5_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ldst = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ldst : issue_slots_5_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_lrs1 = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_lrs1 : issue_slots_5_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_lrs2 = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_lrs2 : issue_slots_5_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_lrs3 = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_lrs3 : issue_slots_5_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ldst_val = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_ldst_val :
    issue_slots_5_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_dst_rtype = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_dst_rtype :
    issue_slots_5_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_lrs1_rtype = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_lrs1_rtype :
    issue_slots_5_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_lrs2_rtype = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_lrs2_rtype :
    issue_slots_5_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_frs3_en = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_frs3_en :
    issue_slots_5_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_fp_val = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_fp_val :
    issue_slots_5_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_fp_single = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_fp_single :
    issue_slots_5_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_xcpt_pf_if = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_xcpt_pf_if :
    issue_slots_5_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_xcpt_ae_if = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_xcpt_ae_if :
    issue_slots_5_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_xcpt_ma_if = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_xcpt_ma_if :
    issue_slots_5_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_bp_debug_if = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_bp_debug_if :
    issue_slots_5_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_bp_xcpt_if = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_bp_xcpt_if :
    issue_slots_5_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_debug_fsrc = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_debug_fsrc :
    issue_slots_5_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_debug_tsrc = _GEN_21[1:0] == 2'h2 ? issue_slots_6_out_uop_debug_tsrc :
    issue_slots_5_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_clock = clock;
  assign slots_5_reset = reset;
  assign slots_5_io_grant = issue_slots_5_request & _T_346 & ~_T_340; // @[issue-unit-age-ordered.scala 118:56]
  assign slots_5_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_5_io_kill = io_flush_pipeline; // @[issue-unit.scala 154:28 issue-unit.scala 162:37]
  assign slots_5_io_clear = _GEN_19[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_5_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 154:28 issue-unit.scala 160:37]
  assign slots_5_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_5_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_5_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_5_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_5_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_5_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_5_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_5_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_5_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_5_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_5_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_5_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_5_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_5_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_5_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_5_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_5_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_5_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_5_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_5_io_in_uop_valid = _GEN_23[1:0] == 2'h2 ? issue_slots_7_will_be_valid : _GEN_836; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_5_io_in_uop_bits_uopc = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_uopc : issue_slots_6_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_inst = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_inst : issue_slots_6_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_debug_inst = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_debug_inst :
    issue_slots_6_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_rvc = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_is_rvc :
    issue_slots_6_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_debug_pc = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_debug_pc :
    issue_slots_6_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_iq_type = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_iq_type :
    issue_slots_6_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_fu_code = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_fu_code :
    issue_slots_6_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_br_type = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_br_type :
    issue_slots_6_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_op1_sel = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_op1_sel :
    issue_slots_6_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_op2_sel = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_op2_sel :
    issue_slots_6_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_imm_sel = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_imm_sel :
    issue_slots_6_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_op_fcn = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_op_fcn :
    issue_slots_6_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_fcn_dw = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_fcn_dw :
    issue_slots_6_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_csr_cmd = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_csr_cmd :
    issue_slots_6_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_is_load = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_is_load :
    issue_slots_6_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_is_sta = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_is_sta :
    issue_slots_6_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_is_std = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_is_std :
    issue_slots_6_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_iw_state = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_iw_state :
    issue_slots_6_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_iw_p1_poisoned = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_iw_p1_poisoned :
    issue_slots_6_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_iw_p2_poisoned = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_iw_p2_poisoned :
    issue_slots_6_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_br = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_is_br : issue_slots_6_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_jalr = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_is_jalr :
    issue_slots_6_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_jal = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_is_jal :
    issue_slots_6_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_sfb = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_is_sfb :
    issue_slots_6_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_br_mask = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_br_mask :
    issue_slots_6_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_br_tag = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_br_tag :
    issue_slots_6_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ftq_idx = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ftq_idx :
    issue_slots_6_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_edge_inst = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_edge_inst :
    issue_slots_6_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_pc_lob = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_pc_lob :
    issue_slots_6_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_taken = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_taken : issue_slots_6_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_imm_packed = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_imm_packed :
    issue_slots_6_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_csr_addr = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_csr_addr :
    issue_slots_6_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_rob_idx = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_rob_idx :
    issue_slots_6_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ldq_idx = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ldq_idx :
    issue_slots_6_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_stq_idx = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_stq_idx :
    issue_slots_6_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_rxq_idx = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_rxq_idx :
    issue_slots_6_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_pdst = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_pdst : issue_slots_6_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_prs1 = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_prs1 : issue_slots_6_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_prs2 = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_prs2 : issue_slots_6_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_prs3 = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_prs3 : issue_slots_6_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ppred = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ppred : issue_slots_6_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_prs1_busy = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_prs1_busy :
    issue_slots_6_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_prs2_busy = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_prs2_busy :
    issue_slots_6_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_prs3_busy = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_prs3_busy :
    issue_slots_6_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ppred_busy = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ppred_busy :
    issue_slots_6_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_stale_pdst = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_stale_pdst :
    issue_slots_6_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_exception = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_exception :
    issue_slots_6_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_exc_cause = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_exc_cause :
    issue_slots_6_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_bypassable = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_bypassable :
    issue_slots_6_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_mem_cmd = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_mem_cmd :
    issue_slots_6_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_mem_size = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_mem_size :
    issue_slots_6_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_mem_signed = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_mem_signed :
    issue_slots_6_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_fence = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_is_fence :
    issue_slots_6_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_fencei = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_is_fencei :
    issue_slots_6_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_amo = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_is_amo :
    issue_slots_6_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_uses_ldq = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_uses_ldq :
    issue_slots_6_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_uses_stq = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_uses_stq :
    issue_slots_6_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_sys_pc2epc = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_is_sys_pc2epc :
    issue_slots_6_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_unique = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_is_unique :
    issue_slots_6_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_flush_on_commit = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_flush_on_commit :
    issue_slots_6_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ldst_is_rs1 = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ldst_is_rs1 :
    issue_slots_6_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ldst = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ldst : issue_slots_6_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_lrs1 = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_lrs1 : issue_slots_6_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_lrs2 = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_lrs2 : issue_slots_6_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_lrs3 = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_lrs3 : issue_slots_6_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ldst_val = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_ldst_val :
    issue_slots_6_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_dst_rtype = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_dst_rtype :
    issue_slots_6_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_lrs1_rtype = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_lrs1_rtype :
    issue_slots_6_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_lrs2_rtype = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_lrs2_rtype :
    issue_slots_6_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_frs3_en = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_frs3_en :
    issue_slots_6_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_fp_val = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_fp_val :
    issue_slots_6_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_fp_single = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_fp_single :
    issue_slots_6_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_xcpt_pf_if = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_xcpt_pf_if :
    issue_slots_6_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_xcpt_ae_if = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_xcpt_ae_if :
    issue_slots_6_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_xcpt_ma_if = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_xcpt_ma_if :
    issue_slots_6_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_bp_debug_if = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_bp_debug_if :
    issue_slots_6_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_bp_xcpt_if = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_bp_xcpt_if :
    issue_slots_6_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_debug_fsrc = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_debug_fsrc :
    issue_slots_6_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_debug_tsrc = _GEN_23[1:0] == 2'h2 ? issue_slots_7_out_uop_debug_tsrc :
    issue_slots_6_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_clock = clock;
  assign slots_6_reset = reset;
  assign slots_6_io_grant = _T_369 & ~_T_355; // @[issue-unit-age-ordered.scala 118:56]
  assign slots_6_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_6_io_kill = io_flush_pipeline; // @[issue-unit.scala 154:28 issue-unit.scala 162:37]
  assign slots_6_io_clear = _GEN_21[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_6_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 154:28 issue-unit.scala 160:37]
  assign slots_6_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_6_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_6_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_6_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_6_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_6_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_6_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_6_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_6_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_6_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_6_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_6_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_6_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_6_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_6_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_6_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_6_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_6_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_6_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_6_io_in_uop_valid = _GEN_25[1:0] == 2'h2 ? issue_slots_8_will_be_valid : _GEN_996; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_6_io_in_uop_bits_uopc = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_uopc : issue_slots_7_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_inst = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_inst : issue_slots_7_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_debug_inst = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_debug_inst :
    issue_slots_7_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_rvc = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_is_rvc :
    issue_slots_7_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_debug_pc = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_debug_pc :
    issue_slots_7_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_iq_type = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_iq_type :
    issue_slots_7_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_fu_code = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_fu_code :
    issue_slots_7_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_br_type = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_br_type :
    issue_slots_7_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_op1_sel = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_op1_sel :
    issue_slots_7_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_op2_sel = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_op2_sel :
    issue_slots_7_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_imm_sel = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_imm_sel :
    issue_slots_7_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_op_fcn = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_op_fcn :
    issue_slots_7_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_fcn_dw = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_fcn_dw :
    issue_slots_7_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_csr_cmd = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_csr_cmd :
    issue_slots_7_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_is_load = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_is_load :
    issue_slots_7_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_is_sta = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_is_sta :
    issue_slots_7_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_is_std = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_is_std :
    issue_slots_7_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_iw_state = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_iw_state :
    issue_slots_7_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_iw_p1_poisoned = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_iw_p1_poisoned :
    issue_slots_7_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_iw_p2_poisoned = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_iw_p2_poisoned :
    issue_slots_7_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_br = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_is_br : issue_slots_7_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_jalr = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_is_jalr :
    issue_slots_7_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_jal = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_is_jal :
    issue_slots_7_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_sfb = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_is_sfb :
    issue_slots_7_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_br_mask = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_br_mask :
    issue_slots_7_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_br_tag = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_br_tag :
    issue_slots_7_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ftq_idx = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ftq_idx :
    issue_slots_7_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_edge_inst = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_edge_inst :
    issue_slots_7_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_pc_lob = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_pc_lob :
    issue_slots_7_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_taken = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_taken : issue_slots_7_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_imm_packed = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_imm_packed :
    issue_slots_7_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_csr_addr = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_csr_addr :
    issue_slots_7_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_rob_idx = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_rob_idx :
    issue_slots_7_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ldq_idx = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ldq_idx :
    issue_slots_7_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_stq_idx = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_stq_idx :
    issue_slots_7_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_rxq_idx = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_rxq_idx :
    issue_slots_7_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_pdst = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_pdst : issue_slots_7_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_prs1 = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_prs1 : issue_slots_7_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_prs2 = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_prs2 : issue_slots_7_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_prs3 = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_prs3 : issue_slots_7_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ppred = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ppred : issue_slots_7_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_prs1_busy = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_prs1_busy :
    issue_slots_7_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_prs2_busy = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_prs2_busy :
    issue_slots_7_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_prs3_busy = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_prs3_busy :
    issue_slots_7_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ppred_busy = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ppred_busy :
    issue_slots_7_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_stale_pdst = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_stale_pdst :
    issue_slots_7_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_exception = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_exception :
    issue_slots_7_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_exc_cause = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_exc_cause :
    issue_slots_7_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_bypassable = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_bypassable :
    issue_slots_7_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_mem_cmd = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_mem_cmd :
    issue_slots_7_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_mem_size = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_mem_size :
    issue_slots_7_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_mem_signed = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_mem_signed :
    issue_slots_7_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_fence = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_is_fence :
    issue_slots_7_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_fencei = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_is_fencei :
    issue_slots_7_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_amo = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_is_amo :
    issue_slots_7_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_uses_ldq = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_uses_ldq :
    issue_slots_7_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_uses_stq = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_uses_stq :
    issue_slots_7_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_sys_pc2epc = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_is_sys_pc2epc :
    issue_slots_7_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_unique = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_is_unique :
    issue_slots_7_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_flush_on_commit = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_flush_on_commit :
    issue_slots_7_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ldst_is_rs1 = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ldst_is_rs1 :
    issue_slots_7_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ldst = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ldst : issue_slots_7_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_lrs1 = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_lrs1 : issue_slots_7_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_lrs2 = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_lrs2 : issue_slots_7_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_lrs3 = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_lrs3 : issue_slots_7_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ldst_val = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_ldst_val :
    issue_slots_7_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_dst_rtype = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_dst_rtype :
    issue_slots_7_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_lrs1_rtype = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_lrs1_rtype :
    issue_slots_7_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_lrs2_rtype = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_lrs2_rtype :
    issue_slots_7_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_frs3_en = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_frs3_en :
    issue_slots_7_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_fp_val = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_fp_val :
    issue_slots_7_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_fp_single = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_fp_single :
    issue_slots_7_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_xcpt_pf_if = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_xcpt_pf_if :
    issue_slots_7_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_xcpt_ae_if = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_xcpt_ae_if :
    issue_slots_7_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_xcpt_ma_if = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_xcpt_ma_if :
    issue_slots_7_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_bp_debug_if = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_bp_debug_if :
    issue_slots_7_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_bp_xcpt_if = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_bp_xcpt_if :
    issue_slots_7_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_debug_fsrc = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_debug_fsrc :
    issue_slots_7_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_debug_tsrc = _GEN_25[1:0] == 2'h2 ? issue_slots_8_out_uop_debug_tsrc :
    issue_slots_7_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_clock = clock;
  assign slots_7_reset = reset;
  assign slots_7_io_grant = issue_slots_7_request & _T_376 & ~_T_370; // @[issue-unit-age-ordered.scala 118:56]
  assign slots_7_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_7_io_kill = io_flush_pipeline; // @[issue-unit.scala 154:28 issue-unit.scala 162:37]
  assign slots_7_io_clear = _GEN_23[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_7_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 154:28 issue-unit.scala 160:37]
  assign slots_7_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_7_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_7_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_7_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_7_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_7_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_7_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_7_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_7_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_7_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_7_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_7_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_7_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_7_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_7_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_7_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_7_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_7_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_7_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_7_io_in_uop_valid = _GEN_27[1:0] == 2'h2 ? issue_slots_9_will_be_valid : _GEN_1156; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_7_io_in_uop_bits_uopc = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_uopc : issue_slots_8_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_inst = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_inst : issue_slots_8_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_debug_inst = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_debug_inst :
    issue_slots_8_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_rvc = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_is_rvc :
    issue_slots_8_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_debug_pc = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_debug_pc :
    issue_slots_8_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_iq_type = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_iq_type :
    issue_slots_8_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_fu_code = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_fu_code :
    issue_slots_8_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_br_type = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_br_type :
    issue_slots_8_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_op1_sel = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_op1_sel :
    issue_slots_8_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_op2_sel = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_op2_sel :
    issue_slots_8_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_imm_sel = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_imm_sel :
    issue_slots_8_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_op_fcn = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_op_fcn :
    issue_slots_8_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_fcn_dw = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_fcn_dw :
    issue_slots_8_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_csr_cmd = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_csr_cmd :
    issue_slots_8_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_is_load = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_is_load :
    issue_slots_8_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_is_sta = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_is_sta :
    issue_slots_8_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_is_std = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_is_std :
    issue_slots_8_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_iw_state = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_iw_state :
    issue_slots_8_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_iw_p1_poisoned = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_iw_p1_poisoned :
    issue_slots_8_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_iw_p2_poisoned = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_iw_p2_poisoned :
    issue_slots_8_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_br = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_is_br : issue_slots_8_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_jalr = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_is_jalr :
    issue_slots_8_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_jal = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_is_jal :
    issue_slots_8_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_sfb = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_is_sfb :
    issue_slots_8_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_br_mask = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_br_mask :
    issue_slots_8_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_br_tag = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_br_tag :
    issue_slots_8_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ftq_idx = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ftq_idx :
    issue_slots_8_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_edge_inst = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_edge_inst :
    issue_slots_8_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_pc_lob = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_pc_lob :
    issue_slots_8_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_taken = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_taken : issue_slots_8_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_imm_packed = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_imm_packed :
    issue_slots_8_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_csr_addr = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_csr_addr :
    issue_slots_8_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_rob_idx = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_rob_idx :
    issue_slots_8_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ldq_idx = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ldq_idx :
    issue_slots_8_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_stq_idx = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_stq_idx :
    issue_slots_8_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_rxq_idx = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_rxq_idx :
    issue_slots_8_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_pdst = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_pdst : issue_slots_8_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_prs1 = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_prs1 : issue_slots_8_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_prs2 = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_prs2 : issue_slots_8_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_prs3 = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_prs3 : issue_slots_8_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ppred = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ppred : issue_slots_8_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_prs1_busy = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_prs1_busy :
    issue_slots_8_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_prs2_busy = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_prs2_busy :
    issue_slots_8_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_prs3_busy = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_prs3_busy :
    issue_slots_8_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ppred_busy = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ppred_busy :
    issue_slots_8_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_stale_pdst = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_stale_pdst :
    issue_slots_8_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_exception = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_exception :
    issue_slots_8_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_exc_cause = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_exc_cause :
    issue_slots_8_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_bypassable = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_bypassable :
    issue_slots_8_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_mem_cmd = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_mem_cmd :
    issue_slots_8_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_mem_size = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_mem_size :
    issue_slots_8_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_mem_signed = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_mem_signed :
    issue_slots_8_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_fence = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_is_fence :
    issue_slots_8_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_fencei = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_is_fencei :
    issue_slots_8_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_amo = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_is_amo :
    issue_slots_8_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_uses_ldq = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_uses_ldq :
    issue_slots_8_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_uses_stq = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_uses_stq :
    issue_slots_8_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_sys_pc2epc = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_is_sys_pc2epc :
    issue_slots_8_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_unique = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_is_unique :
    issue_slots_8_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_flush_on_commit = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_flush_on_commit :
    issue_slots_8_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ldst_is_rs1 = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ldst_is_rs1 :
    issue_slots_8_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ldst = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ldst : issue_slots_8_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_lrs1 = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_lrs1 : issue_slots_8_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_lrs2 = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_lrs2 : issue_slots_8_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_lrs3 = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_lrs3 : issue_slots_8_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ldst_val = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_ldst_val :
    issue_slots_8_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_dst_rtype = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_dst_rtype :
    issue_slots_8_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_lrs1_rtype = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_lrs1_rtype :
    issue_slots_8_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_lrs2_rtype = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_lrs2_rtype :
    issue_slots_8_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_frs3_en = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_frs3_en :
    issue_slots_8_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_fp_val = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_fp_val :
    issue_slots_8_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_fp_single = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_fp_single :
    issue_slots_8_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_xcpt_pf_if = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_xcpt_pf_if :
    issue_slots_8_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_xcpt_ae_if = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_xcpt_ae_if :
    issue_slots_8_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_xcpt_ma_if = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_xcpt_ma_if :
    issue_slots_8_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_bp_debug_if = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_bp_debug_if :
    issue_slots_8_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_bp_xcpt_if = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_bp_xcpt_if :
    issue_slots_8_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_debug_fsrc = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_debug_fsrc :
    issue_slots_8_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_debug_tsrc = _GEN_27[1:0] == 2'h2 ? issue_slots_9_out_uop_debug_tsrc :
    issue_slots_8_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_clock = clock;
  assign slots_8_reset = reset;
  assign slots_8_io_grant = issue_slots_8_request & _T_391 & ~_T_385; // @[issue-unit-age-ordered.scala 118:56]
  assign slots_8_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_8_io_kill = io_flush_pipeline; // @[issue-unit.scala 154:28 issue-unit.scala 162:37]
  assign slots_8_io_clear = _GEN_25[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_8_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 154:28 issue-unit.scala 160:37]
  assign slots_8_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_8_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_8_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_8_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_8_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_8_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_8_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_8_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_8_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_8_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_8_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_8_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_8_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_8_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_8_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_8_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_8_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_8_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_8_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_8_io_in_uop_valid = _GEN_29[1:0] == 2'h2 ? issue_slots_10_will_be_valid : _GEN_1316; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_8_io_in_uop_bits_uopc = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_uopc : issue_slots_9_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_inst = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_inst : issue_slots_9_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_debug_inst = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_debug_inst :
    issue_slots_9_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_rvc = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_is_rvc :
    issue_slots_9_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_debug_pc = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_debug_pc :
    issue_slots_9_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_iq_type = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_iq_type :
    issue_slots_9_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_fu_code = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_fu_code :
    issue_slots_9_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_br_type = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_br_type :
    issue_slots_9_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_op1_sel = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_op1_sel :
    issue_slots_9_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_op2_sel = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_op2_sel :
    issue_slots_9_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_imm_sel = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_imm_sel :
    issue_slots_9_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_op_fcn = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_op_fcn :
    issue_slots_9_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_fcn_dw = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_fcn_dw :
    issue_slots_9_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_csr_cmd = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_csr_cmd :
    issue_slots_9_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_is_load = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_is_load :
    issue_slots_9_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_is_sta = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_is_sta :
    issue_slots_9_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_is_std = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_is_std :
    issue_slots_9_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_iw_state = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_iw_state :
    issue_slots_9_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_iw_p1_poisoned = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_iw_p1_poisoned :
    issue_slots_9_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_iw_p2_poisoned = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_iw_p2_poisoned :
    issue_slots_9_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_br = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_is_br :
    issue_slots_9_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_jalr = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_is_jalr :
    issue_slots_9_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_jal = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_is_jal :
    issue_slots_9_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_sfb = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_is_sfb :
    issue_slots_9_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_br_mask = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_br_mask :
    issue_slots_9_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_br_tag = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_br_tag :
    issue_slots_9_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ftq_idx = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ftq_idx :
    issue_slots_9_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_edge_inst = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_edge_inst :
    issue_slots_9_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_pc_lob = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_pc_lob :
    issue_slots_9_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_taken = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_taken :
    issue_slots_9_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_imm_packed = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_imm_packed :
    issue_slots_9_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_csr_addr = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_csr_addr :
    issue_slots_9_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_rob_idx = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_rob_idx :
    issue_slots_9_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ldq_idx = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ldq_idx :
    issue_slots_9_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_stq_idx = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_stq_idx :
    issue_slots_9_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_rxq_idx = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_rxq_idx :
    issue_slots_9_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_pdst = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_pdst : issue_slots_9_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_prs1 = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_prs1 : issue_slots_9_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_prs2 = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_prs2 : issue_slots_9_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_prs3 = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_prs3 : issue_slots_9_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ppred = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ppred :
    issue_slots_9_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_prs1_busy = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_prs1_busy :
    issue_slots_9_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_prs2_busy = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_prs2_busy :
    issue_slots_9_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_prs3_busy = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_prs3_busy :
    issue_slots_9_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ppred_busy = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ppred_busy :
    issue_slots_9_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_stale_pdst = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_stale_pdst :
    issue_slots_9_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_exception = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_exception :
    issue_slots_9_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_exc_cause = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_exc_cause :
    issue_slots_9_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_bypassable = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_bypassable :
    issue_slots_9_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_mem_cmd = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_mem_cmd :
    issue_slots_9_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_mem_size = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_mem_size :
    issue_slots_9_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_mem_signed = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_mem_signed :
    issue_slots_9_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_fence = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_is_fence :
    issue_slots_9_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_fencei = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_is_fencei :
    issue_slots_9_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_amo = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_is_amo :
    issue_slots_9_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_uses_ldq = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_uses_ldq :
    issue_slots_9_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_uses_stq = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_uses_stq :
    issue_slots_9_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_sys_pc2epc = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_is_sys_pc2epc :
    issue_slots_9_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_unique = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_is_unique :
    issue_slots_9_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_flush_on_commit = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_flush_on_commit :
    issue_slots_9_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ldst_is_rs1 = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ldst_is_rs1 :
    issue_slots_9_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ldst = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ldst : issue_slots_9_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_lrs1 = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_lrs1 : issue_slots_9_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_lrs2 = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_lrs2 : issue_slots_9_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_lrs3 = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_lrs3 : issue_slots_9_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ldst_val = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_ldst_val :
    issue_slots_9_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_dst_rtype = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_dst_rtype :
    issue_slots_9_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_lrs1_rtype = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_lrs1_rtype :
    issue_slots_9_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_lrs2_rtype = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_lrs2_rtype :
    issue_slots_9_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_frs3_en = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_frs3_en :
    issue_slots_9_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_fp_val = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_fp_val :
    issue_slots_9_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_fp_single = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_fp_single :
    issue_slots_9_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_xcpt_pf_if = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_xcpt_pf_if :
    issue_slots_9_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_xcpt_ae_if = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_xcpt_ae_if :
    issue_slots_9_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_xcpt_ma_if = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_xcpt_ma_if :
    issue_slots_9_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_bp_debug_if = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_bp_debug_if :
    issue_slots_9_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_bp_xcpt_if = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_bp_xcpt_if :
    issue_slots_9_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_debug_fsrc = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_debug_fsrc :
    issue_slots_9_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_debug_tsrc = _GEN_29[1:0] == 2'h2 ? issue_slots_10_out_uop_debug_tsrc :
    issue_slots_9_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_clock = clock;
  assign slots_9_reset = reset;
  assign slots_9_io_grant = _T_414 & ~_T_400; // @[issue-unit-age-ordered.scala 118:56]
  assign slots_9_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_9_io_kill = io_flush_pipeline; // @[issue-unit.scala 154:28 issue-unit.scala 162:37]
  assign slots_9_io_clear = _GEN_27[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_9_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 154:28 issue-unit.scala 160:37]
  assign slots_9_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_9_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_9_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_9_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_9_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_9_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_9_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_9_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_9_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_9_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_9_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_9_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_9_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_9_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_9_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_9_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_9_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_9_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_9_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_9_io_in_uop_valid = _GEN_31[1:0] == 2'h2 ? issue_slots_11_will_be_valid : _GEN_1476; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_9_io_in_uop_bits_uopc = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_uopc : issue_slots_10_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_inst = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_inst : issue_slots_10_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_debug_inst = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_debug_inst :
    issue_slots_10_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_rvc = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_is_rvc :
    issue_slots_10_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_debug_pc = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_debug_pc :
    issue_slots_10_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_iq_type = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_iq_type :
    issue_slots_10_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_fu_code = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_fu_code :
    issue_slots_10_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_br_type = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_br_type :
    issue_slots_10_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_op1_sel = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_op1_sel :
    issue_slots_10_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_op2_sel = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_op2_sel :
    issue_slots_10_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_imm_sel = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_imm_sel :
    issue_slots_10_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_op_fcn = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_op_fcn :
    issue_slots_10_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_fcn_dw = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_fcn_dw :
    issue_slots_10_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_csr_cmd = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_csr_cmd :
    issue_slots_10_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_is_load = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_is_load :
    issue_slots_10_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_is_sta = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_is_sta :
    issue_slots_10_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_is_std = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_is_std :
    issue_slots_10_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_iw_state = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_iw_state :
    issue_slots_10_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_iw_p1_poisoned = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_iw_p1_poisoned :
    issue_slots_10_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_iw_p2_poisoned = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_iw_p2_poisoned :
    issue_slots_10_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_br = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_is_br :
    issue_slots_10_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_jalr = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_is_jalr :
    issue_slots_10_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_jal = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_is_jal :
    issue_slots_10_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_sfb = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_is_sfb :
    issue_slots_10_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_br_mask = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_br_mask :
    issue_slots_10_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_br_tag = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_br_tag :
    issue_slots_10_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ftq_idx = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ftq_idx :
    issue_slots_10_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_edge_inst = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_edge_inst :
    issue_slots_10_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_pc_lob = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_pc_lob :
    issue_slots_10_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_taken = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_taken :
    issue_slots_10_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_imm_packed = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_imm_packed :
    issue_slots_10_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_csr_addr = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_csr_addr :
    issue_slots_10_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_rob_idx = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_rob_idx :
    issue_slots_10_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ldq_idx = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ldq_idx :
    issue_slots_10_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_stq_idx = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_stq_idx :
    issue_slots_10_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_rxq_idx = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_rxq_idx :
    issue_slots_10_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_pdst = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_pdst : issue_slots_10_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_prs1 = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_prs1 : issue_slots_10_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_prs2 = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_prs2 : issue_slots_10_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_prs3 = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_prs3 : issue_slots_10_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ppred = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ppred :
    issue_slots_10_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_prs1_busy = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_prs1_busy :
    issue_slots_10_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_prs2_busy = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_prs2_busy :
    issue_slots_10_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_prs3_busy = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_prs3_busy :
    issue_slots_10_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ppred_busy = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ppred_busy :
    issue_slots_10_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_stale_pdst = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_stale_pdst :
    issue_slots_10_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_exception = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_exception :
    issue_slots_10_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_exc_cause = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_exc_cause :
    issue_slots_10_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_bypassable = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_bypassable :
    issue_slots_10_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_mem_cmd = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_mem_cmd :
    issue_slots_10_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_mem_size = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_mem_size :
    issue_slots_10_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_mem_signed = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_mem_signed :
    issue_slots_10_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_fence = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_is_fence :
    issue_slots_10_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_fencei = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_is_fencei :
    issue_slots_10_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_amo = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_is_amo :
    issue_slots_10_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_uses_ldq = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_uses_ldq :
    issue_slots_10_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_uses_stq = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_uses_stq :
    issue_slots_10_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_sys_pc2epc = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_is_sys_pc2epc :
    issue_slots_10_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_unique = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_is_unique :
    issue_slots_10_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_flush_on_commit = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_flush_on_commit :
    issue_slots_10_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ldst_is_rs1 = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ldst_is_rs1 :
    issue_slots_10_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ldst = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ldst : issue_slots_10_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_lrs1 = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_lrs1 : issue_slots_10_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_lrs2 = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_lrs2 : issue_slots_10_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_lrs3 = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_lrs3 : issue_slots_10_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ldst_val = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_ldst_val :
    issue_slots_10_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_dst_rtype = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_dst_rtype :
    issue_slots_10_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_lrs1_rtype = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_lrs1_rtype :
    issue_slots_10_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_lrs2_rtype = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_lrs2_rtype :
    issue_slots_10_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_frs3_en = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_frs3_en :
    issue_slots_10_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_fp_val = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_fp_val :
    issue_slots_10_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_fp_single = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_fp_single :
    issue_slots_10_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_xcpt_pf_if = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_xcpt_pf_if :
    issue_slots_10_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_xcpt_ae_if = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_xcpt_ae_if :
    issue_slots_10_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_xcpt_ma_if = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_xcpt_ma_if :
    issue_slots_10_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_bp_debug_if = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_bp_debug_if :
    issue_slots_10_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_bp_xcpt_if = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_bp_xcpt_if :
    issue_slots_10_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_debug_fsrc = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_debug_fsrc :
    issue_slots_10_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_debug_tsrc = _GEN_31[1:0] == 2'h2 ? issue_slots_11_out_uop_debug_tsrc :
    issue_slots_10_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_clock = clock;
  assign slots_10_reset = reset;
  assign slots_10_io_grant = issue_slots_10_request & _T_421 & ~_T_415; // @[issue-unit-age-ordered.scala 118:56]
  assign slots_10_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_10_io_kill = io_flush_pipeline; // @[issue-unit.scala 154:28 issue-unit.scala 162:37]
  assign slots_10_io_clear = _GEN_29[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_10_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 154:28 issue-unit.scala 160:37]
  assign slots_10_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_10_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_10_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_10_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_10_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_10_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_10_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_10_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_10_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_10_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_10_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_10_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_10_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_10_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_10_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_10_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_10_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_10_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_10_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_10_io_in_uop_valid = _GEN_33[1:0] == 2'h2 ? will_be_valid_12 : _GEN_1636; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_10_io_in_uop_bits_uopc = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_uopc : issue_slots_11_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_inst = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_inst : issue_slots_11_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_debug_inst = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_debug_inst :
    issue_slots_11_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_rvc = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_is_rvc :
    issue_slots_11_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_debug_pc = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_debug_pc :
    issue_slots_11_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_iq_type = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_iq_type :
    issue_slots_11_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_fu_code = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_fu_code :
    issue_slots_11_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_br_type = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_br_type :
    issue_slots_11_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_op1_sel = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_op1_sel :
    issue_slots_11_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_op2_sel = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_op2_sel :
    issue_slots_11_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_imm_sel = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_imm_sel :
    issue_slots_11_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_op_fcn = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_op_fcn :
    issue_slots_11_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_fcn_dw = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_fcn_dw :
    issue_slots_11_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_csr_cmd = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_csr_cmd :
    issue_slots_11_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_is_load = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_is_load :
    issue_slots_11_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_is_sta = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_is_sta :
    issue_slots_11_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_is_std = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_is_std :
    issue_slots_11_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_iw_state = _GEN_33[1:0] == 2'h2 ? uops_12_iw_state : issue_slots_11_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_iw_p1_poisoned = _GEN_33[1:0] == 2'h2 ? 1'h0 : issue_slots_11_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_iw_p2_poisoned = _GEN_33[1:0] == 2'h2 ? 1'h0 : issue_slots_11_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_br = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_is_br : issue_slots_11_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_jalr = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_is_jalr :
    issue_slots_11_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_jal = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_is_jal :
    issue_slots_11_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_sfb = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_is_sfb :
    issue_slots_11_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_br_mask = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_br_mask :
    issue_slots_11_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_br_tag = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_br_tag :
    issue_slots_11_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ftq_idx = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_ftq_idx :
    issue_slots_11_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_edge_inst = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_edge_inst :
    issue_slots_11_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_pc_lob = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_pc_lob :
    issue_slots_11_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_taken = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_taken : issue_slots_11_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_imm_packed = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_imm_packed :
    issue_slots_11_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_csr_addr = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_csr_addr :
    issue_slots_11_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_rob_idx = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_rob_idx :
    issue_slots_11_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ldq_idx = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_ldq_idx :
    issue_slots_11_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_stq_idx = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_stq_idx :
    issue_slots_11_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_rxq_idx = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_rxq_idx :
    issue_slots_11_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_pdst = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_pdst : issue_slots_11_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_prs1 = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_prs1 : issue_slots_11_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_prs2 = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_prs2 : issue_slots_11_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_prs3 = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_prs3 : issue_slots_11_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ppred = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_ppred : issue_slots_11_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_prs1_busy = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_prs1_busy :
    issue_slots_11_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_prs2_busy = _GEN_33[1:0] == 2'h2 ? uops_12_prs2_busy : issue_slots_11_out_uop_prs2_busy
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_prs3_busy = _GEN_33[1:0] == 2'h2 ? 1'h0 : issue_slots_11_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ppred_busy = _GEN_33[1:0] == 2'h2 ? 1'h0 : issue_slots_11_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_stale_pdst = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_stale_pdst :
    issue_slots_11_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_exception = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_exception :
    issue_slots_11_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_exc_cause = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_exc_cause :
    issue_slots_11_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_bypassable = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_bypassable :
    issue_slots_11_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_mem_cmd = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_mem_cmd :
    issue_slots_11_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_mem_size = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_mem_size :
    issue_slots_11_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_mem_signed = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_mem_signed :
    issue_slots_11_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_fence = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_is_fence :
    issue_slots_11_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_fencei = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_is_fencei :
    issue_slots_11_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_amo = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_is_amo :
    issue_slots_11_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_uses_ldq = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_uses_ldq :
    issue_slots_11_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_uses_stq = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_uses_stq :
    issue_slots_11_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_sys_pc2epc = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_is_sys_pc2epc :
    issue_slots_11_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_unique = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_is_unique :
    issue_slots_11_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_flush_on_commit = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_flush_on_commit :
    issue_slots_11_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ldst_is_rs1 = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_ldst_is_rs1 :
    issue_slots_11_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ldst = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_ldst : issue_slots_11_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_lrs1 = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_lrs1 : issue_slots_11_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_lrs2 = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_lrs2 : issue_slots_11_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_lrs3 = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_lrs3 : issue_slots_11_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ldst_val = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_ldst_val :
    issue_slots_11_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_dst_rtype = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_dst_rtype :
    issue_slots_11_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_lrs1_rtype = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_lrs1_rtype :
    issue_slots_11_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_lrs2_rtype = _GEN_33[1:0] == 2'h2 ? uops_12_lrs2_rtype :
    issue_slots_11_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_frs3_en = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_frs3_en :
    issue_slots_11_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_fp_val = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_fp_val :
    issue_slots_11_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_fp_single = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_fp_single :
    issue_slots_11_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_xcpt_pf_if = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_xcpt_pf_if :
    issue_slots_11_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_xcpt_ae_if = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_xcpt_ae_if :
    issue_slots_11_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_xcpt_ma_if = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_xcpt_ma_if :
    issue_slots_11_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_bp_debug_if = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_bp_debug_if :
    issue_slots_11_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_bp_xcpt_if = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_bp_xcpt_if :
    issue_slots_11_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_debug_fsrc = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_debug_fsrc :
    issue_slots_11_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_debug_tsrc = _GEN_33[1:0] == 2'h2 ? io_dis_uops_0_bits_debug_tsrc :
    issue_slots_11_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_clock = clock;
  assign slots_11_reset = reset;
  assign slots_11_io_grant = issue_slots_11_request & _T_436 & ~_T_430; // @[issue-unit-age-ordered.scala 118:56]
  assign slots_11_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 154:28 issue-unit.scala 161:37]
  assign slots_11_io_kill = io_flush_pipeline; // @[issue-unit.scala 154:28 issue-unit.scala 162:37]
  assign slots_11_io_clear = _GEN_31[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_11_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 154:28 issue-unit.scala 160:37]
  assign slots_11_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_11_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_11_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_11_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_11_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_11_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_11_io_wakeup_ports_2_valid = io_wakeup_ports_2_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_11_io_wakeup_ports_2_bits_pdst = io_wakeup_ports_2_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_11_io_wakeup_ports_2_bits_poisoned = io_wakeup_ports_2_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_11_io_wakeup_ports_3_valid = io_wakeup_ports_3_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_11_io_wakeup_ports_3_bits_pdst = io_wakeup_ports_3_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_11_io_wakeup_ports_3_bits_poisoned = io_wakeup_ports_3_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_11_io_wakeup_ports_4_valid = io_wakeup_ports_4_valid; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_11_io_wakeup_ports_4_bits_pdst = io_wakeup_ports_4_bits_pdst; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_11_io_wakeup_ports_4_bits_poisoned = io_wakeup_ports_4_bits_poisoned; // @[issue-unit.scala 154:28 issue-unit.scala 157:37]
  assign slots_11_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_11_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 154:28 issue-unit.scala 158:37]
  assign slots_11_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_11_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 154:28 issue-unit.scala 159:37]
  assign slots_11_io_in_uop_valid = _GEN_35[1:0] == 2'h2 ? will_be_valid_13 : _GEN_1796; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_11_io_in_uop_bits_uopc = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_uopc : io_dis_uops_0_bits_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_inst = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_inst : io_dis_uops_0_bits_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_debug_inst = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_debug_inst :
    io_dis_uops_0_bits_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_rvc = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_is_rvc : io_dis_uops_0_bits_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_debug_pc = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_debug_pc :
    io_dis_uops_0_bits_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_iq_type = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_iq_type :
    io_dis_uops_0_bits_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_fu_code = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_fu_code :
    io_dis_uops_0_bits_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_br_type = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_br_type :
    io_dis_uops_0_bits_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_op1_sel = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_op1_sel :
    io_dis_uops_0_bits_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_op2_sel = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_op2_sel :
    io_dis_uops_0_bits_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_imm_sel = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_imm_sel :
    io_dis_uops_0_bits_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_op_fcn = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_op_fcn :
    io_dis_uops_0_bits_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_fcn_dw = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_fcn_dw :
    io_dis_uops_0_bits_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_csr_cmd = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_csr_cmd :
    io_dis_uops_0_bits_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_is_load = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_is_load :
    io_dis_uops_0_bits_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_is_sta = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_is_sta :
    io_dis_uops_0_bits_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_is_std = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_is_std :
    io_dis_uops_0_bits_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_iw_state = _GEN_35[1:0] == 2'h2 ? uops_13_iw_state : uops_12_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_iw_p1_poisoned = 1'h0; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_iw_p2_poisoned = 1'h0; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_br = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_is_br : io_dis_uops_0_bits_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_jalr = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_is_jalr :
    io_dis_uops_0_bits_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_jal = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_is_jal : io_dis_uops_0_bits_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_sfb = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_is_sfb : io_dis_uops_0_bits_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_br_mask = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_br_mask :
    io_dis_uops_0_bits_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_br_tag = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_br_tag : io_dis_uops_0_bits_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ftq_idx = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_ftq_idx :
    io_dis_uops_0_bits_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_edge_inst = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_edge_inst :
    io_dis_uops_0_bits_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_pc_lob = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_pc_lob : io_dis_uops_0_bits_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_taken = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_taken : io_dis_uops_0_bits_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_imm_packed = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_imm_packed :
    io_dis_uops_0_bits_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_csr_addr = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_csr_addr :
    io_dis_uops_0_bits_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_rob_idx = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_rob_idx :
    io_dis_uops_0_bits_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ldq_idx = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_ldq_idx :
    io_dis_uops_0_bits_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_stq_idx = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_stq_idx :
    io_dis_uops_0_bits_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_rxq_idx = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_rxq_idx :
    io_dis_uops_0_bits_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_pdst = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_pdst : io_dis_uops_0_bits_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_prs1 = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_prs1 : io_dis_uops_0_bits_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_prs2 = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_prs2 : io_dis_uops_0_bits_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_prs3 = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_prs3 : io_dis_uops_0_bits_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ppred = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_ppred : io_dis_uops_0_bits_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_prs1_busy = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_prs1_busy :
    io_dis_uops_0_bits_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_prs2_busy = _GEN_35[1:0] == 2'h2 ? uops_13_prs2_busy : uops_12_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_prs3_busy = 1'h0; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ppred_busy = 1'h0; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_stale_pdst = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_stale_pdst :
    io_dis_uops_0_bits_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_exception = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_exception :
    io_dis_uops_0_bits_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_exc_cause = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_exc_cause :
    io_dis_uops_0_bits_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_bypassable = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_bypassable :
    io_dis_uops_0_bits_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_mem_cmd = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_mem_cmd :
    io_dis_uops_0_bits_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_mem_size = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_mem_size :
    io_dis_uops_0_bits_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_mem_signed = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_mem_signed :
    io_dis_uops_0_bits_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_fence = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_is_fence :
    io_dis_uops_0_bits_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_fencei = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_is_fencei :
    io_dis_uops_0_bits_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_amo = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_is_amo : io_dis_uops_0_bits_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_uses_ldq = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_uses_ldq :
    io_dis_uops_0_bits_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_uses_stq = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_uses_stq :
    io_dis_uops_0_bits_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_sys_pc2epc = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_is_sys_pc2epc :
    io_dis_uops_0_bits_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_unique = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_is_unique :
    io_dis_uops_0_bits_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_flush_on_commit = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_flush_on_commit :
    io_dis_uops_0_bits_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ldst_is_rs1 = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_ldst_is_rs1 :
    io_dis_uops_0_bits_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ldst = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_ldst : io_dis_uops_0_bits_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_lrs1 = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_lrs1 : io_dis_uops_0_bits_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_lrs2 = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_lrs2 : io_dis_uops_0_bits_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_lrs3 = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_lrs3 : io_dis_uops_0_bits_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ldst_val = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_ldst_val :
    io_dis_uops_0_bits_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_dst_rtype = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_dst_rtype :
    io_dis_uops_0_bits_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_lrs1_rtype = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_lrs1_rtype :
    io_dis_uops_0_bits_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_lrs2_rtype = _GEN_35[1:0] == 2'h2 ? uops_13_lrs2_rtype : uops_12_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_frs3_en = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_frs3_en :
    io_dis_uops_0_bits_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_fp_val = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_fp_val : io_dis_uops_0_bits_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_fp_single = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_fp_single :
    io_dis_uops_0_bits_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_xcpt_pf_if = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_xcpt_pf_if :
    io_dis_uops_0_bits_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_xcpt_ae_if = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_xcpt_ae_if :
    io_dis_uops_0_bits_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_xcpt_ma_if = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_xcpt_ma_if :
    io_dis_uops_0_bits_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_bp_debug_if = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_bp_debug_if :
    io_dis_uops_0_bits_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_bp_xcpt_if = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_bp_xcpt_if :
    io_dis_uops_0_bits_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_debug_fsrc = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_debug_fsrc :
    io_dis_uops_0_bits_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_debug_tsrc = _GEN_35[1:0] == 2'h2 ? io_dis_uops_1_bits_debug_tsrc :
    io_dis_uops_0_bits_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  always @(posedge clock) begin
    REG <= num_available > 4'h0; // @[issue-unit-age-ordered.scala 87:51]
    REG_1 <= num_available > 4'h1; // @[issue-unit-age-ordered.scala 87:51]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_dis_uops_0_bits_ppred_busy & io_dis_uops_0_valid) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at issue-unit.scala:145 assert(!(io.dis_uops(w).bits.ppred_busy && io.dis_uops(w).valid))\n"
            ); // @[issue-unit.scala 145:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_dis_uops_0_bits_ppred_busy & io_dis_uops_0_valid) | reset)) begin
          $fatal; // @[issue-unit.scala 145:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_dis_uops_1_bits_ppred_busy & io_dis_uops_1_valid) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at issue-unit.scala:145 assert(!(io.dis_uops(w).bits.ppred_busy && io.dis_uops(w).valid))\n"
            ); // @[issue-unit.scala 145:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_dis_uops_1_bits_ppred_busy & io_dis_uops_1_valid) | reset)) begin
          $fatal; // @[issue-unit.scala 145:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_79 <= 4'h1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [issue] window giving out too many grants.\n    at issue-unit.scala:172 assert (PopCount(issue_slots.map(s => s.grant)) <= issueWidth.U, \"[issue] window giving out too many grants.\")\n"
            ); // @[issue-unit.scala 172:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_79 <= 4'h1 | reset)) begin
          $fatal; // @[issue-unit.scala 172:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG_1 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
