module BundleBridgeNexus_15(
  input         clock,
  input         reset,
  input         auto_in_group_0_iretire,
  input  [31:0] auto_in_group_0_iaddr,
  input  [3:0]  auto_in_group_0_itype,
  input         auto_in_group_0_ilastsize,
  input  [3:0]  auto_in_priv,
  input  [31:0] auto_in_tval,
  input  [31:0] auto_in_cause
);
endmodule
