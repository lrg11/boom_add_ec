module RoundAnyRawFNToRecFN_7(
  input         io_invalidExc,
  input         io_infiniteExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [12:0] io_in_sExp,
  input  [55:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags
);
  wire  roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  roundMagUp = roundingMode_min & io_in_sign | roundingMode_max & ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:42]
  wire [11:0] _roundMask_T_1 = ~io_in_sExp[11:0]; // @[primitives.scala 51:21]
  wire  roundMask_msb = _roundMask_T_1[11]; // @[primitives.scala 57:25]
  wire [10:0] roundMask_lsbs = _roundMask_T_1[10:0]; // @[primitives.scala 58:26]
  wire  roundMask_msb_1 = roundMask_lsbs[10]; // @[primitives.scala 57:25]
  wire [9:0] roundMask_lsbs_1 = roundMask_lsbs[9:0]; // @[primitives.scala 58:26]
  wire  roundMask_msb_2 = roundMask_lsbs_1[9]; // @[primitives.scala 57:25]
  wire [8:0] roundMask_lsbs_2 = roundMask_lsbs_1[8:0]; // @[primitives.scala 58:26]
  wire  roundMask_msb_3 = roundMask_lsbs_2[8]; // @[primitives.scala 57:25]
  wire [7:0] roundMask_lsbs_3 = roundMask_lsbs_2[7:0]; // @[primitives.scala 58:26]
  wire  roundMask_msb_4 = roundMask_lsbs_3[7]; // @[primitives.scala 57:25]
  wire [6:0] roundMask_lsbs_4 = roundMask_lsbs_3[6:0]; // @[primitives.scala 58:26]
  wire  roundMask_msb_5 = roundMask_lsbs_4[6]; // @[primitives.scala 57:25]
  wire [5:0] roundMask_lsbs_5 = roundMask_lsbs_4[5:0]; // @[primitives.scala 58:26]
  wire [64:0] roundMask_shift = 65'sh10000000000000000 >>> roundMask_lsbs_5; // @[primitives.scala 77:58]
  wire [31:0] _roundMask_T_7 = {{16'd0}, roundMask_shift[44:29]}; // @[Bitwise.scala 103:31]
  wire [31:0] _roundMask_T_9 = {roundMask_shift[28:13], 16'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _roundMask_T_11 = _roundMask_T_9 & 32'hffff0000; // @[Bitwise.scala 103:75]
  wire [31:0] _roundMask_T_12 = _roundMask_T_7 | _roundMask_T_11; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_0 = {{8'd0}, _roundMask_T_12[31:8]}; // @[Bitwise.scala 103:31]
  wire [31:0] _roundMask_T_17 = _GEN_0 & 32'hff00ff; // @[Bitwise.scala 103:31]
  wire [31:0] _roundMask_T_19 = {_roundMask_T_12[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _roundMask_T_21 = _roundMask_T_19 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  wire [31:0] _roundMask_T_22 = _roundMask_T_17 | _roundMask_T_21; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1 = {{4'd0}, _roundMask_T_22[31:4]}; // @[Bitwise.scala 103:31]
  wire [31:0] _roundMask_T_27 = _GEN_1 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  wire [31:0] _roundMask_T_29 = {_roundMask_T_22[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _roundMask_T_31 = _roundMask_T_29 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  wire [31:0] _roundMask_T_32 = _roundMask_T_27 | _roundMask_T_31; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_2 = {{2'd0}, _roundMask_T_32[31:2]}; // @[Bitwise.scala 103:31]
  wire [31:0] _roundMask_T_37 = _GEN_2 & 32'h33333333; // @[Bitwise.scala 103:31]
  wire [31:0] _roundMask_T_39 = {_roundMask_T_32[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _roundMask_T_41 = _roundMask_T_39 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  wire [31:0] _roundMask_T_42 = _roundMask_T_37 | _roundMask_T_41; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_3 = {{1'd0}, _roundMask_T_42[31:1]}; // @[Bitwise.scala 103:31]
  wire [31:0] _roundMask_T_47 = _GEN_3 & 32'h55555555; // @[Bitwise.scala 103:31]
  wire [31:0] _roundMask_T_49 = {_roundMask_T_42[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _roundMask_T_51 = _roundMask_T_49 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  wire [31:0] roundMask_hi = _roundMask_T_47 | _roundMask_T_51; // @[Bitwise.scala 103:39]
  wire [15:0] _roundMask_T_57 = {{8'd0}, roundMask_shift[60:53]}; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_59 = {roundMask_shift[52:45], 8'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _roundMask_T_61 = _roundMask_T_59 & 16'hff00; // @[Bitwise.scala 103:75]
  wire [15:0] _roundMask_T_62 = _roundMask_T_57 | _roundMask_T_61; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_4 = {{4'd0}, _roundMask_T_62[15:4]}; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_67 = _GEN_4 & 16'hf0f; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_69 = {_roundMask_T_62[11:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _roundMask_T_71 = _roundMask_T_69 & 16'hf0f0; // @[Bitwise.scala 103:75]
  wire [15:0] _roundMask_T_72 = _roundMask_T_67 | _roundMask_T_71; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_5 = {{2'd0}, _roundMask_T_72[15:2]}; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_77 = _GEN_5 & 16'h3333; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_79 = {_roundMask_T_72[13:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _roundMask_T_81 = _roundMask_T_79 & 16'hcccc; // @[Bitwise.scala 103:75]
  wire [15:0] _roundMask_T_82 = _roundMask_T_77 | _roundMask_T_81; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_6 = {{1'd0}, _roundMask_T_82[15:1]}; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_87 = _GEN_6 & 16'h5555; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_89 = {_roundMask_T_82[14:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _roundMask_T_91 = _roundMask_T_89 & 16'haaaa; // @[Bitwise.scala 103:75]
  wire [15:0] roundMask_hi_1 = _roundMask_T_87 | _roundMask_T_91; // @[Bitwise.scala 103:39]
  wire  roundMask_hi_2 = roundMask_shift[61]; // @[Bitwise.scala 109:18]
  wire  roundMask_lo = roundMask_shift[62]; // @[Bitwise.scala 109:44]
  wire  roundMask_lo_1 = roundMask_shift[63]; // @[Bitwise.scala 109:44]
  wire [50:0] _roundMask_T_94 = {roundMask_hi,roundMask_hi_1,roundMask_hi_2,roundMask_lo,roundMask_lo_1}; // @[Cat.scala 30:58]
  wire [50:0] _roundMask_T_95 = ~_roundMask_T_94; // @[primitives.scala 74:36]
  wire [50:0] _roundMask_T_96 = roundMask_msb_5 ? 51'h0 : _roundMask_T_95; // @[primitives.scala 74:21]
  wire [50:0] _roundMask_T_97 = ~_roundMask_T_96; // @[primitives.scala 74:17]
  wire [50:0] _roundMask_T_98 = ~_roundMask_T_97; // @[primitives.scala 74:36]
  wire [50:0] _roundMask_T_99 = roundMask_msb_4 ? 51'h0 : _roundMask_T_98; // @[primitives.scala 74:21]
  wire [50:0] _roundMask_T_100 = ~_roundMask_T_99; // @[primitives.scala 74:17]
  wire [50:0] _roundMask_T_101 = ~_roundMask_T_100; // @[primitives.scala 74:36]
  wire [50:0] _roundMask_T_102 = roundMask_msb_3 ? 51'h0 : _roundMask_T_101; // @[primitives.scala 74:21]
  wire [50:0] _roundMask_T_103 = ~_roundMask_T_102; // @[primitives.scala 74:17]
  wire [50:0] _roundMask_T_104 = ~_roundMask_T_103; // @[primitives.scala 74:36]
  wire [50:0] _roundMask_T_105 = roundMask_msb_2 ? 51'h0 : _roundMask_T_104; // @[primitives.scala 74:21]
  wire [50:0] roundMask_hi_4 = ~_roundMask_T_105; // @[primitives.scala 74:17]
  wire [53:0] _roundMask_T_106 = {roundMask_hi_4,3'h7}; // @[Cat.scala 30:58]
  wire  roundMask_hi_5 = roundMask_shift[0]; // @[Bitwise.scala 109:18]
  wire  roundMask_lo_4 = roundMask_shift[1]; // @[Bitwise.scala 109:44]
  wire  roundMask_lo_5 = roundMask_shift[2]; // @[Bitwise.scala 109:44]
  wire [2:0] _roundMask_T_109 = {roundMask_hi_5,roundMask_lo_4,roundMask_lo_5}; // @[Cat.scala 30:58]
  wire [2:0] _roundMask_T_110 = roundMask_msb_5 ? _roundMask_T_109 : 3'h0; // @[primitives.scala 61:24]
  wire [2:0] _roundMask_T_111 = roundMask_msb_4 ? _roundMask_T_110 : 3'h0; // @[primitives.scala 61:24]
  wire [2:0] _roundMask_T_112 = roundMask_msb_3 ? _roundMask_T_111 : 3'h0; // @[primitives.scala 61:24]
  wire [2:0] _roundMask_T_113 = roundMask_msb_2 ? _roundMask_T_112 : 3'h0; // @[primitives.scala 61:24]
  wire [53:0] _roundMask_T_114 = roundMask_msb_1 ? _roundMask_T_106 : {{51'd0}, _roundMask_T_113}; // @[primitives.scala 66:24]
  wire [53:0] roundMask_hi_7 = roundMask_msb ? _roundMask_T_114 : 54'h0; // @[primitives.scala 61:24]
  wire [55:0] roundMask = {roundMask_hi_7,2'h3}; // @[Cat.scala 30:58]
  wire [54:0] shiftedRoundMask_lo = roundMask[55:1]; // @[RoundAnyRawFNToRecFN.scala 160:57]
  wire [55:0] shiftedRoundMask = {1'h0,shiftedRoundMask_lo}; // @[Cat.scala 30:58]
  wire [55:0] _roundPosMask_T = ~shiftedRoundMask; // @[RoundAnyRawFNToRecFN.scala 161:28]
  wire [55:0] roundPosMask = _roundPosMask_T & roundMask; // @[RoundAnyRawFNToRecFN.scala 161:46]
  wire [55:0] _roundPosBit_T = io_in_sig & roundPosMask; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  roundPosBit = |_roundPosBit_T; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [55:0] _anyRoundExtra_T = io_in_sig & shiftedRoundMask; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  anyRoundExtra = |_anyRoundExtra_T; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  anyRound = roundPosBit | anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _roundIncr_T = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _roundIncr_T_1 = (roundingMode_near_even | roundingMode_near_maxMag) & roundPosBit; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _roundIncr_T_2 = roundMagUp & anyRound; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  roundIncr = _roundIncr_T_1 | _roundIncr_T_2; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [55:0] _roundedSig_T = io_in_sig | roundMask; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [54:0] _roundedSig_T_2 = _roundedSig_T[55:2] + 54'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _roundedSig_T_4 = ~anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 174:30]
  wire [54:0] _roundedSig_T_7 = roundingMode_near_even & roundPosBit & _roundedSig_T_4 ? shiftedRoundMask_lo : 55'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [54:0] _roundedSig_T_8 = ~_roundedSig_T_7; // @[RoundAnyRawFNToRecFN.scala 173:21]
  wire [54:0] _roundedSig_T_9 = _roundedSig_T_2 & _roundedSig_T_8; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [55:0] _roundedSig_T_10 = ~roundMask; // @[RoundAnyRawFNToRecFN.scala 178:32]
  wire [55:0] _roundedSig_T_11 = io_in_sig & _roundedSig_T_10; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire [54:0] _roundedSig_T_15 = roundingMode_odd & anyRound ? roundPosMask[55:1] : 55'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [54:0] _GEN_7 = {{1'd0}, _roundedSig_T_11[55:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [54:0] _roundedSig_T_16 = _GEN_7 | _roundedSig_T_15; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [54:0] roundedSig = roundIncr ? _roundedSig_T_9 : _roundedSig_T_16; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _sRoundedExp_T_1 = {1'b0,$signed(roundedSig[54:53])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [12:0] _GEN_8 = {{10{_sRoundedExp_T_1[2]}},_sRoundedExp_T_1}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [13:0] sRoundedExp = $signed(io_in_sExp) + $signed(_GEN_8); // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [11:0] common_expOut = sRoundedExp[11:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [51:0] common_fractOut = roundedSig[51:0]; // @[RoundAnyRawFNToRecFN.scala 189:27]
  wire [3:0] _common_overflow_T = sRoundedExp[13:10]; // @[RoundAnyRawFNToRecFN.scala 194:30]
  wire  common_overflow = $signed(_common_overflow_T) >= 4'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50]
  wire  common_totalUnderflow = $signed(sRoundedExp) < 14'sh3ce; // @[RoundAnyRawFNToRecFN.scala 198:31]
  wire  unboundedRange_roundPosBit = io_in_sig[1]; // @[RoundAnyRawFNToRecFN.scala 201:61]
  wire  unboundedRange_anyRound = |io_in_sig[1:0]; // @[RoundAnyRawFNToRecFN.scala 203:70]
  wire  _unboundedRange_roundIncr_T_1 = _roundIncr_T & unboundedRange_roundPosBit; // @[RoundAnyRawFNToRecFN.scala 205:67]
  wire  _unboundedRange_roundIncr_T_2 = roundMagUp & unboundedRange_anyRound; // @[RoundAnyRawFNToRecFN.scala 207:29]
  wire  unboundedRange_roundIncr = _unboundedRange_roundIncr_T_1 | _unboundedRange_roundIncr_T_2; // @[RoundAnyRawFNToRecFN.scala 206:46]
  wire  roundCarry = roundedSig[53]; // @[RoundAnyRawFNToRecFN.scala 211:27]
  wire [1:0] _common_underflow_T = io_in_sExp[12:11]; // @[RoundAnyRawFNToRecFN.scala 218:48]
  wire  _common_underflow_T_6 = anyRound & $signed(_common_underflow_T) <= 2'sh0 & roundMask[2]; // @[RoundAnyRawFNToRecFN.scala 218:74]
  wire  _common_underflow_T_11 = ~roundMask[3]; // @[RoundAnyRawFNToRecFN.scala 221:34]
  wire  _common_underflow_T_12 = io_detectTininess & _common_underflow_T_11; // @[RoundAnyRawFNToRecFN.scala 220:77]
  wire  _common_underflow_T_13 = _common_underflow_T_12 & roundCarry; // @[RoundAnyRawFNToRecFN.scala 224:38]
  wire  _common_underflow_T_15 = _common_underflow_T_13 & roundPosBit & unboundedRange_roundIncr; // @[RoundAnyRawFNToRecFN.scala 225:60]
  wire  _common_underflow_T_16 = ~_common_underflow_T_15; // @[RoundAnyRawFNToRecFN.scala 220:27]
  wire  _common_underflow_T_17 = _common_underflow_T_6 & _common_underflow_T_16; // @[RoundAnyRawFNToRecFN.scala 219:76]
  wire  common_underflow = common_totalUnderflow | _common_underflow_T_17; // @[RoundAnyRawFNToRecFN.scala 215:40]
  wire  common_inexact = common_totalUnderflow | anyRound; // @[RoundAnyRawFNToRecFN.scala 228:49]
  wire  isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  notNaN_isSpecialInfOut = io_infiniteExc | io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 234:49]
  wire  commonCase = ~isNaNOut & ~notNaN_isSpecialInfOut & ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:61]
  wire  overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  wire  underflow = commonCase & common_underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  wire  inexact = overflow | commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:28]
  wire  overflow_roundMagUp = _roundIncr_T | roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  wire  pegMinNonzeroMagOut = commonCase & common_totalUnderflow & (roundMagUp | roundingMode_odd); // @[RoundAnyRawFNToRecFN.scala 243:45]
  wire  pegMaxFiniteMagOut = overflow & ~overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 244:39]
  wire  notNaN_isInfOut = notNaN_isSpecialInfOut | overflow & overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 246:32]
  wire  signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire [11:0] _expOut_T_1 = io_in_isZero | common_totalUnderflow ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [11:0] _expOut_T_2 = ~_expOut_T_1; // @[RoundAnyRawFNToRecFN.scala 251:14]
  wire [11:0] _expOut_T_3 = common_expOut & _expOut_T_2; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [11:0] _expOut_T_5 = pegMinNonzeroMagOut ? 12'hc31 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 255:18]
  wire [11:0] _expOut_T_6 = ~_expOut_T_5; // @[RoundAnyRawFNToRecFN.scala 255:14]
  wire [11:0] _expOut_T_7 = _expOut_T_3 & _expOut_T_6; // @[RoundAnyRawFNToRecFN.scala 254:17]
  wire [11:0] _expOut_T_8 = pegMaxFiniteMagOut ? 12'h400 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 259:18]
  wire [11:0] _expOut_T_9 = ~_expOut_T_8; // @[RoundAnyRawFNToRecFN.scala 259:14]
  wire [11:0] _expOut_T_10 = _expOut_T_7 & _expOut_T_9; // @[RoundAnyRawFNToRecFN.scala 258:17]
  wire [11:0] _expOut_T_11 = notNaN_isInfOut ? 12'h200 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [11:0] _expOut_T_12 = ~_expOut_T_11; // @[RoundAnyRawFNToRecFN.scala 263:14]
  wire [11:0] _expOut_T_13 = _expOut_T_10 & _expOut_T_12; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [11:0] _expOut_T_14 = pegMinNonzeroMagOut ? 12'h3ce : 12'h0; // @[RoundAnyRawFNToRecFN.scala 267:16]
  wire [11:0] _expOut_T_15 = _expOut_T_13 | _expOut_T_14; // @[RoundAnyRawFNToRecFN.scala 266:18]
  wire [11:0] _expOut_T_16 = pegMaxFiniteMagOut ? 12'hbff : 12'h0; // @[RoundAnyRawFNToRecFN.scala 271:16]
  wire [11:0] _expOut_T_17 = _expOut_T_15 | _expOut_T_16; // @[RoundAnyRawFNToRecFN.scala 270:15]
  wire [11:0] _expOut_T_18 = notNaN_isInfOut ? 12'hc00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [11:0] _expOut_T_19 = _expOut_T_17 | _expOut_T_18; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [11:0] _expOut_T_20 = isNaNOut ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [11:0] expOut = _expOut_T_19 | _expOut_T_20; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire [51:0] _fractOut_T_2 = isNaNOut ? 52'h8000000000000 : 52'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [51:0] _fractOut_T_3 = isNaNOut | io_in_isZero | common_totalUnderflow ? _fractOut_T_2 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [51:0] _fractOut_T_5 = pegMaxFiniteMagOut ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [51:0] fractOut = _fractOut_T_3 | _fractOut_T_5; // @[RoundAnyRawFNToRecFN.scala 281:11]
  wire [12:0] io_out_hi = {signOut,expOut}; // @[Cat.scala 30:58]
  wire [1:0] io_exceptionFlags_lo = {underflow,inexact}; // @[Cat.scala 30:58]
  wire [2:0] io_exceptionFlags_hi = {io_invalidExc,io_infiniteExc,overflow}; // @[Cat.scala 30:58]
  assign io_out = {io_out_hi,fractOut}; // @[Cat.scala 30:58]
  assign io_exceptionFlags = {io_exceptionFlags_hi,io_exceptionFlags_lo}; // @[Cat.scala 30:58]
endmodule
