module BranchDecode(
  input         clock,
  input         reset,
  input  [31:0] io_inst,
  input  [39:0] io_pc,
  output        io_out_is_ret,
  output        io_out_is_call,
  output [39:0] io_out_target,
  output [2:0]  io_out_cfi_type,
  output        io_out_sfb_offset_valid,
  output [5:0]  io_out_sfb_offset_bits,
  output        io_out_shadowable
);
  wire [31:0] _bit_T = io_inst & 32'h707f; // @[Decode.scala 14:65]
  wire  _bit_T_1 = _bit_T == 32'h63; // @[Decode.scala 14:121]
  wire  _bit_T_3 = _bit_T == 32'h1063; // @[Decode.scala 14:121]
  wire  _bit_T_5 = _bit_T == 32'h5063; // @[Decode.scala 14:121]
  wire  _bit_T_7 = _bit_T == 32'h7063; // @[Decode.scala 14:121]
  wire  _bit_T_9 = _bit_T == 32'h4063; // @[Decode.scala 14:121]
  wire  _bit_T_11 = _bit_T == 32'h6063; // @[Decode.scala 14:121]
  wire  bpd_csignals_0 = _bit_T_1 | _bit_T_3 | _bit_T_5 | _bit_T_7 | _bit_T_9 | _bit_T_11; // @[Decode.scala 15:30]
  wire [31:0] _bit_T_17 = io_inst & 32'h7f; // @[Decode.scala 14:65]
  wire  bpd_csignals_1 = _bit_T_17 == 32'h6f; // @[Decode.scala 14:121]
  wire  bpd_csignals_2 = _bit_T == 32'h67; // @[Decode.scala 14:121]
  wire [31:0] _bit_T_21 = io_inst & 32'hfc00707f; // @[Decode.scala 14:65]
  wire  _bit_T_22 = _bit_T_21 == 32'h1013; // @[Decode.scala 14:121]
  wire  _bit_T_24 = _bit_T_21 == 32'h5013; // @[Decode.scala 14:121]
  wire  _bit_T_26 = _bit_T_21 == 32'h40005013; // @[Decode.scala 14:121]
  wire  _bit_T_28 = _bit_T == 32'h1b; // @[Decode.scala 14:121]
  wire [31:0] _bit_T_29 = io_inst & 32'hfe00707f; // @[Decode.scala 14:65]
  wire  _bit_T_30 = _bit_T_29 == 32'h101b; // @[Decode.scala 14:121]
  wire  _bit_T_32 = _bit_T_29 == 32'h4000501b; // @[Decode.scala 14:121]
  wire  _bit_T_34 = _bit_T_29 == 32'h501b; // @[Decode.scala 14:121]
  wire  _bit_T_36 = _bit_T_29 == 32'h3b; // @[Decode.scala 14:121]
  wire  _bit_T_38 = _bit_T_29 == 32'h4000003b; // @[Decode.scala 14:121]
  wire  _bit_T_40 = _bit_T_29 == 32'h103b; // @[Decode.scala 14:121]
  wire  _bit_T_42 = _bit_T_29 == 32'h4000503b; // @[Decode.scala 14:121]
  wire  _bit_T_44 = _bit_T_29 == 32'h503b; // @[Decode.scala 14:121]
  wire  _bit_T_46 = _bit_T_17 == 32'h37; // @[Decode.scala 14:121]
  wire  _bit_T_48 = _bit_T == 32'h13; // @[Decode.scala 14:121]
  wire  _bit_T_50 = _bit_T == 32'h7013; // @[Decode.scala 14:121]
  wire  _bit_T_52 = _bit_T == 32'h6013; // @[Decode.scala 14:121]
  wire  _bit_T_54 = _bit_T == 32'h4013; // @[Decode.scala 14:121]
  wire  _bit_T_56 = _bit_T == 32'h2013; // @[Decode.scala 14:121]
  wire  _bit_T_58 = _bit_T == 32'h3013; // @[Decode.scala 14:121]
  wire  _bit_T_60 = _bit_T_29 == 32'h1033; // @[Decode.scala 14:121]
  wire  _bit_T_62 = _bit_T_29 == 32'h33; // @[Decode.scala 14:121]
  wire  _bit_T_64 = _bit_T_29 == 32'h40000033; // @[Decode.scala 14:121]
  wire  _bit_T_66 = _bit_T_29 == 32'h2033; // @[Decode.scala 14:121]
  wire  _bit_T_68 = _bit_T_29 == 32'h3033; // @[Decode.scala 14:121]
  wire  _bit_T_70 = _bit_T_29 == 32'h7033; // @[Decode.scala 14:121]
  wire  _bit_T_72 = _bit_T_29 == 32'h6033; // @[Decode.scala 14:121]
  wire  _bit_T_74 = _bit_T_29 == 32'h4033; // @[Decode.scala 14:121]
  wire  _bit_T_76 = _bit_T_29 == 32'h40005033; // @[Decode.scala 14:121]
  wire  _bit_T_78 = _bit_T_29 == 32'h5033; // @[Decode.scala 14:121]
  wire  bpd_csignals_3 = _bit_T_22 | _bit_T_24 | _bit_T_26 | _bit_T_28 | _bit_T_30 | _bit_T_32 | _bit_T_34 | _bit_T_36
     | _bit_T_38 | _bit_T_40 | _bit_T_42 | _bit_T_44 | _bit_T_46 | _bit_T_48 | _bit_T_50 | _bit_T_52 | _bit_T_54 |
    _bit_T_56 | _bit_T_58 | _bit_T_60 | _bit_T_62 | _bit_T_64 | _bit_T_66 | _bit_T_68 | _bit_T_70 | _bit_T_72 |
    _bit_T_74 | _bit_T_76 | _bit_T_78; // @[Decode.scala 15:30]
  wire [31:0] _T = io_inst & 32'h24; // @[Decode.scala 14:65]
  wire  bpd_csignals_4 = _T == 32'h20; // @[Decode.scala 14:121]
  wire [4:0] _T_7 = io_inst[19:15] & 5'h1b; // @[decode.scala 686:51]
  wire [19:0] hi_hi_hi = io_inst[31] ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12]
  wire  hi_hi_lo = io_inst[7]; // @[consts.scala 337:46]
  wire [5:0] hi_lo = io_inst[30:25]; // @[consts.scala 337:55]
  wire [3:0] lo_hi = io_inst[11:8]; // @[consts.scala 337:68]
  wire [31:0] _T_17 = {hi_hi_hi,hi_hi_lo,hi_lo,lo_hi,1'h0}; // @[consts.scala 338:27]
  wire [39:0] _GEN_0 = {{8{_T_17[31]}},_T_17}; // @[consts.scala 338:17]
  wire [39:0] _T_20 = $signed(io_pc) + $signed(_GEN_0); // @[consts.scala 338:17]
  wire [39:0] _T_23 = $signed(_T_20) & -40'sh2; // @[consts.scala 338:52]
  wire [11:0] hi_hi_hi_1 = io_inst[31] ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [7:0] hi_hi_lo_1 = io_inst[19:12]; // @[consts.scala 343:46]
  wire  hi_lo_1 = io_inst[20]; // @[consts.scala 343:59]
  wire [3:0] lo_hi_lo = io_inst[24:21]; // @[consts.scala 343:82]
  wire [31:0] _T_28 = {hi_hi_hi_1,hi_hi_lo_1,hi_lo_1,hi_lo,lo_hi_lo,1'h0}; // @[consts.scala 344:27]
  wire [39:0] _GEN_1 = {{8{_T_28[31]}},_T_28}; // @[consts.scala 344:17]
  wire [39:0] _T_31 = $signed(io_pc) + $signed(_GEN_1); // @[consts.scala 344:17]
  wire [39:0] _T_34 = $signed(_T_31) & -40'sh2; // @[consts.scala 344:52]
  wire [2:0] _T_36 = bpd_csignals_0 ? 3'h1 : 3'h0; // @[decode.scala 695:8]
  wire [2:0] _T_37 = bpd_csignals_1 ? 3'h2 : _T_36; // @[decode.scala 693:8]
  wire [11:0] br_offset = {hi_hi_lo,hi_lo,lo_hi,1'h0}; // @[Cat.scala 30:58]
  wire  _T_50 = io_inst[19:15] == io_inst[11:7]; // @[decode.scala 705:22]
  wire  _T_51 = ~bpd_csignals_4 | _T_50; // @[decode.scala 704:17]
  wire  _T_56 = 32'h33 == _bit_T_29 & io_inst[19:15] == 5'h0; // @[decode.scala 706:22]
  wire  _T_57 = _T_51 | _T_56; // @[decode.scala 705:42]
  assign io_out_is_ret = bpd_csignals_2 & 5'h1 == _T_7 & io_inst[11:7] == 5'h0; // @[decode.scala 686:72]
  assign io_out_is_call = (bpd_csignals_1 | bpd_csignals_2) & io_inst[11:7] == 5'h1; // @[decode.scala 685:47]
  assign io_out_target = bpd_csignals_0 ? _T_23 : _T_34; // @[decode.scala 688:23]
  assign io_out_cfi_type = bpd_csignals_2 ? 3'h3 : _T_37; // @[decode.scala 691:8]
  assign io_out_sfb_offset_valid = bpd_csignals_0 & ~io_inst[31] & br_offset != 12'h0 & br_offset[11:6] == 6'h0; // @[decode.scala 701:76]
  assign io_out_sfb_offset_bits = br_offset[5:0]; // @[decode.scala 702:27]
  assign io_out_shadowable = bpd_csignals_3 & _T_57; // @[decode.scala 703:41]
endmodule
