module TLXbar_8(
  input   clock,
  input   reset
);
endmodule
