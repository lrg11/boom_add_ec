module BranchDecode(
  input         clock,
  input         reset,
  input  [31:0] io_inst,
  input  [39:0] io_pc,
  input         io_is_unicore,
  output        io_out_is_ret,
  output        io_out_is_call,
  output [39:0] io_out_target,
  output [2:0]  io_out_cfi_type,
  output        io_out_sfb_offset_valid,
  output [5:0]  io_out_sfb_offset_bits,
  output        io_out_shadowable
);
  wire [31:0] _bit_T = io_inst & 32'h707f; // @[Decode.scala 14:65]
  wire  _bit_T_1 = _bit_T == 32'h63; // @[Decode.scala 14:121]
  wire  _bit_T_3 = _bit_T == 32'h1063; // @[Decode.scala 14:121]
  wire  _bit_T_5 = _bit_T == 32'h5063; // @[Decode.scala 14:121]
  wire  _bit_T_7 = _bit_T == 32'h7063; // @[Decode.scala 14:121]
  wire  _bit_T_9 = _bit_T == 32'h4063; // @[Decode.scala 14:121]
  wire  _bit_T_11 = _bit_T == 32'h6063; // @[Decode.scala 14:121]
  wire  bpd_csignals_0 = _bit_T_1 | _bit_T_3 | _bit_T_5 | _bit_T_7 | _bit_T_9 | _bit_T_11; // @[Decode.scala 15:30]
  wire [31:0] _bit_T_17 = io_inst & 32'h7f; // @[Decode.scala 14:65]
  wire  bpd_csignals_1 = _bit_T_17 == 32'h6f; // @[Decode.scala 14:121]
  wire  bpd_csignals_2 = _bit_T == 32'h67; // @[Decode.scala 14:121]
  wire [31:0] _bit_T_21 = io_inst & 32'hfc00707f; // @[Decode.scala 14:65]
  wire  _bit_T_22 = _bit_T_21 == 32'h1013; // @[Decode.scala 14:121]
  wire  _bit_T_24 = _bit_T_21 == 32'h5013; // @[Decode.scala 14:121]
  wire  _bit_T_26 = _bit_T_21 == 32'h40005013; // @[Decode.scala 14:121]
  wire  _bit_T_28 = _bit_T == 32'h1b; // @[Decode.scala 14:121]
  wire [31:0] _bit_T_29 = io_inst & 32'hfe00707f; // @[Decode.scala 14:65]
  wire  _bit_T_30 = _bit_T_29 == 32'h101b; // @[Decode.scala 14:121]
  wire  _bit_T_32 = _bit_T_29 == 32'h4000501b; // @[Decode.scala 14:121]
  wire  _bit_T_34 = _bit_T_29 == 32'h501b; // @[Decode.scala 14:121]
  wire  _bit_T_36 = _bit_T_29 == 32'h3b; // @[Decode.scala 14:121]
  wire  _bit_T_38 = _bit_T_29 == 32'h4000003b; // @[Decode.scala 14:121]
  wire  _bit_T_40 = _bit_T_29 == 32'h103b; // @[Decode.scala 14:121]
  wire  _bit_T_42 = _bit_T_29 == 32'h4000503b; // @[Decode.scala 14:121]
  wire  _bit_T_44 = _bit_T_29 == 32'h503b; // @[Decode.scala 14:121]
  wire  _bit_T_46 = _bit_T_17 == 32'h37; // @[Decode.scala 14:121]
  wire  _bit_T_48 = _bit_T == 32'h13; // @[Decode.scala 14:121]
  wire  _bit_T_50 = _bit_T == 32'h7013; // @[Decode.scala 14:121]
  wire  _bit_T_52 = _bit_T == 32'h6013; // @[Decode.scala 14:121]
  wire  _bit_T_54 = _bit_T == 32'h4013; // @[Decode.scala 14:121]
  wire  _bit_T_56 = _bit_T == 32'h2013; // @[Decode.scala 14:121]
  wire  _bit_T_58 = _bit_T == 32'h3013; // @[Decode.scala 14:121]
  wire  _bit_T_60 = _bit_T_29 == 32'h1033; // @[Decode.scala 14:121]
  wire  _bit_T_62 = _bit_T_29 == 32'h33; // @[Decode.scala 14:121]
  wire  _bit_T_64 = _bit_T_29 == 32'h40000033; // @[Decode.scala 14:121]
  wire  _bit_T_66 = _bit_T_29 == 32'h2033; // @[Decode.scala 14:121]
  wire  _bit_T_68 = _bit_T_29 == 32'h3033; // @[Decode.scala 14:121]
  wire  _bit_T_70 = _bit_T_29 == 32'h7033; // @[Decode.scala 14:121]
  wire  _bit_T_72 = _bit_T_29 == 32'h6033; // @[Decode.scala 14:121]
  wire  _bit_T_74 = _bit_T_29 == 32'h4033; // @[Decode.scala 14:121]
  wire  _bit_T_76 = _bit_T_29 == 32'h40005033; // @[Decode.scala 14:121]
  wire  _bit_T_78 = _bit_T_29 == 32'h5033; // @[Decode.scala 14:121]
  wire  bpd_csignals_3 = _bit_T_22 | _bit_T_24 | _bit_T_26 | _bit_T_28 | _bit_T_30 | _bit_T_32 | _bit_T_34 | _bit_T_36
     | _bit_T_38 | _bit_T_40 | _bit_T_42 | _bit_T_44 | _bit_T_46 | _bit_T_48 | _bit_T_50 | _bit_T_52 | _bit_T_54 |
    _bit_T_56 | _bit_T_58 | _bit_T_60 | _bit_T_62 | _bit_T_64 | _bit_T_66 | _bit_T_68 | _bit_T_70 | _bit_T_72 |
    _bit_T_74 | _bit_T_76 | _bit_T_78; // @[Decode.scala 15:30]
  wire [31:0] _T = io_inst & 32'h24; // @[Decode.scala 14:65]
  wire  bpd_csignals_4 = _T == 32'h20; // @[Decode.scala 14:121]
  wire [31:0] _bit_T_107 = io_inst & 32'he9000000; // @[Decode.scala 14:65]
  wire  _bit_T_108 = _bit_T_107 == 32'ha0000000; // @[Decode.scala 14:121]
  wire [31:0] _bit_T_109 = io_inst & 32'hfd000000; // @[Decode.scala 14:65]
  wire  _bit_T_110 = _bit_T_109 == 32'hb8000000; // @[Decode.scala 14:121]
  wire  _bit_T_112 = _bit_T_107 == 32'ha1000000; // @[Decode.scala 14:121]
  wire  _bit_T_114 = _bit_T_109 == 32'hb9000000; // @[Decode.scala 14:121]
  wire  bpd_csignals_unicore_0 = _bit_T_108 | _bit_T_110 | _bit_T_112 | _bit_T_114; // @[Decode.scala 15:30]
  wire [31:0] _bit_T_118 = io_inst & 32'hff000000; // @[Decode.scala 14:65]
  wire  _bit_T_119 = _bit_T_118 == 32'hbc000000; // @[Decode.scala 14:121]
  wire  _bit_T_121 = _bit_T_118 == 32'hbd000000; // @[Decode.scala 14:121]
  wire  bpd_csignals_unicore_1 = _bit_T_119 | _bit_T_121; // @[Decode.scala 15:30]
  wire [31:0] _bit_T_123 = io_inst & 32'hffffffe0; // @[Decode.scala 14:65]
  wire  _bit_T_124 = _bit_T_123 == 32'h10ffc120; // @[Decode.scala 14:121]
  wire  _bit_T_126 = _bit_T_123 == 32'h11ffc120; // @[Decode.scala 14:121]
  wire  bpd_csignals_unicore_2 = _bit_T_124 | _bit_T_126; // @[Decode.scala 15:30]
  wire  cs_is_br = io_is_unicore ? bpd_csignals_unicore_0 : bpd_csignals_0; // @[decode.scala 956:24]
  wire  cs_is_jal = io_is_unicore ? bpd_csignals_unicore_1 : bpd_csignals_1; // @[decode.scala 957:24]
  wire  cs_is_jalr = io_is_unicore ? bpd_csignals_unicore_2 : bpd_csignals_2; // @[decode.scala 958:24]
  wire  is_call_riscv = (cs_is_jal | cs_is_jalr) & io_inst[11:7] == 5'h1; // @[decode.scala 959:49]
  wire [4:0] _T_6 = io_inst[19:15] & 5'h1b; // @[decode.scala 960:52]
  wire  is_ret_riscv = cs_is_jalr & 5'h1 == _T_6 & io_inst[11:7] == 5'h0; // @[decode.scala 960:73]
  wire [19:0] hi_hi_hi = io_inst[31] ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12]
  wire  hi_hi_lo = io_inst[7]; // @[consts.scala 470:46]
  wire [5:0] hi_lo = io_inst[30:25]; // @[consts.scala 470:55]
  wire [3:0] lo_hi = io_inst[11:8]; // @[consts.scala 470:68]
  wire [31:0] _T_15 = {hi_hi_hi,hi_hi_lo,hi_lo,lo_hi,1'h0}; // @[consts.scala 471:27]
  wire [39:0] _GEN_0 = {{8{_T_15[31]}},_T_15}; // @[consts.scala 471:17]
  wire [39:0] _T_18 = $signed(io_pc) + $signed(_GEN_0); // @[consts.scala 471:17]
  wire [39:0] _T_21 = $signed(_T_18) & -40'sh2; // @[consts.scala 471:52]
  wire [11:0] hi_hi_hi_1 = io_inst[31] ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [7:0] hi_hi_lo_1 = io_inst[19:12]; // @[consts.scala 476:46]
  wire  hi_lo_1 = io_inst[20]; // @[consts.scala 476:59]
  wire [3:0] lo_hi_lo = io_inst[24:21]; // @[consts.scala 476:82]
  wire [31:0] _T_26 = {hi_hi_hi_1,hi_hi_lo_1,hi_lo_1,hi_lo,lo_hi_lo,1'h0}; // @[consts.scala 477:27]
  wire [39:0] _GEN_1 = {{8{_T_26[31]}},_T_26}; // @[consts.scala 477:17]
  wire [39:0] _T_29 = $signed(io_pc) + $signed(_GEN_1); // @[consts.scala 477:17]
  wire [39:0] _T_32 = $signed(_T_29) & -40'sh2; // @[consts.scala 477:52]
  wire [39:0] target_riscv = cs_is_br ? _T_21 : _T_32; // @[decode.scala 961:25]
  wire [5:0] hi_hi_2 = io_inst[23] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [23:0] hi_lo_2 = io_inst[23:0]; // @[consts.scala 464:45]
  wire [31:0] _T_37 = {hi_hi_2,hi_lo_2,2'h0}; // @[consts.scala 465:27]
  wire [39:0] _GEN_2 = {{8{_T_37[31]}},_T_37}; // @[consts.scala 465:17]
  wire [39:0] _T_40 = $signed(io_pc) + $signed(_GEN_2); // @[consts.scala 465:17]
  wire [39:0] _T_43 = $signed(_T_40) + 40'sh4; // @[consts.scala 465:34]
  wire [39:0] target_unicore = $signed(_T_43) & -40'sh2; // @[consts.scala 465:51]
  wire [2:0] _T_49 = cs_is_br ? 3'h1 : 3'h0; // @[decode.scala 968:75]
  wire [2:0] _T_50 = cs_is_jal ? 3'h2 : _T_49; // @[decode.scala 968:51]
  wire [11:0] br_offset = {hi_hi_lo,hi_lo,lo_hi,1'h0}; // @[Cat.scala 30:58]
  wire  sfb_offset_valid_riscv = cs_is_br & ~io_inst[31] & br_offset != 12'h0 & br_offset[11:6] == 6'h0; // @[decode.scala 971:78]
  wire  _T_68 = 32'h33 == _bit_T_29 & io_inst[19:15] == 5'h0; // @[decode.scala 974:24]
  wire  _T_69 = ~bpd_csignals_4 | io_inst[19:15] == io_inst[11:7] | _T_68; // @[decode.scala 973:59]
  wire  shadowable_riscv = bpd_csignals_3 & _T_69; // @[decode.scala 972:43]
  assign io_out_is_ret = io_is_unicore ? 1'h0 : is_ret_riscv; // @[decode.scala 966:24]
  assign io_out_is_call = io_is_unicore ? 1'h0 : is_call_riscv; // @[decode.scala 965:24]
  assign io_out_target = io_is_unicore ? target_unicore : target_riscv; // @[decode.scala 967:23]
  assign io_out_cfi_type = cs_is_jalr ? 3'h3 : _T_50; // @[decode.scala 968:25]
  assign io_out_sfb_offset_valid = io_is_unicore ? 1'h0 : sfb_offset_valid_riscv; // @[decode.scala 976:33]
  assign io_out_sfb_offset_bits = br_offset[5:0]; // @[decode.scala 977:27]
  assign io_out_shadowable = io_is_unicore ? 1'h0 : shadowable_riscv; // @[decode.scala 978:27]
endmodule
