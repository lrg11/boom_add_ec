module BundleBridgeNexus_11(
  input   clock,
  input   reset,
  output  auto_out_enable,
  output  auto_out_stall
);
  assign auto_out_enable = 1'h0; // @[BaseTile.scala 271:19 BaseTile.scala 273:16]
  assign auto_out_stall = 1'h0; // @[BaseTile.scala 271:19 BaseTile.scala 272:16]
endmodule
