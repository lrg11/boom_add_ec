module BoomTile(
  input         clock,
  input         reset,
  output        auto_trace_out_0_valid,
  output [39:0] auto_trace_out_0_iaddr,
  output [31:0] auto_trace_out_0_insn,
  output [2:0]  auto_trace_out_0_priv,
  output        auto_trace_out_0_exception,
  output        auto_trace_out_0_interrupt,
  output [63:0] auto_trace_out_0_cause,
  output [39:0] auto_trace_out_0_tval,
  output [63:0] auto_trace_out_0_wdata,
  output        auto_trace_out_1_valid,
  output [39:0] auto_trace_out_1_iaddr,
  output [31:0] auto_trace_out_1_insn,
  output [2:0]  auto_trace_out_1_priv,
  output        auto_trace_out_1_exception,
  output        auto_trace_out_1_interrupt,
  output [63:0] auto_trace_out_1_cause,
  output [39:0] auto_trace_out_1_tval,
  output [63:0] auto_trace_out_1_wdata,
  output        auto_broadcast_out_0_valid,
  output [39:0] auto_broadcast_out_0_iaddr,
  output [31:0] auto_broadcast_out_0_insn,
  output [2:0]  auto_broadcast_out_0_priv,
  output        auto_broadcast_out_0_exception,
  output        auto_broadcast_out_0_interrupt,
  output [63:0] auto_broadcast_out_0_cause,
  output [39:0] auto_broadcast_out_0_tval,
  output        auto_broadcast_out_1_valid,
  output [39:0] auto_broadcast_out_1_iaddr,
  output [31:0] auto_broadcast_out_1_insn,
  output [2:0]  auto_broadcast_out_1_priv,
  output        auto_broadcast_out_1_exception,
  output        auto_broadcast_out_1_interrupt,
  output [63:0] auto_broadcast_out_1_cause,
  output [39:0] auto_broadcast_out_1_tval,
  output        auto_wfi_out_0,
  output        auto_cease_out_0,
  output        auto_halt_out_0,
  input         auto_int_local_in_3_0,
  input         auto_int_local_in_2_0,
  input         auto_int_local_in_1_0,
  input         auto_int_local_in_1_1,
  input         auto_int_local_in_0_0,
  output        auto_trace_core_source_out_group_0_iretire,
  output [31:0] auto_trace_core_source_out_group_0_iaddr,
  output [3:0]  auto_trace_core_source_out_group_0_itype,
  output        auto_trace_core_source_out_group_0_ilastsize,
  output [3:0]  auto_trace_core_source_out_priv,
  output [31:0] auto_trace_core_source_out_tval,
  output [31:0] auto_trace_core_source_out_cause,
  input         auto_nmi_in_rnmi,
  input  [31:0] auto_nmi_in_rnmi_interrupt_vector,
  input  [31:0] auto_nmi_in_rnmi_exception_vector,
  input         auto_nmi_in_unmi,
  input  [31:0] auto_nmi_in_unmi_interrupt_vector,
  input  [31:0] auto_nmi_in_unmi_exception_vector,
  input  [31:0] auto_reset_vector_in,
  input         auto_hartid_in,
  input         auto_tl_other_masters_out_a_ready,
  output        auto_tl_other_masters_out_a_valid,
  output [2:0]  auto_tl_other_masters_out_a_bits_opcode,
  output [2:0]  auto_tl_other_masters_out_a_bits_param,
  output [3:0]  auto_tl_other_masters_out_a_bits_size,
  output [2:0]  auto_tl_other_masters_out_a_bits_source,
  output [31:0] auto_tl_other_masters_out_a_bits_address,
  output [7:0]  auto_tl_other_masters_out_a_bits_mask,
  output [63:0] auto_tl_other_masters_out_a_bits_data,
  output        auto_tl_other_masters_out_a_bits_corrupt,
  output        auto_tl_other_masters_out_b_ready,
  input         auto_tl_other_masters_out_b_valid,
  input  [2:0]  auto_tl_other_masters_out_b_bits_opcode,
  input  [1:0]  auto_tl_other_masters_out_b_bits_param,
  input  [3:0]  auto_tl_other_masters_out_b_bits_size,
  input  [2:0]  auto_tl_other_masters_out_b_bits_source,
  input  [31:0] auto_tl_other_masters_out_b_bits_address,
  input  [7:0]  auto_tl_other_masters_out_b_bits_mask,
  input  [63:0] auto_tl_other_masters_out_b_bits_data,
  input         auto_tl_other_masters_out_b_bits_corrupt,
  input         auto_tl_other_masters_out_c_ready,
  output        auto_tl_other_masters_out_c_valid,
  output [2:0]  auto_tl_other_masters_out_c_bits_opcode,
  output [2:0]  auto_tl_other_masters_out_c_bits_param,
  output [3:0]  auto_tl_other_masters_out_c_bits_size,
  output [2:0]  auto_tl_other_masters_out_c_bits_source,
  output [31:0] auto_tl_other_masters_out_c_bits_address,
  output [63:0] auto_tl_other_masters_out_c_bits_data,
  output        auto_tl_other_masters_out_c_bits_corrupt,
  output        auto_tl_other_masters_out_d_ready,
  input         auto_tl_other_masters_out_d_valid,
  input  [2:0]  auto_tl_other_masters_out_d_bits_opcode,
  input  [1:0]  auto_tl_other_masters_out_d_bits_param,
  input  [3:0]  auto_tl_other_masters_out_d_bits_size,
  input  [2:0]  auto_tl_other_masters_out_d_bits_source,
  input  [1:0]  auto_tl_other_masters_out_d_bits_sink,
  input         auto_tl_other_masters_out_d_bits_denied,
  input  [63:0] auto_tl_other_masters_out_d_bits_data,
  input         auto_tl_other_masters_out_d_bits_corrupt,
  input         auto_tl_other_masters_out_e_ready,
  output        auto_tl_other_masters_out_e_valid,
  output [1:0]  auto_tl_other_masters_out_e_bits_sink
);
  wire  tlMasterXbar_clock; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_reset; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_1_a_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_1_a_valid; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_in_1_a_bits_opcode; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_in_1_a_bits_param; // @[BaseTile.scala 195:42]
  wire [3:0] tlMasterXbar_auto_in_1_a_bits_size; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_1_a_bits_source; // @[BaseTile.scala 195:42]
  wire [31:0] tlMasterXbar_auto_in_1_a_bits_address; // @[BaseTile.scala 195:42]
  wire [7:0] tlMasterXbar_auto_in_1_a_bits_mask; // @[BaseTile.scala 195:42]
  wire [63:0] tlMasterXbar_auto_in_1_a_bits_data; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_1_a_bits_corrupt; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_1_d_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_1_d_valid; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_in_1_d_bits_opcode; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_in_1_d_bits_param; // @[BaseTile.scala 195:42]
  wire [3:0] tlMasterXbar_auto_in_1_d_bits_size; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_1_d_bits_source; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_in_1_d_bits_sink; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_1_d_bits_denied; // @[BaseTile.scala 195:42]
  wire [63:0] tlMasterXbar_auto_in_1_d_bits_data; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_1_d_bits_corrupt; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_a_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_a_valid; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_in_0_a_bits_opcode; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_in_0_a_bits_param; // @[BaseTile.scala 195:42]
  wire [3:0] tlMasterXbar_auto_in_0_a_bits_size; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_in_0_a_bits_source; // @[BaseTile.scala 195:42]
  wire [31:0] tlMasterXbar_auto_in_0_a_bits_address; // @[BaseTile.scala 195:42]
  wire [7:0] tlMasterXbar_auto_in_0_a_bits_mask; // @[BaseTile.scala 195:42]
  wire [63:0] tlMasterXbar_auto_in_0_a_bits_data; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_a_bits_corrupt; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_b_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_b_valid; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_in_0_b_bits_opcode; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_in_0_b_bits_param; // @[BaseTile.scala 195:42]
  wire [3:0] tlMasterXbar_auto_in_0_b_bits_size; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_in_0_b_bits_source; // @[BaseTile.scala 195:42]
  wire [31:0] tlMasterXbar_auto_in_0_b_bits_address; // @[BaseTile.scala 195:42]
  wire [7:0] tlMasterXbar_auto_in_0_b_bits_mask; // @[BaseTile.scala 195:42]
  wire [63:0] tlMasterXbar_auto_in_0_b_bits_data; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_b_bits_corrupt; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_c_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_c_valid; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_in_0_c_bits_opcode; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_in_0_c_bits_param; // @[BaseTile.scala 195:42]
  wire [3:0] tlMasterXbar_auto_in_0_c_bits_size; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_in_0_c_bits_source; // @[BaseTile.scala 195:42]
  wire [31:0] tlMasterXbar_auto_in_0_c_bits_address; // @[BaseTile.scala 195:42]
  wire [63:0] tlMasterXbar_auto_in_0_c_bits_data; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_c_bits_corrupt; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_d_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_d_valid; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_in_0_d_bits_opcode; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_in_0_d_bits_param; // @[BaseTile.scala 195:42]
  wire [3:0] tlMasterXbar_auto_in_0_d_bits_size; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_in_0_d_bits_source; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_in_0_d_bits_sink; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_d_bits_denied; // @[BaseTile.scala 195:42]
  wire [63:0] tlMasterXbar_auto_in_0_d_bits_data; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_d_bits_corrupt; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_e_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_e_valid; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_in_0_e_bits_sink; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_a_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_a_valid; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_out_a_bits_opcode; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_out_a_bits_param; // @[BaseTile.scala 195:42]
  wire [3:0] tlMasterXbar_auto_out_a_bits_size; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_out_a_bits_source; // @[BaseTile.scala 195:42]
  wire [31:0] tlMasterXbar_auto_out_a_bits_address; // @[BaseTile.scala 195:42]
  wire [7:0] tlMasterXbar_auto_out_a_bits_mask; // @[BaseTile.scala 195:42]
  wire [63:0] tlMasterXbar_auto_out_a_bits_data; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_a_bits_corrupt; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_b_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_b_valid; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_out_b_bits_opcode; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_out_b_bits_param; // @[BaseTile.scala 195:42]
  wire [3:0] tlMasterXbar_auto_out_b_bits_size; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_out_b_bits_source; // @[BaseTile.scala 195:42]
  wire [31:0] tlMasterXbar_auto_out_b_bits_address; // @[BaseTile.scala 195:42]
  wire [7:0] tlMasterXbar_auto_out_b_bits_mask; // @[BaseTile.scala 195:42]
  wire [63:0] tlMasterXbar_auto_out_b_bits_data; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_b_bits_corrupt; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_c_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_c_valid; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_out_c_bits_opcode; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_out_c_bits_param; // @[BaseTile.scala 195:42]
  wire [3:0] tlMasterXbar_auto_out_c_bits_size; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_out_c_bits_source; // @[BaseTile.scala 195:42]
  wire [31:0] tlMasterXbar_auto_out_c_bits_address; // @[BaseTile.scala 195:42]
  wire [63:0] tlMasterXbar_auto_out_c_bits_data; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_c_bits_corrupt; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_d_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_d_valid; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_out_d_bits_opcode; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_out_d_bits_param; // @[BaseTile.scala 195:42]
  wire [3:0] tlMasterXbar_auto_out_d_bits_size; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_out_d_bits_source; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_out_d_bits_sink; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_d_bits_denied; // @[BaseTile.scala 195:42]
  wire [63:0] tlMasterXbar_auto_out_d_bits_data; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_d_bits_corrupt; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_e_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_e_valid; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_out_e_bits_sink; // @[BaseTile.scala 195:42]
  wire  tlSlaveXbar_clock; // @[BaseTile.scala 196:41]
  wire  tlSlaveXbar_reset; // @[BaseTile.scala 196:41]
  wire  intXbar_clock; // @[BaseTile.scala 197:37]
  wire  intXbar_reset; // @[BaseTile.scala 197:37]
  wire  intXbar_auto_int_in_3_0; // @[BaseTile.scala 197:37]
  wire  intXbar_auto_int_in_2_0; // @[BaseTile.scala 197:37]
  wire  intXbar_auto_int_in_1_0; // @[BaseTile.scala 197:37]
  wire  intXbar_auto_int_in_1_1; // @[BaseTile.scala 197:37]
  wire  intXbar_auto_int_in_0_0; // @[BaseTile.scala 197:37]
  wire  intXbar_auto_int_out_0; // @[BaseTile.scala 197:37]
  wire  intXbar_auto_int_out_1; // @[BaseTile.scala 197:37]
  wire  intXbar_auto_int_out_2; // @[BaseTile.scala 197:37]
  wire  intXbar_auto_int_out_3; // @[BaseTile.scala 197:37]
  wire  intXbar_auto_int_out_4; // @[BaseTile.scala 197:37]
  wire  broadcast_clock; // @[BundleBridge.scala 196:31]
  wire  broadcast_reset; // @[BundleBridge.scala 196:31]
  wire  broadcast_auto_in; // @[BundleBridge.scala 196:31]
  wire  broadcast_auto_out; // @[BundleBridge.scala 196:31]
  wire  broadcast_1_clock; // @[BundleBridge.scala 196:31]
  wire  broadcast_1_reset; // @[BundleBridge.scala 196:31]
  wire [31:0] broadcast_1_auto_in; // @[BundleBridge.scala 196:31]
  wire [31:0] broadcast_1_auto_out_1; // @[BundleBridge.scala 196:31]
  wire [31:0] broadcast_1_auto_out_0; // @[BundleBridge.scala 196:31]
  wire  broadcast_2_clock; // @[BundleBridge.scala 196:31]
  wire  broadcast_2_reset; // @[BundleBridge.scala 196:31]
  wire  broadcast_2_auto_in_rnmi; // @[BundleBridge.scala 196:31]
  wire [31:0] broadcast_2_auto_in_rnmi_interrupt_vector; // @[BundleBridge.scala 196:31]
  wire [31:0] broadcast_2_auto_in_rnmi_exception_vector; // @[BundleBridge.scala 196:31]
  wire  broadcast_2_auto_in_unmi; // @[BundleBridge.scala 196:31]
  wire [31:0] broadcast_2_auto_in_unmi_interrupt_vector; // @[BundleBridge.scala 196:31]
  wire [31:0] broadcast_2_auto_in_unmi_exception_vector; // @[BundleBridge.scala 196:31]
  wire  broadcast_2_auto_out_rnmi; // @[BundleBridge.scala 196:31]
  wire [31:0] broadcast_2_auto_out_rnmi_interrupt_vector; // @[BundleBridge.scala 196:31]
  wire [31:0] broadcast_2_auto_out_rnmi_exception_vector; // @[BundleBridge.scala 196:31]
  wire  broadcast_2_auto_out_unmi; // @[BundleBridge.scala 196:31]
  wire [31:0] broadcast_2_auto_out_unmi_interrupt_vector; // @[BundleBridge.scala 196:31]
  wire [31:0] broadcast_2_auto_out_unmi_exception_vector; // @[BundleBridge.scala 196:31]
  wire  nexus_clock; // @[BundleBridge.scala 183:27]
  wire  nexus_reset; // @[BundleBridge.scala 183:27]
  wire  broadcast_3_clock; // @[BundleBridge.scala 196:31]
  wire  broadcast_3_reset; // @[BundleBridge.scala 196:31]
  wire  broadcast_3_auto_in_0_valid; // @[BundleBridge.scala 196:31]
  wire [39:0] broadcast_3_auto_in_0_iaddr; // @[BundleBridge.scala 196:31]
  wire [31:0] broadcast_3_auto_in_0_insn; // @[BundleBridge.scala 196:31]
  wire [2:0] broadcast_3_auto_in_0_priv; // @[BundleBridge.scala 196:31]
  wire  broadcast_3_auto_in_0_exception; // @[BundleBridge.scala 196:31]
  wire  broadcast_3_auto_in_0_interrupt; // @[BundleBridge.scala 196:31]
  wire [63:0] broadcast_3_auto_in_0_cause; // @[BundleBridge.scala 196:31]
  wire [39:0] broadcast_3_auto_in_0_tval; // @[BundleBridge.scala 196:31]
  wire  broadcast_3_auto_in_1_valid; // @[BundleBridge.scala 196:31]
  wire [39:0] broadcast_3_auto_in_1_iaddr; // @[BundleBridge.scala 196:31]
  wire [31:0] broadcast_3_auto_in_1_insn; // @[BundleBridge.scala 196:31]
  wire [2:0] broadcast_3_auto_in_1_priv; // @[BundleBridge.scala 196:31]
  wire  broadcast_3_auto_in_1_exception; // @[BundleBridge.scala 196:31]
  wire  broadcast_3_auto_in_1_interrupt; // @[BundleBridge.scala 196:31]
  wire [63:0] broadcast_3_auto_in_1_cause; // @[BundleBridge.scala 196:31]
  wire [39:0] broadcast_3_auto_in_1_tval; // @[BundleBridge.scala 196:31]
  wire  broadcast_3_auto_out_0_valid; // @[BundleBridge.scala 196:31]
  wire [39:0] broadcast_3_auto_out_0_iaddr; // @[BundleBridge.scala 196:31]
  wire [31:0] broadcast_3_auto_out_0_insn; // @[BundleBridge.scala 196:31]
  wire [2:0] broadcast_3_auto_out_0_priv; // @[BundleBridge.scala 196:31]
  wire  broadcast_3_auto_out_0_exception; // @[BundleBridge.scala 196:31]
  wire  broadcast_3_auto_out_0_interrupt; // @[BundleBridge.scala 196:31]
  wire [63:0] broadcast_3_auto_out_0_cause; // @[BundleBridge.scala 196:31]
  wire [39:0] broadcast_3_auto_out_0_tval; // @[BundleBridge.scala 196:31]
  wire  broadcast_3_auto_out_1_valid; // @[BundleBridge.scala 196:31]
  wire [39:0] broadcast_3_auto_out_1_iaddr; // @[BundleBridge.scala 196:31]
  wire [31:0] broadcast_3_auto_out_1_insn; // @[BundleBridge.scala 196:31]
  wire [2:0] broadcast_3_auto_out_1_priv; // @[BundleBridge.scala 196:31]
  wire  broadcast_3_auto_out_1_exception; // @[BundleBridge.scala 196:31]
  wire  broadcast_3_auto_out_1_interrupt; // @[BundleBridge.scala 196:31]
  wire [63:0] broadcast_3_auto_out_1_cause; // @[BundleBridge.scala 196:31]
  wire [39:0] broadcast_3_auto_out_1_tval; // @[BundleBridge.scala 196:31]
  wire  nexus_1_clock; // @[BundleBridge.scala 183:27]
  wire  nexus_1_reset; // @[BundleBridge.scala 183:27]
  wire  nexus_1_auto_out_enable; // @[BundleBridge.scala 183:27]
  wire  nexus_1_auto_out_stall; // @[BundleBridge.scala 183:27]
  wire  broadcast_4_clock; // @[BundleBridge.scala 196:31]
  wire  broadcast_4_reset; // @[BundleBridge.scala 196:31]
  wire  trace_clock; // @[BundleBridge.scala 196:31]
  wire  trace_reset; // @[BundleBridge.scala 196:31]
  wire  trace_auto_in_0_valid; // @[BundleBridge.scala 196:31]
  wire [39:0] trace_auto_in_0_iaddr; // @[BundleBridge.scala 196:31]
  wire [31:0] trace_auto_in_0_insn; // @[BundleBridge.scala 196:31]
  wire [2:0] trace_auto_in_0_priv; // @[BundleBridge.scala 196:31]
  wire  trace_auto_in_0_exception; // @[BundleBridge.scala 196:31]
  wire  trace_auto_in_0_interrupt; // @[BundleBridge.scala 196:31]
  wire [63:0] trace_auto_in_0_cause; // @[BundleBridge.scala 196:31]
  wire [39:0] trace_auto_in_0_tval; // @[BundleBridge.scala 196:31]
  wire [63:0] trace_auto_in_0_wdata; // @[BundleBridge.scala 196:31]
  wire  trace_auto_in_1_valid; // @[BundleBridge.scala 196:31]
  wire [39:0] trace_auto_in_1_iaddr; // @[BundleBridge.scala 196:31]
  wire [31:0] trace_auto_in_1_insn; // @[BundleBridge.scala 196:31]
  wire [2:0] trace_auto_in_1_priv; // @[BundleBridge.scala 196:31]
  wire  trace_auto_in_1_exception; // @[BundleBridge.scala 196:31]
  wire  trace_auto_in_1_interrupt; // @[BundleBridge.scala 196:31]
  wire [63:0] trace_auto_in_1_cause; // @[BundleBridge.scala 196:31]
  wire [39:0] trace_auto_in_1_tval; // @[BundleBridge.scala 196:31]
  wire [63:0] trace_auto_in_1_wdata; // @[BundleBridge.scala 196:31]
  wire  trace_auto_out_0_valid; // @[BundleBridge.scala 196:31]
  wire [39:0] trace_auto_out_0_iaddr; // @[BundleBridge.scala 196:31]
  wire [31:0] trace_auto_out_0_insn; // @[BundleBridge.scala 196:31]
  wire [2:0] trace_auto_out_0_priv; // @[BundleBridge.scala 196:31]
  wire  trace_auto_out_0_exception; // @[BundleBridge.scala 196:31]
  wire  trace_auto_out_0_interrupt; // @[BundleBridge.scala 196:31]
  wire [63:0] trace_auto_out_0_cause; // @[BundleBridge.scala 196:31]
  wire [39:0] trace_auto_out_0_tval; // @[BundleBridge.scala 196:31]
  wire [63:0] trace_auto_out_0_wdata; // @[BundleBridge.scala 196:31]
  wire  trace_auto_out_1_valid; // @[BundleBridge.scala 196:31]
  wire [39:0] trace_auto_out_1_iaddr; // @[BundleBridge.scala 196:31]
  wire [31:0] trace_auto_out_1_insn; // @[BundleBridge.scala 196:31]
  wire [2:0] trace_auto_out_1_priv; // @[BundleBridge.scala 196:31]
  wire  trace_auto_out_1_exception; // @[BundleBridge.scala 196:31]
  wire  trace_auto_out_1_interrupt; // @[BundleBridge.scala 196:31]
  wire [63:0] trace_auto_out_1_cause; // @[BundleBridge.scala 196:31]
  wire [39:0] trace_auto_out_1_tval; // @[BundleBridge.scala 196:31]
  wire [63:0] trace_auto_out_1_wdata; // @[BundleBridge.scala 196:31]
  wire  dcache_clock; // @[tile.scala 134:54]
  wire  dcache_reset; // @[tile.scala 134:54]
  wire  dcache_auto_out_a_ready; // @[tile.scala 134:54]
  wire  dcache_auto_out_a_valid; // @[tile.scala 134:54]
  wire [2:0] dcache_auto_out_a_bits_opcode; // @[tile.scala 134:54]
  wire [2:0] dcache_auto_out_a_bits_param; // @[tile.scala 134:54]
  wire [3:0] dcache_auto_out_a_bits_size; // @[tile.scala 134:54]
  wire [1:0] dcache_auto_out_a_bits_source; // @[tile.scala 134:54]
  wire [31:0] dcache_auto_out_a_bits_address; // @[tile.scala 134:54]
  wire [7:0] dcache_auto_out_a_bits_mask; // @[tile.scala 134:54]
  wire [63:0] dcache_auto_out_a_bits_data; // @[tile.scala 134:54]
  wire  dcache_auto_out_a_bits_corrupt; // @[tile.scala 134:54]
  wire  dcache_auto_out_b_ready; // @[tile.scala 134:54]
  wire  dcache_auto_out_b_valid; // @[tile.scala 134:54]
  wire [2:0] dcache_auto_out_b_bits_opcode; // @[tile.scala 134:54]
  wire [1:0] dcache_auto_out_b_bits_param; // @[tile.scala 134:54]
  wire [3:0] dcache_auto_out_b_bits_size; // @[tile.scala 134:54]
  wire [1:0] dcache_auto_out_b_bits_source; // @[tile.scala 134:54]
  wire [31:0] dcache_auto_out_b_bits_address; // @[tile.scala 134:54]
  wire [7:0] dcache_auto_out_b_bits_mask; // @[tile.scala 134:54]
  wire [63:0] dcache_auto_out_b_bits_data; // @[tile.scala 134:54]
  wire  dcache_auto_out_b_bits_corrupt; // @[tile.scala 134:54]
  wire  dcache_auto_out_c_ready; // @[tile.scala 134:54]
  wire  dcache_auto_out_c_valid; // @[tile.scala 134:54]
  wire [2:0] dcache_auto_out_c_bits_opcode; // @[tile.scala 134:54]
  wire [2:0] dcache_auto_out_c_bits_param; // @[tile.scala 134:54]
  wire [3:0] dcache_auto_out_c_bits_size; // @[tile.scala 134:54]
  wire [1:0] dcache_auto_out_c_bits_source; // @[tile.scala 134:54]
  wire [31:0] dcache_auto_out_c_bits_address; // @[tile.scala 134:54]
  wire [63:0] dcache_auto_out_c_bits_data; // @[tile.scala 134:54]
  wire  dcache_auto_out_c_bits_corrupt; // @[tile.scala 134:54]
  wire  dcache_auto_out_d_ready; // @[tile.scala 134:54]
  wire  dcache_auto_out_d_valid; // @[tile.scala 134:54]
  wire [2:0] dcache_auto_out_d_bits_opcode; // @[tile.scala 134:54]
  wire [1:0] dcache_auto_out_d_bits_param; // @[tile.scala 134:54]
  wire [3:0] dcache_auto_out_d_bits_size; // @[tile.scala 134:54]
  wire [1:0] dcache_auto_out_d_bits_source; // @[tile.scala 134:54]
  wire [1:0] dcache_auto_out_d_bits_sink; // @[tile.scala 134:54]
  wire  dcache_auto_out_d_bits_denied; // @[tile.scala 134:54]
  wire [63:0] dcache_auto_out_d_bits_data; // @[tile.scala 134:54]
  wire  dcache_auto_out_d_bits_corrupt; // @[tile.scala 134:54]
  wire  dcache_auto_out_e_ready; // @[tile.scala 134:54]
  wire  dcache_auto_out_e_valid; // @[tile.scala 134:54]
  wire [1:0] dcache_auto_out_e_bits_sink; // @[tile.scala 134:54]
  wire  dcache_io_errors_bus_valid; // @[tile.scala 134:54]
  wire [31:0] dcache_io_errors_bus_bits; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_ready; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_valid; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_valid; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_switch; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_switch_off; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_is_unicore; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_req_bits_0_bits_uop_shift; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_req_bits_0_bits_uop_lrs3_rtype; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_rflag; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_wflag; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_req_bits_0_bits_uop_prflag; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_req_bits_0_bits_uop_pwflag; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_pflag_busy; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_req_bits_0_bits_uop_stale_pflag; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_req_bits_0_bits_uop_op1_sel; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_req_bits_0_bits_uop_op2_sel; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_req_bits_0_bits_uop_split_num; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_req_bits_0_bits_uop_self_index; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_req_bits_0_bits_uop_rob_inst_idx; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_req_bits_0_bits_uop_address_num; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_req_bits_0_bits_uop_uopc; // @[tile.scala 134:54]
  wire [31:0] dcache_io_lsu_req_bits_0_bits_uop_inst; // @[tile.scala 134:54]
  wire [31:0] dcache_io_lsu_req_bits_0_bits_uop_debug_inst; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_is_rvc; // @[tile.scala 134:54]
  wire [39:0] dcache_io_lsu_req_bits_0_bits_uop_debug_pc; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_req_bits_0_bits_uop_iq_type; // @[tile.scala 134:54]
  wire [9:0] dcache_io_lsu_req_bits_0_bits_uop_fu_code; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_req_bits_0_bits_uop_ctrl_br_type; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_req_bits_0_bits_uop_ctrl_op1_sel; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_req_bits_0_bits_uop_ctrl_op2_sel; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_req_bits_0_bits_uop_ctrl_imm_sel; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_req_bits_0_bits_uop_ctrl_op_fcn; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_ctrl_fcn_dw; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_req_bits_0_bits_uop_ctrl_csr_cmd; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_ctrl_is_load; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_ctrl_is_sta; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_ctrl_is_std; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_req_bits_0_bits_uop_ctrl_op3_sel; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_req_bits_0_bits_uop_iw_state; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_iw_p1_poisoned; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_iw_p2_poisoned; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_is_br; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_is_jalr; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_is_jal; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_is_sfb; // @[tile.scala 134:54]
  wire [11:0] dcache_io_lsu_req_bits_0_bits_uop_br_mask; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_req_bits_0_bits_uop_br_tag; // @[tile.scala 134:54]
  wire [4:0] dcache_io_lsu_req_bits_0_bits_uop_ftq_idx; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_edge_inst; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_req_bits_0_bits_uop_pc_lob; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_taken; // @[tile.scala 134:54]
  wire [19:0] dcache_io_lsu_req_bits_0_bits_uop_imm_packed; // @[tile.scala 134:54]
  wire [11:0] dcache_io_lsu_req_bits_0_bits_uop_csr_addr; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_req_bits_0_bits_uop_rob_idx; // @[tile.scala 134:54]
  wire [4:0] dcache_io_lsu_req_bits_0_bits_uop_ldq_idx; // @[tile.scala 134:54]
  wire [4:0] dcache_io_lsu_req_bits_0_bits_uop_stq_idx; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_req_bits_0_bits_uop_rxq_idx; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_req_bits_0_bits_uop_pdst; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_req_bits_0_bits_uop_prs1; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_req_bits_0_bits_uop_prs2; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_req_bits_0_bits_uop_prs3; // @[tile.scala 134:54]
  wire [4:0] dcache_io_lsu_req_bits_0_bits_uop_ppred; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_prs1_busy; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_prs2_busy; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_prs3_busy; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_ppred_busy; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_req_bits_0_bits_uop_stale_pdst; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_exception; // @[tile.scala 134:54]
  wire [63:0] dcache_io_lsu_req_bits_0_bits_uop_exc_cause; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_bypassable; // @[tile.scala 134:54]
  wire [4:0] dcache_io_lsu_req_bits_0_bits_uop_mem_cmd; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_req_bits_0_bits_uop_mem_size; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_mem_signed; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_is_fence; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_is_fencei; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_is_amo; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_uses_ldq; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_uses_stq; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_is_sys_pc2epc; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_is_unique; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_flush_on_commit; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_ldst_is_rs1; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_req_bits_0_bits_uop_ldst; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_req_bits_0_bits_uop_lrs1; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_req_bits_0_bits_uop_lrs2; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_req_bits_0_bits_uop_lrs3; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_ldst_val; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_req_bits_0_bits_uop_dst_rtype; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_req_bits_0_bits_uop_lrs1_rtype; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_req_bits_0_bits_uop_lrs2_rtype; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_frs3_en; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_fp_val; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_fp_single; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_xcpt_pf_if; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_xcpt_ae_if; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_xcpt_ma_if; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_bp_debug_if; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_uop_bp_xcpt_if; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_req_bits_0_bits_uop_debug_fsrc; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_req_bits_0_bits_uop_debug_tsrc; // @[tile.scala 134:54]
  wire [39:0] dcache_io_lsu_req_bits_0_bits_addr; // @[tile.scala 134:54]
  wire [63:0] dcache_io_lsu_req_bits_0_bits_data; // @[tile.scala 134:54]
  wire  dcache_io_lsu_req_bits_0_bits_is_hella; // @[tile.scala 134:54]
  wire  dcache_io_lsu_s1_kill_0; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_valid; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_switch; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_switch_off; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_is_unicore; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_resp_0_bits_uop_shift; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_resp_0_bits_uop_lrs3_rtype; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_rflag; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_wflag; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_resp_0_bits_uop_prflag; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_resp_0_bits_uop_pwflag; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_pflag_busy; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_resp_0_bits_uop_stale_pflag; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_resp_0_bits_uop_op1_sel; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_resp_0_bits_uop_op2_sel; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_resp_0_bits_uop_split_num; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_resp_0_bits_uop_self_index; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_resp_0_bits_uop_rob_inst_idx; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_resp_0_bits_uop_address_num; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_resp_0_bits_uop_uopc; // @[tile.scala 134:54]
  wire [31:0] dcache_io_lsu_resp_0_bits_uop_inst; // @[tile.scala 134:54]
  wire [31:0] dcache_io_lsu_resp_0_bits_uop_debug_inst; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_is_rvc; // @[tile.scala 134:54]
  wire [39:0] dcache_io_lsu_resp_0_bits_uop_debug_pc; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_resp_0_bits_uop_iq_type; // @[tile.scala 134:54]
  wire [9:0] dcache_io_lsu_resp_0_bits_uop_fu_code; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_resp_0_bits_uop_ctrl_br_type; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_resp_0_bits_uop_ctrl_op1_sel; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_resp_0_bits_uop_ctrl_op2_sel; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_resp_0_bits_uop_ctrl_imm_sel; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_resp_0_bits_uop_ctrl_op_fcn; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_ctrl_fcn_dw; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_resp_0_bits_uop_ctrl_csr_cmd; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_ctrl_is_load; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_ctrl_is_sta; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_ctrl_is_std; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_resp_0_bits_uop_ctrl_op3_sel; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_resp_0_bits_uop_iw_state; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_iw_p1_poisoned; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_iw_p2_poisoned; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_is_br; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_is_jalr; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_is_jal; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_is_sfb; // @[tile.scala 134:54]
  wire [11:0] dcache_io_lsu_resp_0_bits_uop_br_mask; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_resp_0_bits_uop_br_tag; // @[tile.scala 134:54]
  wire [4:0] dcache_io_lsu_resp_0_bits_uop_ftq_idx; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_edge_inst; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_resp_0_bits_uop_pc_lob; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_taken; // @[tile.scala 134:54]
  wire [19:0] dcache_io_lsu_resp_0_bits_uop_imm_packed; // @[tile.scala 134:54]
  wire [11:0] dcache_io_lsu_resp_0_bits_uop_csr_addr; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_resp_0_bits_uop_rob_idx; // @[tile.scala 134:54]
  wire [4:0] dcache_io_lsu_resp_0_bits_uop_ldq_idx; // @[tile.scala 134:54]
  wire [4:0] dcache_io_lsu_resp_0_bits_uop_stq_idx; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_resp_0_bits_uop_rxq_idx; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_resp_0_bits_uop_pdst; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_resp_0_bits_uop_prs1; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_resp_0_bits_uop_prs2; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_resp_0_bits_uop_prs3; // @[tile.scala 134:54]
  wire [4:0] dcache_io_lsu_resp_0_bits_uop_ppred; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_prs1_busy; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_prs2_busy; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_prs3_busy; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_ppred_busy; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_resp_0_bits_uop_stale_pdst; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_exception; // @[tile.scala 134:54]
  wire [63:0] dcache_io_lsu_resp_0_bits_uop_exc_cause; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_bypassable; // @[tile.scala 134:54]
  wire [4:0] dcache_io_lsu_resp_0_bits_uop_mem_cmd; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_resp_0_bits_uop_mem_size; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_mem_signed; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_is_fence; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_is_fencei; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_is_amo; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_uses_ldq; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_uses_stq; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_is_sys_pc2epc; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_is_unique; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_flush_on_commit; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_ldst_is_rs1; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_resp_0_bits_uop_ldst; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_resp_0_bits_uop_lrs1; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_resp_0_bits_uop_lrs2; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_resp_0_bits_uop_lrs3; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_ldst_val; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_resp_0_bits_uop_dst_rtype; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_resp_0_bits_uop_lrs1_rtype; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_resp_0_bits_uop_lrs2_rtype; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_frs3_en; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_fp_val; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_fp_single; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_xcpt_pf_if; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_xcpt_ae_if; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_xcpt_ma_if; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_bp_debug_if; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_uop_bp_xcpt_if; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_resp_0_bits_uop_debug_fsrc; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_resp_0_bits_uop_debug_tsrc; // @[tile.scala 134:54]
  wire [63:0] dcache_io_lsu_resp_0_bits_data; // @[tile.scala 134:54]
  wire  dcache_io_lsu_resp_0_bits_is_hella; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_valid; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_switch; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_switch_off; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_is_unicore; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_nack_0_bits_uop_shift; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_nack_0_bits_uop_lrs3_rtype; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_rflag; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_wflag; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_nack_0_bits_uop_prflag; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_nack_0_bits_uop_pwflag; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_pflag_busy; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_nack_0_bits_uop_stale_pflag; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_nack_0_bits_uop_op1_sel; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_nack_0_bits_uop_op2_sel; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_nack_0_bits_uop_split_num; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_nack_0_bits_uop_self_index; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_nack_0_bits_uop_rob_inst_idx; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_nack_0_bits_uop_address_num; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_nack_0_bits_uop_uopc; // @[tile.scala 134:54]
  wire [31:0] dcache_io_lsu_nack_0_bits_uop_inst; // @[tile.scala 134:54]
  wire [31:0] dcache_io_lsu_nack_0_bits_uop_debug_inst; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_is_rvc; // @[tile.scala 134:54]
  wire [39:0] dcache_io_lsu_nack_0_bits_uop_debug_pc; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_nack_0_bits_uop_iq_type; // @[tile.scala 134:54]
  wire [9:0] dcache_io_lsu_nack_0_bits_uop_fu_code; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_nack_0_bits_uop_ctrl_br_type; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_nack_0_bits_uop_ctrl_op1_sel; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_nack_0_bits_uop_ctrl_op2_sel; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_nack_0_bits_uop_ctrl_imm_sel; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_nack_0_bits_uop_ctrl_op_fcn; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_ctrl_fcn_dw; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_nack_0_bits_uop_ctrl_csr_cmd; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_ctrl_is_load; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_ctrl_is_sta; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_ctrl_is_std; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_nack_0_bits_uop_ctrl_op3_sel; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_nack_0_bits_uop_iw_state; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_iw_p1_poisoned; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_iw_p2_poisoned; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_is_br; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_is_jalr; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_is_jal; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_is_sfb; // @[tile.scala 134:54]
  wire [11:0] dcache_io_lsu_nack_0_bits_uop_br_mask; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_nack_0_bits_uop_br_tag; // @[tile.scala 134:54]
  wire [4:0] dcache_io_lsu_nack_0_bits_uop_ftq_idx; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_edge_inst; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_nack_0_bits_uop_pc_lob; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_taken; // @[tile.scala 134:54]
  wire [19:0] dcache_io_lsu_nack_0_bits_uop_imm_packed; // @[tile.scala 134:54]
  wire [11:0] dcache_io_lsu_nack_0_bits_uop_csr_addr; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_nack_0_bits_uop_rob_idx; // @[tile.scala 134:54]
  wire [4:0] dcache_io_lsu_nack_0_bits_uop_ldq_idx; // @[tile.scala 134:54]
  wire [4:0] dcache_io_lsu_nack_0_bits_uop_stq_idx; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_nack_0_bits_uop_rxq_idx; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_nack_0_bits_uop_pdst; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_nack_0_bits_uop_prs1; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_nack_0_bits_uop_prs2; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_nack_0_bits_uop_prs3; // @[tile.scala 134:54]
  wire [4:0] dcache_io_lsu_nack_0_bits_uop_ppred; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_prs1_busy; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_prs2_busy; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_prs3_busy; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_ppred_busy; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_nack_0_bits_uop_stale_pdst; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_exception; // @[tile.scala 134:54]
  wire [63:0] dcache_io_lsu_nack_0_bits_uop_exc_cause; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_bypassable; // @[tile.scala 134:54]
  wire [4:0] dcache_io_lsu_nack_0_bits_uop_mem_cmd; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_nack_0_bits_uop_mem_size; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_mem_signed; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_is_fence; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_is_fencei; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_is_amo; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_uses_ldq; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_uses_stq; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_is_sys_pc2epc; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_is_unique; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_flush_on_commit; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_ldst_is_rs1; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_nack_0_bits_uop_ldst; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_nack_0_bits_uop_lrs1; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_nack_0_bits_uop_lrs2; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_nack_0_bits_uop_lrs3; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_ldst_val; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_nack_0_bits_uop_dst_rtype; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_nack_0_bits_uop_lrs1_rtype; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_nack_0_bits_uop_lrs2_rtype; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_frs3_en; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_fp_val; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_fp_single; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_xcpt_pf_if; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_xcpt_ae_if; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_xcpt_ma_if; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_bp_debug_if; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_uop_bp_xcpt_if; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_nack_0_bits_uop_debug_fsrc; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_nack_0_bits_uop_debug_tsrc; // @[tile.scala 134:54]
  wire [39:0] dcache_io_lsu_nack_0_bits_addr; // @[tile.scala 134:54]
  wire [63:0] dcache_io_lsu_nack_0_bits_data; // @[tile.scala 134:54]
  wire  dcache_io_lsu_nack_0_bits_is_hella; // @[tile.scala 134:54]
  wire [11:0] dcache_io_lsu_brupdate_b1_resolve_mask; // @[tile.scala 134:54]
  wire [11:0] dcache_io_lsu_brupdate_b1_mispredict_mask; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_switch; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_switch_off; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_is_unicore; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_brupdate_b2_uop_shift; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_brupdate_b2_uop_lrs3_rtype; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_rflag; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_wflag; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_brupdate_b2_uop_prflag; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_brupdate_b2_uop_pwflag; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_pflag_busy; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_brupdate_b2_uop_stale_pflag; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_brupdate_b2_uop_op1_sel; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_brupdate_b2_uop_op2_sel; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_brupdate_b2_uop_split_num; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_brupdate_b2_uop_self_index; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_brupdate_b2_uop_rob_inst_idx; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_brupdate_b2_uop_address_num; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_brupdate_b2_uop_uopc; // @[tile.scala 134:54]
  wire [31:0] dcache_io_lsu_brupdate_b2_uop_inst; // @[tile.scala 134:54]
  wire [31:0] dcache_io_lsu_brupdate_b2_uop_debug_inst; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_is_rvc; // @[tile.scala 134:54]
  wire [39:0] dcache_io_lsu_brupdate_b2_uop_debug_pc; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_brupdate_b2_uop_iq_type; // @[tile.scala 134:54]
  wire [9:0] dcache_io_lsu_brupdate_b2_uop_fu_code; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_brupdate_b2_uop_ctrl_br_type; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_brupdate_b2_uop_ctrl_op1_sel; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_brupdate_b2_uop_ctrl_op2_sel; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_brupdate_b2_uop_ctrl_imm_sel; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_brupdate_b2_uop_ctrl_op_fcn; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_ctrl_fcn_dw; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_brupdate_b2_uop_ctrl_csr_cmd; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_ctrl_is_load; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_ctrl_is_sta; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_ctrl_is_std; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_brupdate_b2_uop_ctrl_op3_sel; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_brupdate_b2_uop_iw_state; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_iw_p1_poisoned; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_iw_p2_poisoned; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_is_br; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_is_jalr; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_is_jal; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_is_sfb; // @[tile.scala 134:54]
  wire [11:0] dcache_io_lsu_brupdate_b2_uop_br_mask; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_brupdate_b2_uop_br_tag; // @[tile.scala 134:54]
  wire [4:0] dcache_io_lsu_brupdate_b2_uop_ftq_idx; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_edge_inst; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_brupdate_b2_uop_pc_lob; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_taken; // @[tile.scala 134:54]
  wire [19:0] dcache_io_lsu_brupdate_b2_uop_imm_packed; // @[tile.scala 134:54]
  wire [11:0] dcache_io_lsu_brupdate_b2_uop_csr_addr; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_brupdate_b2_uop_rob_idx; // @[tile.scala 134:54]
  wire [4:0] dcache_io_lsu_brupdate_b2_uop_ldq_idx; // @[tile.scala 134:54]
  wire [4:0] dcache_io_lsu_brupdate_b2_uop_stq_idx; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_brupdate_b2_uop_rxq_idx; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_brupdate_b2_uop_pdst; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_brupdate_b2_uop_prs1; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_brupdate_b2_uop_prs2; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_brupdate_b2_uop_prs3; // @[tile.scala 134:54]
  wire [4:0] dcache_io_lsu_brupdate_b2_uop_ppred; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_prs1_busy; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_prs2_busy; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_prs3_busy; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_ppred_busy; // @[tile.scala 134:54]
  wire [6:0] dcache_io_lsu_brupdate_b2_uop_stale_pdst; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_exception; // @[tile.scala 134:54]
  wire [63:0] dcache_io_lsu_brupdate_b2_uop_exc_cause; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_bypassable; // @[tile.scala 134:54]
  wire [4:0] dcache_io_lsu_brupdate_b2_uop_mem_cmd; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_brupdate_b2_uop_mem_size; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_mem_signed; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_is_fence; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_is_fencei; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_is_amo; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_uses_ldq; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_uses_stq; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_is_sys_pc2epc; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_is_unique; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_flush_on_commit; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_ldst_is_rs1; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_brupdate_b2_uop_ldst; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_brupdate_b2_uop_lrs1; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_brupdate_b2_uop_lrs2; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_brupdate_b2_uop_lrs3; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_ldst_val; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_brupdate_b2_uop_dst_rtype; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_brupdate_b2_uop_lrs1_rtype; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_brupdate_b2_uop_lrs2_rtype; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_frs3_en; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_fp_val; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_fp_single; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_xcpt_pf_if; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_xcpt_ae_if; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_xcpt_ma_if; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_bp_debug_if; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_uop_bp_xcpt_if; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_brupdate_b2_uop_debug_fsrc; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_brupdate_b2_uop_debug_tsrc; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_valid; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_mispredict; // @[tile.scala 134:54]
  wire  dcache_io_lsu_brupdate_b2_taken; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_brupdate_b2_cfi_type; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_brupdate_b2_pc_sel; // @[tile.scala 134:54]
  wire [39:0] dcache_io_lsu_brupdate_b2_jalr_target; // @[tile.scala 134:54]
  wire [31:0] dcache_io_lsu_brupdate_b2_target_offset; // @[tile.scala 134:54]
  wire  dcache_io_lsu_exception; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_rob_pnr_idx; // @[tile.scala 134:54]
  wire [5:0] dcache_io_lsu_rob_head_idx; // @[tile.scala 134:54]
  wire  dcache_io_lsu_release_ready; // @[tile.scala 134:54]
  wire  dcache_io_lsu_release_valid; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_release_bits_opcode; // @[tile.scala 134:54]
  wire [2:0] dcache_io_lsu_release_bits_param; // @[tile.scala 134:54]
  wire [3:0] dcache_io_lsu_release_bits_size; // @[tile.scala 134:54]
  wire [1:0] dcache_io_lsu_release_bits_source; // @[tile.scala 134:54]
  wire [31:0] dcache_io_lsu_release_bits_address; // @[tile.scala 134:54]
  wire [63:0] dcache_io_lsu_release_bits_data; // @[tile.scala 134:54]
  wire  dcache_io_lsu_release_bits_corrupt; // @[tile.scala 134:54]
  wire  dcache_io_lsu_force_order; // @[tile.scala 134:54]
  wire  dcache_io_lsu_ordered; // @[tile.scala 134:54]
  wire  dcache_io_lsu_perf_acquire; // @[tile.scala 134:54]
  wire  dcache_io_lsu_perf_release; // @[tile.scala 134:54]
  wire  frontend_clock; // @[tile.scala 140:28]
  wire  frontend_reset; // @[tile.scala 140:28]
  wire  frontend_auto_icache_master_out_a_ready; // @[tile.scala 140:28]
  wire  frontend_auto_icache_master_out_a_valid; // @[tile.scala 140:28]
  wire [2:0] frontend_auto_icache_master_out_a_bits_opcode; // @[tile.scala 140:28]
  wire [2:0] frontend_auto_icache_master_out_a_bits_param; // @[tile.scala 140:28]
  wire [3:0] frontend_auto_icache_master_out_a_bits_size; // @[tile.scala 140:28]
  wire  frontend_auto_icache_master_out_a_bits_source; // @[tile.scala 140:28]
  wire [31:0] frontend_auto_icache_master_out_a_bits_address; // @[tile.scala 140:28]
  wire [7:0] frontend_auto_icache_master_out_a_bits_mask; // @[tile.scala 140:28]
  wire [63:0] frontend_auto_icache_master_out_a_bits_data; // @[tile.scala 140:28]
  wire  frontend_auto_icache_master_out_a_bits_corrupt; // @[tile.scala 140:28]
  wire  frontend_auto_icache_master_out_d_ready; // @[tile.scala 140:28]
  wire  frontend_auto_icache_master_out_d_valid; // @[tile.scala 140:28]
  wire [2:0] frontend_auto_icache_master_out_d_bits_opcode; // @[tile.scala 140:28]
  wire [1:0] frontend_auto_icache_master_out_d_bits_param; // @[tile.scala 140:28]
  wire [3:0] frontend_auto_icache_master_out_d_bits_size; // @[tile.scala 140:28]
  wire  frontend_auto_icache_master_out_d_bits_source; // @[tile.scala 140:28]
  wire [1:0] frontend_auto_icache_master_out_d_bits_sink; // @[tile.scala 140:28]
  wire  frontend_auto_icache_master_out_d_bits_denied; // @[tile.scala 140:28]
  wire [63:0] frontend_auto_icache_master_out_d_bits_data; // @[tile.scala 140:28]
  wire  frontend_auto_icache_master_out_d_bits_corrupt; // @[tile.scala 140:28]
  wire [31:0] frontend_auto_reset_vector_sink_in; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_ready; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_valid; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_valid; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_switch; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_switch_off; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_unicore; // @[tile.scala 140:28]
  wire [2:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_shift; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_lrs3_rtype; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_rflag; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_wflag; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_prflag; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_pwflag; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_pflag_busy; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_stale_pflag; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_op1_sel; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_op2_sel; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_split_num; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_self_index; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_rob_inst_idx; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_address_num; // @[tile.scala 140:28]
  wire [6:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_uopc; // @[tile.scala 140:28]
  wire [31:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_inst; // @[tile.scala 140:28]
  wire [31:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_debug_inst; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_rvc; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_debug_pc; // @[tile.scala 140:28]
  wire [2:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_iq_type; // @[tile.scala 140:28]
  wire [9:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_fu_code; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_br_type; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_op1_sel; // @[tile.scala 140:28]
  wire [2:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_op2_sel; // @[tile.scala 140:28]
  wire [2:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_imm_sel; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_op_fcn; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_fcn_dw; // @[tile.scala 140:28]
  wire [2:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_csr_cmd; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_is_load; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_is_sta; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_is_std; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_op3_sel; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_iw_state; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_iw_p1_poisoned; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_iw_p2_poisoned; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_br; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_jalr; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_jal; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_sfb; // @[tile.scala 140:28]
  wire [11:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_br_mask; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_br_tag; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_ftq_idx; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_edge_inst; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_pc_lob; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_taken; // @[tile.scala 140:28]
  wire [19:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_imm_packed; // @[tile.scala 140:28]
  wire [11:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_csr_addr; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_rob_idx; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_ldq_idx; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_stq_idx; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_rxq_idx; // @[tile.scala 140:28]
  wire [6:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_pdst; // @[tile.scala 140:28]
  wire [6:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_prs1; // @[tile.scala 140:28]
  wire [6:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_prs2; // @[tile.scala 140:28]
  wire [6:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_prs3; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_ppred; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_prs1_busy; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_prs2_busy; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_prs3_busy; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_ppred_busy; // @[tile.scala 140:28]
  wire [6:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_stale_pdst; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_exception; // @[tile.scala 140:28]
  wire [63:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_exc_cause; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_bypassable; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_mem_cmd; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_mem_size; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_mem_signed; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_fence; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_fencei; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_amo; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_uses_ldq; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_uses_stq; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_sys_pc2epc; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_unique; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_flush_on_commit; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_ldst_is_rs1; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_ldst; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_lrs1; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_lrs2; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_lrs3; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_ldst_val; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_dst_rtype; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_lrs1_rtype; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_lrs2_rtype; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_frs3_en; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_fp_val; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_fp_single; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_xcpt_pf_if; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_xcpt_ae_if; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_xcpt_ma_if; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_bp_debug_if; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_0_bits_bp_xcpt_if; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_debug_fsrc; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_0_bits_debug_tsrc; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_valid; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_switch; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_switch_off; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_unicore; // @[tile.scala 140:28]
  wire [2:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_shift; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_lrs3_rtype; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_rflag; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_wflag; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_prflag; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_pwflag; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_pflag_busy; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_stale_pflag; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_op1_sel; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_op2_sel; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_split_num; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_self_index; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_rob_inst_idx; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_address_num; // @[tile.scala 140:28]
  wire [6:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_uopc; // @[tile.scala 140:28]
  wire [31:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_inst; // @[tile.scala 140:28]
  wire [31:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_debug_inst; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_rvc; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_debug_pc; // @[tile.scala 140:28]
  wire [2:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_iq_type; // @[tile.scala 140:28]
  wire [9:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_fu_code; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_br_type; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_op1_sel; // @[tile.scala 140:28]
  wire [2:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_op2_sel; // @[tile.scala 140:28]
  wire [2:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_imm_sel; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_op_fcn; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_fcn_dw; // @[tile.scala 140:28]
  wire [2:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_csr_cmd; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_is_load; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_is_sta; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_is_std; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_op3_sel; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_iw_state; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_iw_p1_poisoned; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_iw_p2_poisoned; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_br; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_jalr; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_jal; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_sfb; // @[tile.scala 140:28]
  wire [11:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_br_mask; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_br_tag; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_ftq_idx; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_edge_inst; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_pc_lob; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_taken; // @[tile.scala 140:28]
  wire [19:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_imm_packed; // @[tile.scala 140:28]
  wire [11:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_csr_addr; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_rob_idx; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_ldq_idx; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_stq_idx; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_rxq_idx; // @[tile.scala 140:28]
  wire [6:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_pdst; // @[tile.scala 140:28]
  wire [6:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_prs1; // @[tile.scala 140:28]
  wire [6:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_prs2; // @[tile.scala 140:28]
  wire [6:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_prs3; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_ppred; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_prs1_busy; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_prs2_busy; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_prs3_busy; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_ppred_busy; // @[tile.scala 140:28]
  wire [6:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_stale_pdst; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_exception; // @[tile.scala 140:28]
  wire [63:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_exc_cause; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_bypassable; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_mem_cmd; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_mem_size; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_mem_signed; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_fence; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_fencei; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_amo; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_uses_ldq; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_uses_stq; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_sys_pc2epc; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_unique; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_flush_on_commit; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_ldst_is_rs1; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_ldst; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_lrs1; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_lrs2; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_lrs3; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_ldst_val; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_dst_rtype; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_lrs1_rtype; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_lrs2_rtype; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_frs3_en; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_fp_val; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_fp_single; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_xcpt_pf_if; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_xcpt_ae_if; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_xcpt_ma_if; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_bp_debug_if; // @[tile.scala 140:28]
  wire  frontend_io_cpu_fetchpacket_bits_uops_1_bits_bp_xcpt_if; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_debug_fsrc; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_fetchpacket_bits_uops_1_bits_debug_tsrc; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_get_pc_0_ftq_idx; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_0_entry_cfi_idx_valid; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_get_pc_0_entry_cfi_idx_bits; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_0_entry_cfi_taken; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_0_entry_cfi_mispredicted; // @[tile.scala 140:28]
  wire [2:0] frontend_io_cpu_get_pc_0_entry_cfi_type; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_get_pc_0_entry_br_mask; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_0_entry_cfi_is_call; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_0_entry_cfi_is_ret; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_0_entry_cfi_npc_plus4; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_get_pc_0_entry_ras_top; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_get_pc_0_entry_ras_idx; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_0_entry_start_bank; // @[tile.scala 140:28]
  wire [15:0] frontend_io_cpu_get_pc_0_ghist_old_history; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_0_ghist_current_saw_branch_not_taken; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_0_ghist_new_saw_branch_not_taken; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_0_ghist_new_saw_branch_taken; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_get_pc_0_ghist_ras_idx; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_get_pc_0_pc; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_get_pc_0_com_pc; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_0_next_val; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_get_pc_0_next_pc; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_get_pc_1_ftq_idx; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_1_entry_cfi_idx_valid; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_get_pc_1_entry_cfi_idx_bits; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_1_entry_cfi_taken; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_1_entry_cfi_mispredicted; // @[tile.scala 140:28]
  wire [2:0] frontend_io_cpu_get_pc_1_entry_cfi_type; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_get_pc_1_entry_br_mask; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_1_entry_cfi_is_call; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_1_entry_cfi_is_ret; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_1_entry_cfi_npc_plus4; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_get_pc_1_entry_ras_top; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_get_pc_1_entry_ras_idx; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_1_entry_start_bank; // @[tile.scala 140:28]
  wire [15:0] frontend_io_cpu_get_pc_1_ghist_old_history; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_1_ghist_current_saw_branch_not_taken; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_1_ghist_new_saw_branch_not_taken; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_1_ghist_new_saw_branch_taken; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_get_pc_1_ghist_ras_idx; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_get_pc_1_pc; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_get_pc_1_com_pc; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_1_next_val; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_get_pc_1_next_pc; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_get_pc_2_ftq_idx; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_2_entry_cfi_idx_valid; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_get_pc_2_entry_cfi_idx_bits; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_2_entry_cfi_taken; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_2_entry_cfi_mispredicted; // @[tile.scala 140:28]
  wire [2:0] frontend_io_cpu_get_pc_2_entry_cfi_type; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_get_pc_2_entry_br_mask; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_2_entry_cfi_is_call; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_2_entry_cfi_is_ret; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_2_entry_cfi_npc_plus4; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_get_pc_2_entry_ras_top; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_get_pc_2_entry_ras_idx; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_2_entry_start_bank; // @[tile.scala 140:28]
  wire [15:0] frontend_io_cpu_get_pc_2_ghist_old_history; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_2_ghist_current_saw_branch_not_taken; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_2_ghist_new_saw_branch_not_taken; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_2_ghist_new_saw_branch_taken; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_get_pc_2_ghist_ras_idx; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_get_pc_2_pc; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_get_pc_2_com_pc; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_2_next_val; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_get_pc_2_next_pc; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_get_pc_3_ftq_idx; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_3_entry_cfi_idx_valid; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_get_pc_3_entry_cfi_idx_bits; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_3_entry_cfi_taken; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_3_entry_cfi_mispredicted; // @[tile.scala 140:28]
  wire [2:0] frontend_io_cpu_get_pc_3_entry_cfi_type; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_get_pc_3_entry_br_mask; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_3_entry_cfi_is_call; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_3_entry_cfi_is_ret; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_3_entry_cfi_npc_plus4; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_get_pc_3_entry_ras_top; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_get_pc_3_entry_ras_idx; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_3_entry_start_bank; // @[tile.scala 140:28]
  wire [15:0] frontend_io_cpu_get_pc_3_ghist_old_history; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_3_ghist_current_saw_branch_not_taken; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_3_ghist_new_saw_branch_not_taken; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_3_ghist_new_saw_branch_taken; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_get_pc_3_ghist_ras_idx; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_get_pc_3_pc; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_get_pc_3_com_pc; // @[tile.scala 140:28]
  wire  frontend_io_cpu_get_pc_3_next_val; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_get_pc_3_next_pc; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_debug_ftq_idx_0; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_debug_ftq_idx_1; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_debug_fetch_pc_0; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_debug_fetch_pc_1; // @[tile.scala 140:28]
  wire  frontend_io_cpu_status_debug; // @[tile.scala 140:28]
  wire  frontend_io_cpu_status_cease; // @[tile.scala 140:28]
  wire  frontend_io_cpu_status_wfi; // @[tile.scala 140:28]
  wire [31:0] frontend_io_cpu_status_isa; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_status_dprv; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_status_prv; // @[tile.scala 140:28]
  wire  frontend_io_cpu_status_sd; // @[tile.scala 140:28]
  wire [26:0] frontend_io_cpu_status_zero2; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_status_sxl; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_status_uxl; // @[tile.scala 140:28]
  wire  frontend_io_cpu_status_sd_rv32; // @[tile.scala 140:28]
  wire [7:0] frontend_io_cpu_status_zero1; // @[tile.scala 140:28]
  wire  frontend_io_cpu_status_tsr; // @[tile.scala 140:28]
  wire  frontend_io_cpu_status_tw; // @[tile.scala 140:28]
  wire  frontend_io_cpu_status_tvm; // @[tile.scala 140:28]
  wire  frontend_io_cpu_status_mxr; // @[tile.scala 140:28]
  wire  frontend_io_cpu_status_sum; // @[tile.scala 140:28]
  wire  frontend_io_cpu_status_mprv; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_status_xs; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_status_fs; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_status_mpp; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_status_vs; // @[tile.scala 140:28]
  wire  frontend_io_cpu_status_spp; // @[tile.scala 140:28]
  wire  frontend_io_cpu_status_mpie; // @[tile.scala 140:28]
  wire  frontend_io_cpu_status_hpie; // @[tile.scala 140:28]
  wire  frontend_io_cpu_status_spie; // @[tile.scala 140:28]
  wire  frontend_io_cpu_status_upie; // @[tile.scala 140:28]
  wire  frontend_io_cpu_status_mie; // @[tile.scala 140:28]
  wire  frontend_io_cpu_status_hie; // @[tile.scala 140:28]
  wire  frontend_io_cpu_status_sie; // @[tile.scala 140:28]
  wire  frontend_io_cpu_status_uie; // @[tile.scala 140:28]
  wire  frontend_io_cpu_sfence_valid; // @[tile.scala 140:28]
  wire  frontend_io_cpu_sfence_bits_rs1; // @[tile.scala 140:28]
  wire  frontend_io_cpu_sfence_bits_rs2; // @[tile.scala 140:28]
  wire [38:0] frontend_io_cpu_sfence_bits_addr; // @[tile.scala 140:28]
  wire  frontend_io_cpu_sfence_bits_asid; // @[tile.scala 140:28]
  wire [11:0] frontend_io_cpu_brupdate_b1_resolve_mask; // @[tile.scala 140:28]
  wire [11:0] frontend_io_cpu_brupdate_b1_mispredict_mask; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_switch; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_switch_off; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_is_unicore; // @[tile.scala 140:28]
  wire [2:0] frontend_io_cpu_brupdate_b2_uop_shift; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_brupdate_b2_uop_lrs3_rtype; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_rflag; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_wflag; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_brupdate_b2_uop_prflag; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_brupdate_b2_uop_pwflag; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_pflag_busy; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_brupdate_b2_uop_stale_pflag; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_brupdate_b2_uop_op1_sel; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_brupdate_b2_uop_op2_sel; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_brupdate_b2_uop_split_num; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_brupdate_b2_uop_self_index; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_brupdate_b2_uop_rob_inst_idx; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_brupdate_b2_uop_address_num; // @[tile.scala 140:28]
  wire [6:0] frontend_io_cpu_brupdate_b2_uop_uopc; // @[tile.scala 140:28]
  wire [31:0] frontend_io_cpu_brupdate_b2_uop_inst; // @[tile.scala 140:28]
  wire [31:0] frontend_io_cpu_brupdate_b2_uop_debug_inst; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_is_rvc; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_brupdate_b2_uop_debug_pc; // @[tile.scala 140:28]
  wire [2:0] frontend_io_cpu_brupdate_b2_uop_iq_type; // @[tile.scala 140:28]
  wire [9:0] frontend_io_cpu_brupdate_b2_uop_fu_code; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_brupdate_b2_uop_ctrl_br_type; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_brupdate_b2_uop_ctrl_op1_sel; // @[tile.scala 140:28]
  wire [2:0] frontend_io_cpu_brupdate_b2_uop_ctrl_op2_sel; // @[tile.scala 140:28]
  wire [2:0] frontend_io_cpu_brupdate_b2_uop_ctrl_imm_sel; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_brupdate_b2_uop_ctrl_op_fcn; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_ctrl_fcn_dw; // @[tile.scala 140:28]
  wire [2:0] frontend_io_cpu_brupdate_b2_uop_ctrl_csr_cmd; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_ctrl_is_load; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_ctrl_is_sta; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_ctrl_is_std; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_brupdate_b2_uop_ctrl_op3_sel; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_brupdate_b2_uop_iw_state; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_iw_p1_poisoned; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_iw_p2_poisoned; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_is_br; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_is_jalr; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_is_jal; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_is_sfb; // @[tile.scala 140:28]
  wire [11:0] frontend_io_cpu_brupdate_b2_uop_br_mask; // @[tile.scala 140:28]
  wire [3:0] frontend_io_cpu_brupdate_b2_uop_br_tag; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_brupdate_b2_uop_ftq_idx; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_edge_inst; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_brupdate_b2_uop_pc_lob; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_taken; // @[tile.scala 140:28]
  wire [19:0] frontend_io_cpu_brupdate_b2_uop_imm_packed; // @[tile.scala 140:28]
  wire [11:0] frontend_io_cpu_brupdate_b2_uop_csr_addr; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_brupdate_b2_uop_rob_idx; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_brupdate_b2_uop_ldq_idx; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_brupdate_b2_uop_stq_idx; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_brupdate_b2_uop_rxq_idx; // @[tile.scala 140:28]
  wire [6:0] frontend_io_cpu_brupdate_b2_uop_pdst; // @[tile.scala 140:28]
  wire [6:0] frontend_io_cpu_brupdate_b2_uop_prs1; // @[tile.scala 140:28]
  wire [6:0] frontend_io_cpu_brupdate_b2_uop_prs2; // @[tile.scala 140:28]
  wire [6:0] frontend_io_cpu_brupdate_b2_uop_prs3; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_brupdate_b2_uop_ppred; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_prs1_busy; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_prs2_busy; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_prs3_busy; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_ppred_busy; // @[tile.scala 140:28]
  wire [6:0] frontend_io_cpu_brupdate_b2_uop_stale_pdst; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_exception; // @[tile.scala 140:28]
  wire [63:0] frontend_io_cpu_brupdate_b2_uop_exc_cause; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_bypassable; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_brupdate_b2_uop_mem_cmd; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_brupdate_b2_uop_mem_size; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_mem_signed; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_is_fence; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_is_fencei; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_is_amo; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_uses_ldq; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_uses_stq; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_is_sys_pc2epc; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_is_unique; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_flush_on_commit; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_ldst_is_rs1; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_brupdate_b2_uop_ldst; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_brupdate_b2_uop_lrs1; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_brupdate_b2_uop_lrs2; // @[tile.scala 140:28]
  wire [5:0] frontend_io_cpu_brupdate_b2_uop_lrs3; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_ldst_val; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_brupdate_b2_uop_dst_rtype; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_brupdate_b2_uop_lrs1_rtype; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_brupdate_b2_uop_lrs2_rtype; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_frs3_en; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_fp_val; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_fp_single; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_xcpt_pf_if; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_xcpt_ae_if; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_xcpt_ma_if; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_bp_debug_if; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_uop_bp_xcpt_if; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_brupdate_b2_uop_debug_fsrc; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_brupdate_b2_uop_debug_tsrc; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_valid; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_mispredict; // @[tile.scala 140:28]
  wire  frontend_io_cpu_brupdate_b2_taken; // @[tile.scala 140:28]
  wire [2:0] frontend_io_cpu_brupdate_b2_cfi_type; // @[tile.scala 140:28]
  wire [1:0] frontend_io_cpu_brupdate_b2_pc_sel; // @[tile.scala 140:28]
  wire [39:0] frontend_io_cpu_brupdate_b2_jalr_target; // @[tile.scala 140:28]
  wire [31:0] frontend_io_cpu_brupdate_b2_target_offset; // @[tile.scala 140:28]
  wire  frontend_io_cpu_redirect_flush; // @[tile.scala 140:28]
  wire  frontend_io_cpu_redirect_val; // @[tile.scala 140:28]
  wire [63:0] frontend_io_cpu_redirect_pc; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_redirect_ftq_idx; // @[tile.scala 140:28]
  wire [15:0] frontend_io_cpu_redirect_ghist_old_history; // @[tile.scala 140:28]
  wire  frontend_io_cpu_redirect_ghist_current_saw_branch_not_taken; // @[tile.scala 140:28]
  wire  frontend_io_cpu_redirect_ghist_new_saw_branch_not_taken; // @[tile.scala 140:28]
  wire  frontend_io_cpu_redirect_ghist_new_saw_branch_taken; // @[tile.scala 140:28]
  wire [4:0] frontend_io_cpu_redirect_ghist_ras_idx; // @[tile.scala 140:28]
  wire  frontend_io_cpu_commit_valid; // @[tile.scala 140:28]
  wire [31:0] frontend_io_cpu_commit_bits; // @[tile.scala 140:28]
  wire  frontend_io_cpu_flush_icache; // @[tile.scala 140:28]
  wire  frontend_io_cpu_perf_acquire; // @[tile.scala 140:28]
  wire  frontend_io_cpu_perf_tlbMiss; // @[tile.scala 140:28]
  wire  frontend_io_cpu_is_unicore; // @[tile.scala 140:28]
  wire  frontend_io_ptw_req_ready; // @[tile.scala 140:28]
  wire  frontend_io_ptw_req_valid; // @[tile.scala 140:28]
  wire  frontend_io_ptw_req_bits_valid; // @[tile.scala 140:28]
  wire [26:0] frontend_io_ptw_req_bits_bits_addr; // @[tile.scala 140:28]
  wire  frontend_io_ptw_resp_valid; // @[tile.scala 140:28]
  wire  frontend_io_ptw_resp_bits_ae; // @[tile.scala 140:28]
  wire [53:0] frontend_io_ptw_resp_bits_pte_ppn; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_resp_bits_pte_reserved_for_software; // @[tile.scala 140:28]
  wire  frontend_io_ptw_resp_bits_pte_d; // @[tile.scala 140:28]
  wire  frontend_io_ptw_resp_bits_pte_a; // @[tile.scala 140:28]
  wire  frontend_io_ptw_resp_bits_pte_g; // @[tile.scala 140:28]
  wire  frontend_io_ptw_resp_bits_pte_u; // @[tile.scala 140:28]
  wire  frontend_io_ptw_resp_bits_pte_x; // @[tile.scala 140:28]
  wire  frontend_io_ptw_resp_bits_pte_w; // @[tile.scala 140:28]
  wire  frontend_io_ptw_resp_bits_pte_r; // @[tile.scala 140:28]
  wire  frontend_io_ptw_resp_bits_pte_v; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_resp_bits_level; // @[tile.scala 140:28]
  wire  frontend_io_ptw_resp_bits_fragmented_superpage; // @[tile.scala 140:28]
  wire  frontend_io_ptw_resp_bits_homogeneous; // @[tile.scala 140:28]
  wire [3:0] frontend_io_ptw_ptbr_mode; // @[tile.scala 140:28]
  wire [15:0] frontend_io_ptw_ptbr_asid; // @[tile.scala 140:28]
  wire [43:0] frontend_io_ptw_ptbr_ppn; // @[tile.scala 140:28]
  wire  frontend_io_ptw_status_debug; // @[tile.scala 140:28]
  wire  frontend_io_ptw_status_cease; // @[tile.scala 140:28]
  wire  frontend_io_ptw_status_wfi; // @[tile.scala 140:28]
  wire [31:0] frontend_io_ptw_status_isa; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_status_dprv; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_status_prv; // @[tile.scala 140:28]
  wire  frontend_io_ptw_status_sd; // @[tile.scala 140:28]
  wire [26:0] frontend_io_ptw_status_zero2; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_status_sxl; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_status_uxl; // @[tile.scala 140:28]
  wire  frontend_io_ptw_status_sd_rv32; // @[tile.scala 140:28]
  wire [7:0] frontend_io_ptw_status_zero1; // @[tile.scala 140:28]
  wire  frontend_io_ptw_status_tsr; // @[tile.scala 140:28]
  wire  frontend_io_ptw_status_tw; // @[tile.scala 140:28]
  wire  frontend_io_ptw_status_tvm; // @[tile.scala 140:28]
  wire  frontend_io_ptw_status_mxr; // @[tile.scala 140:28]
  wire  frontend_io_ptw_status_sum; // @[tile.scala 140:28]
  wire  frontend_io_ptw_status_mprv; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_status_xs; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_status_fs; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_status_mpp; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_status_vs; // @[tile.scala 140:28]
  wire  frontend_io_ptw_status_spp; // @[tile.scala 140:28]
  wire  frontend_io_ptw_status_mpie; // @[tile.scala 140:28]
  wire  frontend_io_ptw_status_hpie; // @[tile.scala 140:28]
  wire  frontend_io_ptw_status_spie; // @[tile.scala 140:28]
  wire  frontend_io_ptw_status_upie; // @[tile.scala 140:28]
  wire  frontend_io_ptw_status_mie; // @[tile.scala 140:28]
  wire  frontend_io_ptw_status_hie; // @[tile.scala 140:28]
  wire  frontend_io_ptw_status_sie; // @[tile.scala 140:28]
  wire  frontend_io_ptw_status_uie; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_0_cfg_l; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_pmp_0_cfg_res; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_pmp_0_cfg_a; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_0_cfg_x; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_0_cfg_w; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_0_cfg_r; // @[tile.scala 140:28]
  wire [29:0] frontend_io_ptw_pmp_0_addr; // @[tile.scala 140:28]
  wire [31:0] frontend_io_ptw_pmp_0_mask; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_1_cfg_l; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_pmp_1_cfg_res; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_pmp_1_cfg_a; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_1_cfg_x; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_1_cfg_w; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_1_cfg_r; // @[tile.scala 140:28]
  wire [29:0] frontend_io_ptw_pmp_1_addr; // @[tile.scala 140:28]
  wire [31:0] frontend_io_ptw_pmp_1_mask; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_2_cfg_l; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_pmp_2_cfg_res; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_pmp_2_cfg_a; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_2_cfg_x; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_2_cfg_w; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_2_cfg_r; // @[tile.scala 140:28]
  wire [29:0] frontend_io_ptw_pmp_2_addr; // @[tile.scala 140:28]
  wire [31:0] frontend_io_ptw_pmp_2_mask; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_3_cfg_l; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_pmp_3_cfg_res; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_pmp_3_cfg_a; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_3_cfg_x; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_3_cfg_w; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_3_cfg_r; // @[tile.scala 140:28]
  wire [29:0] frontend_io_ptw_pmp_3_addr; // @[tile.scala 140:28]
  wire [31:0] frontend_io_ptw_pmp_3_mask; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_4_cfg_l; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_pmp_4_cfg_res; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_pmp_4_cfg_a; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_4_cfg_x; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_4_cfg_w; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_4_cfg_r; // @[tile.scala 140:28]
  wire [29:0] frontend_io_ptw_pmp_4_addr; // @[tile.scala 140:28]
  wire [31:0] frontend_io_ptw_pmp_4_mask; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_5_cfg_l; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_pmp_5_cfg_res; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_pmp_5_cfg_a; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_5_cfg_x; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_5_cfg_w; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_5_cfg_r; // @[tile.scala 140:28]
  wire [29:0] frontend_io_ptw_pmp_5_addr; // @[tile.scala 140:28]
  wire [31:0] frontend_io_ptw_pmp_5_mask; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_6_cfg_l; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_pmp_6_cfg_res; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_pmp_6_cfg_a; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_6_cfg_x; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_6_cfg_w; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_6_cfg_r; // @[tile.scala 140:28]
  wire [29:0] frontend_io_ptw_pmp_6_addr; // @[tile.scala 140:28]
  wire [31:0] frontend_io_ptw_pmp_6_mask; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_7_cfg_l; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_pmp_7_cfg_res; // @[tile.scala 140:28]
  wire [1:0] frontend_io_ptw_pmp_7_cfg_a; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_7_cfg_x; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_7_cfg_w; // @[tile.scala 140:28]
  wire  frontend_io_ptw_pmp_7_cfg_r; // @[tile.scala 140:28]
  wire [29:0] frontend_io_ptw_pmp_7_addr; // @[tile.scala 140:28]
  wire [31:0] frontend_io_ptw_pmp_7_mask; // @[tile.scala 140:28]
  wire  frontend_io_ptw_customCSRs_csrs_0_wen; // @[tile.scala 140:28]
  wire [63:0] frontend_io_ptw_customCSRs_csrs_0_wdata; // @[tile.scala 140:28]
  wire [63:0] frontend_io_ptw_customCSRs_csrs_0_value; // @[tile.scala 140:28]
  wire  frontend_io_errors_bus_valid; // @[tile.scala 140:28]
  wire [31:0] frontend_io_errors_bus_bits; // @[tile.scala 140:28]
  wire  core_clock; // @[tile.scala 159:20]
  wire  core_reset; // @[tile.scala 159:20]
  wire  core_io_hartid; // @[tile.scala 159:20]
  wire  core_io_interrupts_debug; // @[tile.scala 159:20]
  wire  core_io_interrupts_mtip; // @[tile.scala 159:20]
  wire  core_io_interrupts_msip; // @[tile.scala 159:20]
  wire  core_io_interrupts_meip; // @[tile.scala 159:20]
  wire  core_io_interrupts_seip; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_ready; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_valid; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_valid; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_switch; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_switch_off; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_is_unicore; // @[tile.scala 159:20]
  wire [2:0] core_io_ifu_fetchpacket_bits_uops_0_bits_shift; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_0_bits_lrs3_rtype; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_rflag; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_wflag; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_fetchpacket_bits_uops_0_bits_prflag; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_fetchpacket_bits_uops_0_bits_pwflag; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_pflag_busy; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_fetchpacket_bits_uops_0_bits_stale_pflag; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_fetchpacket_bits_uops_0_bits_op1_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_fetchpacket_bits_uops_0_bits_op2_sel; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_fetchpacket_bits_uops_0_bits_split_num; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_fetchpacket_bits_uops_0_bits_self_index; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_fetchpacket_bits_uops_0_bits_rob_inst_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_fetchpacket_bits_uops_0_bits_address_num; // @[tile.scala 159:20]
  wire [6:0] core_io_ifu_fetchpacket_bits_uops_0_bits_uopc; // @[tile.scala 159:20]
  wire [31:0] core_io_ifu_fetchpacket_bits_uops_0_bits_inst; // @[tile.scala 159:20]
  wire [31:0] core_io_ifu_fetchpacket_bits_uops_0_bits_debug_inst; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_is_rvc; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_fetchpacket_bits_uops_0_bits_debug_pc; // @[tile.scala 159:20]
  wire [2:0] core_io_ifu_fetchpacket_bits_uops_0_bits_iq_type; // @[tile.scala 159:20]
  wire [9:0] core_io_ifu_fetchpacket_bits_uops_0_bits_fu_code; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_br_type; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_op1_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_op2_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_imm_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_op_fcn; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_fcn_dw; // @[tile.scala 159:20]
  wire [2:0] core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_csr_cmd; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_is_load; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_is_sta; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_is_std; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_op3_sel; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_0_bits_iw_state; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_iw_p1_poisoned; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_iw_p2_poisoned; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_is_br; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_is_jalr; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_is_jal; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_is_sfb; // @[tile.scala 159:20]
  wire [11:0] core_io_ifu_fetchpacket_bits_uops_0_bits_br_mask; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_fetchpacket_bits_uops_0_bits_br_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_fetchpacket_bits_uops_0_bits_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_edge_inst; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_fetchpacket_bits_uops_0_bits_pc_lob; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_taken; // @[tile.scala 159:20]
  wire [19:0] core_io_ifu_fetchpacket_bits_uops_0_bits_imm_packed; // @[tile.scala 159:20]
  wire [11:0] core_io_ifu_fetchpacket_bits_uops_0_bits_csr_addr; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_fetchpacket_bits_uops_0_bits_rob_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_fetchpacket_bits_uops_0_bits_ldq_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_fetchpacket_bits_uops_0_bits_stq_idx; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_0_bits_rxq_idx; // @[tile.scala 159:20]
  wire [6:0] core_io_ifu_fetchpacket_bits_uops_0_bits_pdst; // @[tile.scala 159:20]
  wire [6:0] core_io_ifu_fetchpacket_bits_uops_0_bits_prs1; // @[tile.scala 159:20]
  wire [6:0] core_io_ifu_fetchpacket_bits_uops_0_bits_prs2; // @[tile.scala 159:20]
  wire [6:0] core_io_ifu_fetchpacket_bits_uops_0_bits_prs3; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_fetchpacket_bits_uops_0_bits_ppred; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_prs1_busy; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_prs2_busy; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_prs3_busy; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_ppred_busy; // @[tile.scala 159:20]
  wire [6:0] core_io_ifu_fetchpacket_bits_uops_0_bits_stale_pdst; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_exception; // @[tile.scala 159:20]
  wire [63:0] core_io_ifu_fetchpacket_bits_uops_0_bits_exc_cause; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_bypassable; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_fetchpacket_bits_uops_0_bits_mem_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_0_bits_mem_size; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_mem_signed; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_is_fence; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_is_fencei; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_is_amo; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_uses_ldq; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_uses_stq; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_is_sys_pc2epc; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_is_unique; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_flush_on_commit; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_ldst_is_rs1; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_fetchpacket_bits_uops_0_bits_ldst; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_fetchpacket_bits_uops_0_bits_lrs1; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_fetchpacket_bits_uops_0_bits_lrs2; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_fetchpacket_bits_uops_0_bits_lrs3; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_ldst_val; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_0_bits_dst_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_0_bits_lrs1_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_0_bits_lrs2_rtype; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_frs3_en; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_fp_val; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_fp_single; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_xcpt_pf_if; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_xcpt_ae_if; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_xcpt_ma_if; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_bp_debug_if; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_0_bits_bp_xcpt_if; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_0_bits_debug_fsrc; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_0_bits_debug_tsrc; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_valid; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_switch; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_switch_off; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_is_unicore; // @[tile.scala 159:20]
  wire [2:0] core_io_ifu_fetchpacket_bits_uops_1_bits_shift; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_1_bits_lrs3_rtype; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_rflag; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_wflag; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_fetchpacket_bits_uops_1_bits_prflag; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_fetchpacket_bits_uops_1_bits_pwflag; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_pflag_busy; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_fetchpacket_bits_uops_1_bits_stale_pflag; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_fetchpacket_bits_uops_1_bits_op1_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_fetchpacket_bits_uops_1_bits_op2_sel; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_fetchpacket_bits_uops_1_bits_split_num; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_fetchpacket_bits_uops_1_bits_self_index; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_fetchpacket_bits_uops_1_bits_rob_inst_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_fetchpacket_bits_uops_1_bits_address_num; // @[tile.scala 159:20]
  wire [6:0] core_io_ifu_fetchpacket_bits_uops_1_bits_uopc; // @[tile.scala 159:20]
  wire [31:0] core_io_ifu_fetchpacket_bits_uops_1_bits_inst; // @[tile.scala 159:20]
  wire [31:0] core_io_ifu_fetchpacket_bits_uops_1_bits_debug_inst; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_is_rvc; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_fetchpacket_bits_uops_1_bits_debug_pc; // @[tile.scala 159:20]
  wire [2:0] core_io_ifu_fetchpacket_bits_uops_1_bits_iq_type; // @[tile.scala 159:20]
  wire [9:0] core_io_ifu_fetchpacket_bits_uops_1_bits_fu_code; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_br_type; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_op1_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_op2_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_imm_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_op_fcn; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_fcn_dw; // @[tile.scala 159:20]
  wire [2:0] core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_csr_cmd; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_is_load; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_is_sta; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_is_std; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_op3_sel; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_1_bits_iw_state; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_iw_p1_poisoned; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_iw_p2_poisoned; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_is_br; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_is_jalr; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_is_jal; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_is_sfb; // @[tile.scala 159:20]
  wire [11:0] core_io_ifu_fetchpacket_bits_uops_1_bits_br_mask; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_fetchpacket_bits_uops_1_bits_br_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_fetchpacket_bits_uops_1_bits_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_edge_inst; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_fetchpacket_bits_uops_1_bits_pc_lob; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_taken; // @[tile.scala 159:20]
  wire [19:0] core_io_ifu_fetchpacket_bits_uops_1_bits_imm_packed; // @[tile.scala 159:20]
  wire [11:0] core_io_ifu_fetchpacket_bits_uops_1_bits_csr_addr; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_fetchpacket_bits_uops_1_bits_rob_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_fetchpacket_bits_uops_1_bits_ldq_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_fetchpacket_bits_uops_1_bits_stq_idx; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_1_bits_rxq_idx; // @[tile.scala 159:20]
  wire [6:0] core_io_ifu_fetchpacket_bits_uops_1_bits_pdst; // @[tile.scala 159:20]
  wire [6:0] core_io_ifu_fetchpacket_bits_uops_1_bits_prs1; // @[tile.scala 159:20]
  wire [6:0] core_io_ifu_fetchpacket_bits_uops_1_bits_prs2; // @[tile.scala 159:20]
  wire [6:0] core_io_ifu_fetchpacket_bits_uops_1_bits_prs3; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_fetchpacket_bits_uops_1_bits_ppred; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_prs1_busy; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_prs2_busy; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_prs3_busy; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_ppred_busy; // @[tile.scala 159:20]
  wire [6:0] core_io_ifu_fetchpacket_bits_uops_1_bits_stale_pdst; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_exception; // @[tile.scala 159:20]
  wire [63:0] core_io_ifu_fetchpacket_bits_uops_1_bits_exc_cause; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_bypassable; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_fetchpacket_bits_uops_1_bits_mem_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_1_bits_mem_size; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_mem_signed; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_is_fence; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_is_fencei; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_is_amo; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_uses_ldq; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_uses_stq; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_is_sys_pc2epc; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_is_unique; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_flush_on_commit; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_ldst_is_rs1; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_fetchpacket_bits_uops_1_bits_ldst; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_fetchpacket_bits_uops_1_bits_lrs1; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_fetchpacket_bits_uops_1_bits_lrs2; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_fetchpacket_bits_uops_1_bits_lrs3; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_ldst_val; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_1_bits_dst_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_1_bits_lrs1_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_1_bits_lrs2_rtype; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_frs3_en; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_fp_val; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_fp_single; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_xcpt_pf_if; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_xcpt_ae_if; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_xcpt_ma_if; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_bp_debug_if; // @[tile.scala 159:20]
  wire  core_io_ifu_fetchpacket_bits_uops_1_bits_bp_xcpt_if; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_1_bits_debug_fsrc; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_fetchpacket_bits_uops_1_bits_debug_tsrc; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_get_pc_0_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_0_entry_cfi_idx_valid; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_get_pc_0_entry_cfi_idx_bits; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_0_entry_cfi_taken; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_0_entry_cfi_mispredicted; // @[tile.scala 159:20]
  wire [2:0] core_io_ifu_get_pc_0_entry_cfi_type; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_get_pc_0_entry_br_mask; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_0_entry_cfi_is_call; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_0_entry_cfi_is_ret; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_0_entry_cfi_npc_plus4; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_get_pc_0_entry_ras_top; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_get_pc_0_entry_ras_idx; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_0_entry_start_bank; // @[tile.scala 159:20]
  wire [15:0] core_io_ifu_get_pc_0_ghist_old_history; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_0_ghist_current_saw_branch_not_taken; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_0_ghist_new_saw_branch_not_taken; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_0_ghist_new_saw_branch_taken; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_get_pc_0_ghist_ras_idx; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_get_pc_0_pc; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_get_pc_0_com_pc; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_0_next_val; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_get_pc_0_next_pc; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_get_pc_1_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_1_entry_cfi_idx_valid; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_get_pc_1_entry_cfi_idx_bits; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_1_entry_cfi_taken; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_1_entry_cfi_mispredicted; // @[tile.scala 159:20]
  wire [2:0] core_io_ifu_get_pc_1_entry_cfi_type; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_get_pc_1_entry_br_mask; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_1_entry_cfi_is_call; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_1_entry_cfi_is_ret; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_1_entry_cfi_npc_plus4; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_get_pc_1_entry_ras_top; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_get_pc_1_entry_ras_idx; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_1_entry_start_bank; // @[tile.scala 159:20]
  wire [15:0] core_io_ifu_get_pc_1_ghist_old_history; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_1_ghist_current_saw_branch_not_taken; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_1_ghist_new_saw_branch_not_taken; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_1_ghist_new_saw_branch_taken; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_get_pc_1_ghist_ras_idx; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_get_pc_1_pc; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_get_pc_1_com_pc; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_1_next_val; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_get_pc_1_next_pc; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_get_pc_2_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_2_entry_cfi_idx_valid; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_get_pc_2_entry_cfi_idx_bits; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_2_entry_cfi_taken; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_2_entry_cfi_mispredicted; // @[tile.scala 159:20]
  wire [2:0] core_io_ifu_get_pc_2_entry_cfi_type; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_get_pc_2_entry_br_mask; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_2_entry_cfi_is_call; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_2_entry_cfi_is_ret; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_2_entry_cfi_npc_plus4; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_get_pc_2_entry_ras_top; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_get_pc_2_entry_ras_idx; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_2_entry_start_bank; // @[tile.scala 159:20]
  wire [15:0] core_io_ifu_get_pc_2_ghist_old_history; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_2_ghist_current_saw_branch_not_taken; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_2_ghist_new_saw_branch_not_taken; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_2_ghist_new_saw_branch_taken; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_get_pc_2_ghist_ras_idx; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_get_pc_2_pc; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_get_pc_2_com_pc; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_2_next_val; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_get_pc_2_next_pc; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_get_pc_3_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_3_entry_cfi_idx_valid; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_get_pc_3_entry_cfi_idx_bits; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_3_entry_cfi_taken; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_3_entry_cfi_mispredicted; // @[tile.scala 159:20]
  wire [2:0] core_io_ifu_get_pc_3_entry_cfi_type; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_get_pc_3_entry_br_mask; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_3_entry_cfi_is_call; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_3_entry_cfi_is_ret; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_3_entry_cfi_npc_plus4; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_get_pc_3_entry_ras_top; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_get_pc_3_entry_ras_idx; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_3_entry_start_bank; // @[tile.scala 159:20]
  wire [15:0] core_io_ifu_get_pc_3_ghist_old_history; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_3_ghist_current_saw_branch_not_taken; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_3_ghist_new_saw_branch_not_taken; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_3_ghist_new_saw_branch_taken; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_get_pc_3_ghist_ras_idx; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_get_pc_3_pc; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_get_pc_3_com_pc; // @[tile.scala 159:20]
  wire  core_io_ifu_get_pc_3_next_val; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_get_pc_3_next_pc; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_debug_ftq_idx_0; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_debug_ftq_idx_1; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_debug_fetch_pc_0; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_debug_fetch_pc_1; // @[tile.scala 159:20]
  wire  core_io_ifu_status_debug; // @[tile.scala 159:20]
  wire  core_io_ifu_status_cease; // @[tile.scala 159:20]
  wire  core_io_ifu_status_wfi; // @[tile.scala 159:20]
  wire [31:0] core_io_ifu_status_isa; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_status_dprv; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_status_prv; // @[tile.scala 159:20]
  wire  core_io_ifu_status_sd; // @[tile.scala 159:20]
  wire [26:0] core_io_ifu_status_zero2; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_status_sxl; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_status_uxl; // @[tile.scala 159:20]
  wire  core_io_ifu_status_sd_rv32; // @[tile.scala 159:20]
  wire [7:0] core_io_ifu_status_zero1; // @[tile.scala 159:20]
  wire  core_io_ifu_status_tsr; // @[tile.scala 159:20]
  wire  core_io_ifu_status_tw; // @[tile.scala 159:20]
  wire  core_io_ifu_status_tvm; // @[tile.scala 159:20]
  wire  core_io_ifu_status_mxr; // @[tile.scala 159:20]
  wire  core_io_ifu_status_sum; // @[tile.scala 159:20]
  wire  core_io_ifu_status_mprv; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_status_xs; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_status_fs; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_status_mpp; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_status_vs; // @[tile.scala 159:20]
  wire  core_io_ifu_status_spp; // @[tile.scala 159:20]
  wire  core_io_ifu_status_mpie; // @[tile.scala 159:20]
  wire  core_io_ifu_status_hpie; // @[tile.scala 159:20]
  wire  core_io_ifu_status_spie; // @[tile.scala 159:20]
  wire  core_io_ifu_status_upie; // @[tile.scala 159:20]
  wire  core_io_ifu_status_mie; // @[tile.scala 159:20]
  wire  core_io_ifu_status_hie; // @[tile.scala 159:20]
  wire  core_io_ifu_status_sie; // @[tile.scala 159:20]
  wire  core_io_ifu_status_uie; // @[tile.scala 159:20]
  wire  core_io_ifu_sfence_valid; // @[tile.scala 159:20]
  wire  core_io_ifu_sfence_bits_rs1; // @[tile.scala 159:20]
  wire  core_io_ifu_sfence_bits_rs2; // @[tile.scala 159:20]
  wire [38:0] core_io_ifu_sfence_bits_addr; // @[tile.scala 159:20]
  wire  core_io_ifu_sfence_bits_asid; // @[tile.scala 159:20]
  wire [11:0] core_io_ifu_brupdate_b1_resolve_mask; // @[tile.scala 159:20]
  wire [11:0] core_io_ifu_brupdate_b1_mispredict_mask; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_switch; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_switch_off; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_is_unicore; // @[tile.scala 159:20]
  wire [2:0] core_io_ifu_brupdate_b2_uop_shift; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_brupdate_b2_uop_lrs3_rtype; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_rflag; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_wflag; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_brupdate_b2_uop_prflag; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_brupdate_b2_uop_pwflag; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_pflag_busy; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_brupdate_b2_uop_stale_pflag; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_brupdate_b2_uop_op1_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_brupdate_b2_uop_op2_sel; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_brupdate_b2_uop_split_num; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_brupdate_b2_uop_self_index; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_brupdate_b2_uop_rob_inst_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_brupdate_b2_uop_address_num; // @[tile.scala 159:20]
  wire [6:0] core_io_ifu_brupdate_b2_uop_uopc; // @[tile.scala 159:20]
  wire [31:0] core_io_ifu_brupdate_b2_uop_inst; // @[tile.scala 159:20]
  wire [31:0] core_io_ifu_brupdate_b2_uop_debug_inst; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_is_rvc; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_brupdate_b2_uop_debug_pc; // @[tile.scala 159:20]
  wire [2:0] core_io_ifu_brupdate_b2_uop_iq_type; // @[tile.scala 159:20]
  wire [9:0] core_io_ifu_brupdate_b2_uop_fu_code; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_brupdate_b2_uop_ctrl_br_type; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_brupdate_b2_uop_ctrl_op1_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_ifu_brupdate_b2_uop_ctrl_op2_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_ifu_brupdate_b2_uop_ctrl_imm_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_brupdate_b2_uop_ctrl_op_fcn; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_ctrl_fcn_dw; // @[tile.scala 159:20]
  wire [2:0] core_io_ifu_brupdate_b2_uop_ctrl_csr_cmd; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_ctrl_is_load; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_ctrl_is_sta; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_ctrl_is_std; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_brupdate_b2_uop_ctrl_op3_sel; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_brupdate_b2_uop_iw_state; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_iw_p1_poisoned; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_iw_p2_poisoned; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_is_br; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_is_jalr; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_is_jal; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_is_sfb; // @[tile.scala 159:20]
  wire [11:0] core_io_ifu_brupdate_b2_uop_br_mask; // @[tile.scala 159:20]
  wire [3:0] core_io_ifu_brupdate_b2_uop_br_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_brupdate_b2_uop_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_edge_inst; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_brupdate_b2_uop_pc_lob; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_taken; // @[tile.scala 159:20]
  wire [19:0] core_io_ifu_brupdate_b2_uop_imm_packed; // @[tile.scala 159:20]
  wire [11:0] core_io_ifu_brupdate_b2_uop_csr_addr; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_brupdate_b2_uop_rob_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_brupdate_b2_uop_ldq_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_brupdate_b2_uop_stq_idx; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_brupdate_b2_uop_rxq_idx; // @[tile.scala 159:20]
  wire [6:0] core_io_ifu_brupdate_b2_uop_pdst; // @[tile.scala 159:20]
  wire [6:0] core_io_ifu_brupdate_b2_uop_prs1; // @[tile.scala 159:20]
  wire [6:0] core_io_ifu_brupdate_b2_uop_prs2; // @[tile.scala 159:20]
  wire [6:0] core_io_ifu_brupdate_b2_uop_prs3; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_brupdate_b2_uop_ppred; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_prs1_busy; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_prs2_busy; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_prs3_busy; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_ppred_busy; // @[tile.scala 159:20]
  wire [6:0] core_io_ifu_brupdate_b2_uop_stale_pdst; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_exception; // @[tile.scala 159:20]
  wire [63:0] core_io_ifu_brupdate_b2_uop_exc_cause; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_bypassable; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_brupdate_b2_uop_mem_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_brupdate_b2_uop_mem_size; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_mem_signed; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_is_fence; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_is_fencei; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_is_amo; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_uses_ldq; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_uses_stq; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_is_sys_pc2epc; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_is_unique; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_flush_on_commit; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_ldst_is_rs1; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_brupdate_b2_uop_ldst; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_brupdate_b2_uop_lrs1; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_brupdate_b2_uop_lrs2; // @[tile.scala 159:20]
  wire [5:0] core_io_ifu_brupdate_b2_uop_lrs3; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_ldst_val; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_brupdate_b2_uop_dst_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_brupdate_b2_uop_lrs1_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_brupdate_b2_uop_lrs2_rtype; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_frs3_en; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_fp_val; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_fp_single; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_xcpt_pf_if; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_xcpt_ae_if; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_xcpt_ma_if; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_bp_debug_if; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_uop_bp_xcpt_if; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_brupdate_b2_uop_debug_fsrc; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_brupdate_b2_uop_debug_tsrc; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_valid; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_mispredict; // @[tile.scala 159:20]
  wire  core_io_ifu_brupdate_b2_taken; // @[tile.scala 159:20]
  wire [2:0] core_io_ifu_brupdate_b2_cfi_type; // @[tile.scala 159:20]
  wire [1:0] core_io_ifu_brupdate_b2_pc_sel; // @[tile.scala 159:20]
  wire [39:0] core_io_ifu_brupdate_b2_jalr_target; // @[tile.scala 159:20]
  wire [31:0] core_io_ifu_brupdate_b2_target_offset; // @[tile.scala 159:20]
  wire  core_io_ifu_redirect_flush; // @[tile.scala 159:20]
  wire  core_io_ifu_redirect_val; // @[tile.scala 159:20]
  wire [63:0] core_io_ifu_redirect_pc; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_redirect_ftq_idx; // @[tile.scala 159:20]
  wire [15:0] core_io_ifu_redirect_ghist_old_history; // @[tile.scala 159:20]
  wire  core_io_ifu_redirect_ghist_current_saw_branch_not_taken; // @[tile.scala 159:20]
  wire  core_io_ifu_redirect_ghist_new_saw_branch_not_taken; // @[tile.scala 159:20]
  wire  core_io_ifu_redirect_ghist_new_saw_branch_taken; // @[tile.scala 159:20]
  wire [4:0] core_io_ifu_redirect_ghist_ras_idx; // @[tile.scala 159:20]
  wire  core_io_ifu_commit_valid; // @[tile.scala 159:20]
  wire [31:0] core_io_ifu_commit_bits; // @[tile.scala 159:20]
  wire  core_io_ifu_flush_icache; // @[tile.scala 159:20]
  wire  core_io_ifu_perf_acquire; // @[tile.scala 159:20]
  wire  core_io_ifu_perf_tlbMiss; // @[tile.scala 159:20]
  wire  core_io_ifu_is_unicore; // @[tile.scala 159:20]
  wire [3:0] core_io_ptw_ptbr_mode; // @[tile.scala 159:20]
  wire [15:0] core_io_ptw_ptbr_asid; // @[tile.scala 159:20]
  wire [43:0] core_io_ptw_ptbr_ppn; // @[tile.scala 159:20]
  wire  core_io_ptw_sfence_valid; // @[tile.scala 159:20]
  wire  core_io_ptw_sfence_bits_rs1; // @[tile.scala 159:20]
  wire  core_io_ptw_sfence_bits_rs2; // @[tile.scala 159:20]
  wire [38:0] core_io_ptw_sfence_bits_addr; // @[tile.scala 159:20]
  wire  core_io_ptw_sfence_bits_asid; // @[tile.scala 159:20]
  wire  core_io_ptw_status_debug; // @[tile.scala 159:20]
  wire  core_io_ptw_status_cease; // @[tile.scala 159:20]
  wire  core_io_ptw_status_wfi; // @[tile.scala 159:20]
  wire [31:0] core_io_ptw_status_isa; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_status_dprv; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_status_prv; // @[tile.scala 159:20]
  wire  core_io_ptw_status_sd; // @[tile.scala 159:20]
  wire [26:0] core_io_ptw_status_zero2; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_status_sxl; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_status_uxl; // @[tile.scala 159:20]
  wire  core_io_ptw_status_sd_rv32; // @[tile.scala 159:20]
  wire [7:0] core_io_ptw_status_zero1; // @[tile.scala 159:20]
  wire  core_io_ptw_status_tsr; // @[tile.scala 159:20]
  wire  core_io_ptw_status_tw; // @[tile.scala 159:20]
  wire  core_io_ptw_status_tvm; // @[tile.scala 159:20]
  wire  core_io_ptw_status_mxr; // @[tile.scala 159:20]
  wire  core_io_ptw_status_sum; // @[tile.scala 159:20]
  wire  core_io_ptw_status_mprv; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_status_xs; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_status_fs; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_status_mpp; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_status_vs; // @[tile.scala 159:20]
  wire  core_io_ptw_status_spp; // @[tile.scala 159:20]
  wire  core_io_ptw_status_mpie; // @[tile.scala 159:20]
  wire  core_io_ptw_status_hpie; // @[tile.scala 159:20]
  wire  core_io_ptw_status_spie; // @[tile.scala 159:20]
  wire  core_io_ptw_status_upie; // @[tile.scala 159:20]
  wire  core_io_ptw_status_mie; // @[tile.scala 159:20]
  wire  core_io_ptw_status_hie; // @[tile.scala 159:20]
  wire  core_io_ptw_status_sie; // @[tile.scala 159:20]
  wire  core_io_ptw_status_uie; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_0_cfg_l; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_pmp_0_cfg_res; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_pmp_0_cfg_a; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_0_cfg_x; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_0_cfg_w; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_0_cfg_r; // @[tile.scala 159:20]
  wire [29:0] core_io_ptw_pmp_0_addr; // @[tile.scala 159:20]
  wire [31:0] core_io_ptw_pmp_0_mask; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_1_cfg_l; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_pmp_1_cfg_res; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_pmp_1_cfg_a; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_1_cfg_x; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_1_cfg_w; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_1_cfg_r; // @[tile.scala 159:20]
  wire [29:0] core_io_ptw_pmp_1_addr; // @[tile.scala 159:20]
  wire [31:0] core_io_ptw_pmp_1_mask; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_2_cfg_l; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_pmp_2_cfg_res; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_pmp_2_cfg_a; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_2_cfg_x; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_2_cfg_w; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_2_cfg_r; // @[tile.scala 159:20]
  wire [29:0] core_io_ptw_pmp_2_addr; // @[tile.scala 159:20]
  wire [31:0] core_io_ptw_pmp_2_mask; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_3_cfg_l; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_pmp_3_cfg_res; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_pmp_3_cfg_a; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_3_cfg_x; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_3_cfg_w; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_3_cfg_r; // @[tile.scala 159:20]
  wire [29:0] core_io_ptw_pmp_3_addr; // @[tile.scala 159:20]
  wire [31:0] core_io_ptw_pmp_3_mask; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_4_cfg_l; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_pmp_4_cfg_res; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_pmp_4_cfg_a; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_4_cfg_x; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_4_cfg_w; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_4_cfg_r; // @[tile.scala 159:20]
  wire [29:0] core_io_ptw_pmp_4_addr; // @[tile.scala 159:20]
  wire [31:0] core_io_ptw_pmp_4_mask; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_5_cfg_l; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_pmp_5_cfg_res; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_pmp_5_cfg_a; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_5_cfg_x; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_5_cfg_w; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_5_cfg_r; // @[tile.scala 159:20]
  wire [29:0] core_io_ptw_pmp_5_addr; // @[tile.scala 159:20]
  wire [31:0] core_io_ptw_pmp_5_mask; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_6_cfg_l; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_pmp_6_cfg_res; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_pmp_6_cfg_a; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_6_cfg_x; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_6_cfg_w; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_6_cfg_r; // @[tile.scala 159:20]
  wire [29:0] core_io_ptw_pmp_6_addr; // @[tile.scala 159:20]
  wire [31:0] core_io_ptw_pmp_6_mask; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_7_cfg_l; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_pmp_7_cfg_res; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_pmp_7_cfg_a; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_7_cfg_x; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_7_cfg_w; // @[tile.scala 159:20]
  wire  core_io_ptw_pmp_7_cfg_r; // @[tile.scala 159:20]
  wire [29:0] core_io_ptw_pmp_7_addr; // @[tile.scala 159:20]
  wire [31:0] core_io_ptw_pmp_7_mask; // @[tile.scala 159:20]
  wire  core_io_ptw_perf_l2miss; // @[tile.scala 159:20]
  wire  core_io_ptw_perf_l2hit; // @[tile.scala 159:20]
  wire  core_io_ptw_perf_pte_miss; // @[tile.scala 159:20]
  wire  core_io_ptw_perf_pte_hit; // @[tile.scala 159:20]
  wire  core_io_ptw_customCSRs_csrs_0_wen; // @[tile.scala 159:20]
  wire [63:0] core_io_ptw_customCSRs_csrs_0_wdata; // @[tile.scala 159:20]
  wire [63:0] core_io_ptw_customCSRs_csrs_0_value; // @[tile.scala 159:20]
  wire  core_io_ptw_clock_enabled; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_ready; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_valid; // @[tile.scala 159:20]
  wire [6:0] core_io_rocc_cmd_bits_inst_funct; // @[tile.scala 159:20]
  wire [4:0] core_io_rocc_cmd_bits_inst_rs2; // @[tile.scala 159:20]
  wire [4:0] core_io_rocc_cmd_bits_inst_rs1; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_inst_xd; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_inst_xs1; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_inst_xs2; // @[tile.scala 159:20]
  wire [4:0] core_io_rocc_cmd_bits_inst_rd; // @[tile.scala 159:20]
  wire [6:0] core_io_rocc_cmd_bits_inst_opcode; // @[tile.scala 159:20]
  wire [63:0] core_io_rocc_cmd_bits_rs1; // @[tile.scala 159:20]
  wire [63:0] core_io_rocc_cmd_bits_rs2; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_status_debug; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_status_cease; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_status_wfi; // @[tile.scala 159:20]
  wire [31:0] core_io_rocc_cmd_bits_status_isa; // @[tile.scala 159:20]
  wire [1:0] core_io_rocc_cmd_bits_status_dprv; // @[tile.scala 159:20]
  wire [1:0] core_io_rocc_cmd_bits_status_prv; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_status_sd; // @[tile.scala 159:20]
  wire [26:0] core_io_rocc_cmd_bits_status_zero2; // @[tile.scala 159:20]
  wire [1:0] core_io_rocc_cmd_bits_status_sxl; // @[tile.scala 159:20]
  wire [1:0] core_io_rocc_cmd_bits_status_uxl; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_status_sd_rv32; // @[tile.scala 159:20]
  wire [7:0] core_io_rocc_cmd_bits_status_zero1; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_status_tsr; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_status_tw; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_status_tvm; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_status_mxr; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_status_sum; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_status_mprv; // @[tile.scala 159:20]
  wire [1:0] core_io_rocc_cmd_bits_status_xs; // @[tile.scala 159:20]
  wire [1:0] core_io_rocc_cmd_bits_status_fs; // @[tile.scala 159:20]
  wire [1:0] core_io_rocc_cmd_bits_status_mpp; // @[tile.scala 159:20]
  wire [1:0] core_io_rocc_cmd_bits_status_vs; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_status_spp; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_status_mpie; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_status_hpie; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_status_spie; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_status_upie; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_status_mie; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_status_hie; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_status_sie; // @[tile.scala 159:20]
  wire  core_io_rocc_cmd_bits_status_uie; // @[tile.scala 159:20]
  wire  core_io_rocc_resp_ready; // @[tile.scala 159:20]
  wire  core_io_rocc_resp_valid; // @[tile.scala 159:20]
  wire [4:0] core_io_rocc_resp_bits_rd; // @[tile.scala 159:20]
  wire [63:0] core_io_rocc_resp_bits_data; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_req_ready; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_req_valid; // @[tile.scala 159:20]
  wire [39:0] core_io_rocc_mem_req_bits_addr; // @[tile.scala 159:20]
  wire [6:0] core_io_rocc_mem_req_bits_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_rocc_mem_req_bits_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_rocc_mem_req_bits_size; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_req_bits_signed; // @[tile.scala 159:20]
  wire [1:0] core_io_rocc_mem_req_bits_dprv; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_req_bits_phys; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_req_bits_no_alloc; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_req_bits_no_xcpt; // @[tile.scala 159:20]
  wire [63:0] core_io_rocc_mem_req_bits_data; // @[tile.scala 159:20]
  wire [7:0] core_io_rocc_mem_req_bits_mask; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_s1_kill; // @[tile.scala 159:20]
  wire [63:0] core_io_rocc_mem_s1_data_data; // @[tile.scala 159:20]
  wire [7:0] core_io_rocc_mem_s1_data_mask; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_s2_nack; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_s2_nack_cause_raw; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_s2_kill; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_s2_uncached; // @[tile.scala 159:20]
  wire [31:0] core_io_rocc_mem_s2_paddr; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_resp_valid; // @[tile.scala 159:20]
  wire [39:0] core_io_rocc_mem_resp_bits_addr; // @[tile.scala 159:20]
  wire [6:0] core_io_rocc_mem_resp_bits_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_rocc_mem_resp_bits_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_rocc_mem_resp_bits_size; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_resp_bits_signed; // @[tile.scala 159:20]
  wire [1:0] core_io_rocc_mem_resp_bits_dprv; // @[tile.scala 159:20]
  wire [63:0] core_io_rocc_mem_resp_bits_data; // @[tile.scala 159:20]
  wire [7:0] core_io_rocc_mem_resp_bits_mask; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_resp_bits_replay; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_resp_bits_has_data; // @[tile.scala 159:20]
  wire [63:0] core_io_rocc_mem_resp_bits_data_word_bypass; // @[tile.scala 159:20]
  wire [63:0] core_io_rocc_mem_resp_bits_data_raw; // @[tile.scala 159:20]
  wire [63:0] core_io_rocc_mem_resp_bits_store_data; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_replay_next; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_s2_xcpt_ma_ld; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_s2_xcpt_ma_st; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_s2_xcpt_pf_ld; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_s2_xcpt_pf_st; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_s2_xcpt_ae_ld; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_s2_xcpt_ae_st; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_ordered; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_perf_acquire; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_perf_release; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_perf_grant; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_perf_tlbMiss; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_perf_blocked; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_perf_canAcceptStoreThenLoad; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_perf_canAcceptStoreThenRMW; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_perf_canAcceptLoadThenLoad; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_perf_storeBufferEmptyAfterLoad; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_perf_storeBufferEmptyAfterStore; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_keep_clock_enabled; // @[tile.scala 159:20]
  wire  core_io_rocc_mem_clock_enabled; // @[tile.scala 159:20]
  wire  core_io_rocc_busy; // @[tile.scala 159:20]
  wire  core_io_rocc_interrupt; // @[tile.scala 159:20]
  wire  core_io_rocc_exception; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_valid; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_switch; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_switch_off; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_is_unicore; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_req_bits_uop_shift; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_uop_lrs3_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_rflag; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_wflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_uop_prflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_uop_pwflag; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_pflag_busy; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_uop_stale_pflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_uop_op1_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_uop_op2_sel; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_uop_split_num; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_uop_self_index; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_uop_rob_inst_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_uop_address_num; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_req_bits_uop_uopc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_exe_0_req_bits_uop_inst; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_exe_0_req_bits_uop_debug_inst; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_is_rvc; // @[tile.scala 159:20]
  wire [39:0] core_io_lsu_exe_0_req_bits_uop_debug_pc; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_req_bits_uop_iq_type; // @[tile.scala 159:20]
  wire [9:0] core_io_lsu_exe_0_req_bits_uop_fu_code; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_uop_ctrl_br_type; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_uop_ctrl_op1_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_req_bits_uop_ctrl_op2_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_req_bits_uop_ctrl_imm_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_uop_ctrl_op_fcn; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_ctrl_fcn_dw; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_req_bits_uop_ctrl_csr_cmd; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_ctrl_is_load; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_ctrl_is_sta; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_ctrl_is_std; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_uop_ctrl_op3_sel; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_uop_iw_state; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_iw_p1_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_iw_p2_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_is_br; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_is_jalr; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_is_jal; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_is_sfb; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_exe_0_req_bits_uop_br_mask; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_uop_br_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_req_bits_uop_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_edge_inst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_uop_pc_lob; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_taken; // @[tile.scala 159:20]
  wire [19:0] core_io_lsu_exe_0_req_bits_uop_imm_packed; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_exe_0_req_bits_uop_csr_addr; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_uop_rob_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_req_bits_uop_ldq_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_req_bits_uop_stq_idx; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_uop_rxq_idx; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_req_bits_uop_pdst; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_req_bits_uop_prs1; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_req_bits_uop_prs2; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_req_bits_uop_prs3; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_req_bits_uop_ppred; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_prs1_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_prs2_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_prs3_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_ppred_busy; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_req_bits_uop_stale_pdst; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_exception; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_exe_0_req_bits_uop_exc_cause; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_bypassable; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_req_bits_uop_mem_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_uop_mem_size; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_mem_signed; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_is_fence; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_is_fencei; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_is_amo; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_uses_ldq; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_uses_stq; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_is_sys_pc2epc; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_is_unique; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_flush_on_commit; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_ldst_is_rs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_uop_ldst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_uop_lrs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_uop_lrs2; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_uop_lrs3; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_ldst_val; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_uop_dst_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_uop_lrs1_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_uop_lrs2_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_frs3_en; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_fp_val; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_fp_single; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_xcpt_pf_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_xcpt_ae_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_xcpt_ma_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_bp_debug_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_uop_bp_xcpt_if; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_uop_debug_fsrc; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_uop_debug_tsrc; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_predicated; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_exe_0_req_bits_data; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_valid; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_switch; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_switch_off; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_unicore; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_shift; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_lrs3_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_rflag; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_wflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_prflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_pwflag; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_pflag_busy; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_stale_pflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_op1_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_op2_sel; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_split_num; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_self_index; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_rob_inst_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_address_num; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_uopc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_inst; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_debug_inst; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_rvc; // @[tile.scala 159:20]
  wire [39:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_debug_pc; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_iq_type; // @[tile.scala 159:20]
  wire [9:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_fu_code; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_br_type; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_op1_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_op2_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_imm_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_op_fcn; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_fcn_dw; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_csr_cmd; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_is_load; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_is_sta; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_is_std; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_op3_sel; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_iw_state; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_iw_p1_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_iw_p2_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_br; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_jalr; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_jal; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_sfb; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_br_mask; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_br_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_edge_inst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_pc_lob; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_taken; // @[tile.scala 159:20]
  wire [19:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_imm_packed; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_csr_addr; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_rob_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_ldq_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_stq_idx; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_rxq_idx; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_pdst; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_prs1; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_prs2; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_prs3; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_ppred; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_prs1_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_prs2_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_prs3_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_ppred_busy; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_stale_pdst; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_exception; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_exc_cause; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_bypassable; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_mem_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_mem_size; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_mem_signed; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_fence; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_fencei; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_amo; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_uses_ldq; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_uses_stq; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_sys_pc2epc; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_unique; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_flush_on_commit; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_ldst_is_rs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_ldst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_lrs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_lrs2; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_lrs3; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_ldst_val; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_dst_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_lrs1_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_lrs2_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_frs3_en; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_fp_val; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_fp_single; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_xcpt_pf_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_xcpt_ae_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_xcpt_ma_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_bp_debug_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflags_bits_uop_bp_xcpt_if; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_debug_fsrc; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflags_bits_uop_debug_tsrc; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_req_bits_fflags_bits_flags; // @[tile.scala 159:20]
  wire [39:0] core_io_lsu_exe_0_req_bits_addr; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_mxcpt_valid; // @[tile.scala 159:20]
  wire [16:0] core_io_lsu_exe_0_req_bits_mxcpt_bits; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_sfence_valid; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_sfence_bits_rs1; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_sfence_bits_rs2; // @[tile.scala 159:20]
  wire [38:0] core_io_lsu_exe_0_req_bits_sfence_bits_addr; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_sfence_bits_asid; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_flagdata; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_valid; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_switch; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_switch_off; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_unicore; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_shift; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs3_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_rflag; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_wflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_prflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_pwflag; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_pflag_busy; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_stale_pflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_op1_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_op2_sel; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_split_num; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_self_index; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_rob_inst_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_address_num; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_uopc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_inst; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_debug_inst; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_rvc; // @[tile.scala 159:20]
  wire [39:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_debug_pc; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_iq_type; // @[tile.scala 159:20]
  wire [9:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_fu_code; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_br_type; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_op1_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_op2_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_imm_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_op_fcn; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_fcn_dw; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_csr_cmd; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_load; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_sta; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_std; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_op3_sel; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_iw_state; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_iw_p1_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_iw_p2_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_br; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_jalr; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_jal; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_sfb; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_br_mask; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_br_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_edge_inst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_pc_lob; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_taken; // @[tile.scala 159:20]
  wire [19:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_imm_packed; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_csr_addr; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_rob_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ldq_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_stq_idx; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_rxq_idx; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_pdst; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs1; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs2; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs3; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ppred; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs1_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs2_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs3_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ppred_busy; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_stale_pdst; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_exception; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_exc_cause; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_bypassable; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_mem_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_mem_size; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_mem_signed; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_fence; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_fencei; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_amo; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_uses_ldq; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_uses_stq; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_sys_pc2epc; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_unique; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_flush_on_commit; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ldst_is_rs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ldst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs2; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs3; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ldst_val; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_dst_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs1_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs2_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_frs3_en; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_fp_val; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_fp_single; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_xcpt_pf_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_xcpt_ae_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_xcpt_ma_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_bp_debug_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_bp_xcpt_if; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_debug_fsrc; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_debug_tsrc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_exe_0_req_bits_fflagdata_bits_fflag; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_ready; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_valid; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_switch; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_switch_off; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_is_unicore; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_iresp_bits_uop_shift; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_uop_lrs3_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_rflag; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_wflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_uop_prflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_uop_pwflag; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_pflag_busy; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_uop_stale_pflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_uop_op1_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_uop_op2_sel; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_uop_split_num; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_uop_self_index; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_uop_rob_inst_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_uop_address_num; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_iresp_bits_uop_uopc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_exe_0_iresp_bits_uop_inst; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_exe_0_iresp_bits_uop_debug_inst; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_is_rvc; // @[tile.scala 159:20]
  wire [39:0] core_io_lsu_exe_0_iresp_bits_uop_debug_pc; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_iresp_bits_uop_iq_type; // @[tile.scala 159:20]
  wire [9:0] core_io_lsu_exe_0_iresp_bits_uop_fu_code; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_uop_ctrl_br_type; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_uop_ctrl_op1_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_iresp_bits_uop_ctrl_op2_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_iresp_bits_uop_ctrl_imm_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_uop_ctrl_op_fcn; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_ctrl_fcn_dw; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_iresp_bits_uop_ctrl_csr_cmd; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_ctrl_is_load; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_ctrl_is_sta; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_ctrl_is_std; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_uop_ctrl_op3_sel; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_uop_iw_state; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_iw_p1_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_iw_p2_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_is_br; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_is_jalr; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_is_jal; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_is_sfb; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_exe_0_iresp_bits_uop_br_mask; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_uop_br_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_iresp_bits_uop_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_edge_inst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_uop_pc_lob; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_taken; // @[tile.scala 159:20]
  wire [19:0] core_io_lsu_exe_0_iresp_bits_uop_imm_packed; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_exe_0_iresp_bits_uop_csr_addr; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_uop_rob_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_iresp_bits_uop_ldq_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_iresp_bits_uop_stq_idx; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_uop_rxq_idx; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_iresp_bits_uop_pdst; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_iresp_bits_uop_prs1; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_iresp_bits_uop_prs2; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_iresp_bits_uop_prs3; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_iresp_bits_uop_ppred; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_prs1_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_prs2_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_prs3_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_ppred_busy; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_iresp_bits_uop_stale_pdst; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_exception; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_exe_0_iresp_bits_uop_exc_cause; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_bypassable; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_iresp_bits_uop_mem_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_uop_mem_size; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_mem_signed; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_is_fence; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_is_fencei; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_is_amo; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_uses_ldq; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_uses_stq; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_is_sys_pc2epc; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_is_unique; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_flush_on_commit; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_ldst_is_rs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_uop_ldst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_uop_lrs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_uop_lrs2; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_uop_lrs3; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_ldst_val; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_uop_dst_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_uop_lrs1_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_uop_lrs2_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_frs3_en; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_fp_val; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_fp_single; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_xcpt_pf_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_xcpt_ae_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_xcpt_ma_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_bp_debug_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_uop_bp_xcpt_if; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_uop_debug_fsrc; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_uop_debug_tsrc; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_exe_0_iresp_bits_data; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_predicated; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_valid; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_switch; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_switch_off; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_unicore; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_shift; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs3_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_rflag; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_wflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_prflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_pwflag; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_pflag_busy; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_stale_pflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_op1_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_op2_sel; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_split_num; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_self_index; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_rob_inst_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_address_num; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_uopc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_inst; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_debug_inst; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_rvc; // @[tile.scala 159:20]
  wire [39:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_debug_pc; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_iq_type; // @[tile.scala 159:20]
  wire [9:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_fu_code; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_br_type; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_op1_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_op2_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_imm_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_op_fcn; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_fcn_dw; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_csr_cmd; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_load; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_sta; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_std; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_op3_sel; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_iw_state; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_iw_p1_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_iw_p2_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_br; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_jalr; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_jal; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_sfb; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_br_mask; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_br_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_edge_inst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_pc_lob; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_taken; // @[tile.scala 159:20]
  wire [19:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_imm_packed; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_csr_addr; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_rob_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ldq_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_stq_idx; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_rxq_idx; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_pdst; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs1; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs2; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs3; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ppred; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs1_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs2_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs3_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ppred_busy; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_stale_pdst; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_exception; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_exc_cause; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_bypassable; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_mem_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_mem_size; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_mem_signed; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_fence; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_fencei; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_amo; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_uses_ldq; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_uses_stq; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_sys_pc2epc; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_unique; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_flush_on_commit; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ldst_is_rs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ldst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs2; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs3; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ldst_val; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_dst_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs1_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs2_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_frs3_en; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_fp_val; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_fp_single; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_xcpt_pf_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_xcpt_ae_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_xcpt_ma_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_bp_debug_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_bp_xcpt_if; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_debug_fsrc; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_debug_tsrc; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_iresp_bits_fflags_bits_flags; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_flagdata; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_valid; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_switch; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_switch_off; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_unicore; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_shift; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs3_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_rflag; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_wflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_pwflag; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_pflag_busy; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_stale_pflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_op1_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_op2_sel; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_split_num; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_self_index; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_rob_inst_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_address_num; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_uopc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_inst; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_debug_inst; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_rvc; // @[tile.scala 159:20]
  wire [39:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_debug_pc; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_iq_type; // @[tile.scala 159:20]
  wire [9:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_fu_code; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_br_type; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op1_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op2_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_imm_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op_fcn; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_fcn_dw; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_csr_cmd; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_load; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_sta; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_std; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op3_sel; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_iw_state; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_iw_p1_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_iw_p2_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_br; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_jalr; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_jal; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_sfb; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_br_mask; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_br_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_edge_inst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_pc_lob; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_taken; // @[tile.scala 159:20]
  wire [19:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_imm_packed; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_csr_addr; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_rob_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ldq_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_stq_idx; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_rxq_idx; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_pdst; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs1; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs2; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs3; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ppred; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs1_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs2_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs3_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ppred_busy; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_stale_pdst; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_exception; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_exc_cause; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_bypassable; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_mem_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_mem_size; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_mem_signed; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_fence; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_fencei; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_amo; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_uses_ldq; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_uses_stq; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_sys_pc2epc; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_unique; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_flush_on_commit; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ldst_is_rs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ldst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs2; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs3; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ldst_val; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_dst_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs1_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs2_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_frs3_en; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_fp_val; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_fp_single; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_pf_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_ae_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_ma_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_bp_debug_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_bp_xcpt_if; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_debug_fsrc; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_debug_tsrc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_exe_0_iresp_bits_fflagdata_bits_fflag; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_ready; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_valid; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_switch; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_switch_off; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_is_unicore; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_fresp_bits_uop_shift; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_uop_lrs3_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_rflag; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_wflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_uop_prflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_uop_pwflag; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_pflag_busy; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_uop_stale_pflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_uop_op1_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_uop_op2_sel; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_uop_split_num; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_uop_self_index; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_uop_rob_inst_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_uop_address_num; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_fresp_bits_uop_uopc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_exe_0_fresp_bits_uop_inst; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_exe_0_fresp_bits_uop_debug_inst; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_is_rvc; // @[tile.scala 159:20]
  wire [39:0] core_io_lsu_exe_0_fresp_bits_uop_debug_pc; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_fresp_bits_uop_iq_type; // @[tile.scala 159:20]
  wire [9:0] core_io_lsu_exe_0_fresp_bits_uop_fu_code; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_uop_ctrl_br_type; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_uop_ctrl_op1_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_fresp_bits_uop_ctrl_op2_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_fresp_bits_uop_ctrl_imm_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_uop_ctrl_op_fcn; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_ctrl_fcn_dw; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_fresp_bits_uop_ctrl_csr_cmd; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_ctrl_is_load; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_ctrl_is_sta; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_ctrl_is_std; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_uop_ctrl_op3_sel; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_uop_iw_state; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_iw_p1_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_iw_p2_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_is_br; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_is_jalr; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_is_jal; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_is_sfb; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_exe_0_fresp_bits_uop_br_mask; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_uop_br_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_fresp_bits_uop_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_edge_inst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_uop_pc_lob; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_taken; // @[tile.scala 159:20]
  wire [19:0] core_io_lsu_exe_0_fresp_bits_uop_imm_packed; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_exe_0_fresp_bits_uop_csr_addr; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_uop_rob_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_fresp_bits_uop_ldq_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_fresp_bits_uop_stq_idx; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_uop_rxq_idx; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_fresp_bits_uop_pdst; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_fresp_bits_uop_prs1; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_fresp_bits_uop_prs2; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_fresp_bits_uop_prs3; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_fresp_bits_uop_ppred; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_prs1_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_prs2_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_prs3_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_ppred_busy; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_fresp_bits_uop_stale_pdst; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_exception; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_exe_0_fresp_bits_uop_exc_cause; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_bypassable; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_fresp_bits_uop_mem_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_uop_mem_size; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_mem_signed; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_is_fence; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_is_fencei; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_is_amo; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_uses_ldq; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_uses_stq; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_is_sys_pc2epc; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_is_unique; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_flush_on_commit; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_ldst_is_rs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_uop_ldst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_uop_lrs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_uop_lrs2; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_uop_lrs3; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_ldst_val; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_uop_dst_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_uop_lrs1_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_uop_lrs2_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_frs3_en; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_fp_val; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_fp_single; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_xcpt_pf_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_xcpt_ae_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_xcpt_ma_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_bp_debug_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_uop_bp_xcpt_if; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_uop_debug_fsrc; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_uop_debug_tsrc; // @[tile.scala 159:20]
  wire [64:0] core_io_lsu_exe_0_fresp_bits_data; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_predicated; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_valid; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_switch; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_switch_off; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_unicore; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_shift; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs3_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_rflag; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_wflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_prflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_pwflag; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_pflag_busy; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_stale_pflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_op1_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_op2_sel; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_split_num; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_self_index; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_rob_inst_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_address_num; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_uopc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_inst; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_debug_inst; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_rvc; // @[tile.scala 159:20]
  wire [39:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_debug_pc; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_iq_type; // @[tile.scala 159:20]
  wire [9:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_fu_code; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_br_type; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_op1_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_op2_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_imm_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_op_fcn; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_fcn_dw; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_csr_cmd; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_load; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_sta; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_std; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_op3_sel; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_iw_state; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_iw_p1_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_iw_p2_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_br; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_jalr; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_jal; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_sfb; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_br_mask; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_br_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_edge_inst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_pc_lob; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_taken; // @[tile.scala 159:20]
  wire [19:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_imm_packed; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_csr_addr; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_rob_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ldq_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_stq_idx; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_rxq_idx; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_pdst; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs1; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs2; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs3; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ppred; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs1_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs2_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs3_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ppred_busy; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_stale_pdst; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_exception; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_exc_cause; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_bypassable; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_mem_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_mem_size; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_mem_signed; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_fence; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_fencei; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_amo; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_uses_ldq; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_uses_stq; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_sys_pc2epc; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_unique; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_flush_on_commit; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ldst_is_rs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ldst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs2; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs3; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ldst_val; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_dst_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs1_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs2_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_frs3_en; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_fp_val; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_fp_single; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_xcpt_pf_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_xcpt_ae_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_xcpt_ma_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_bp_debug_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_bp_xcpt_if; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_debug_fsrc; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_debug_tsrc; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_fresp_bits_fflags_bits_flags; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_flagdata; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_valid; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_switch; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_switch_off; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_unicore; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_shift; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs3_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_rflag; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_wflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_pwflag; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_pflag_busy; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_stale_pflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_op1_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_op2_sel; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_split_num; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_self_index; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_rob_inst_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_address_num; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_uopc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_inst; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_debug_inst; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_rvc; // @[tile.scala 159:20]
  wire [39:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_debug_pc; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_iq_type; // @[tile.scala 159:20]
  wire [9:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_fu_code; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_br_type; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op1_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op2_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_imm_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op_fcn; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_fcn_dw; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_csr_cmd; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_load; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_sta; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_std; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op3_sel; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_iw_state; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_iw_p1_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_iw_p2_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_br; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_jalr; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_jal; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_sfb; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_br_mask; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_br_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_edge_inst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_pc_lob; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_taken; // @[tile.scala 159:20]
  wire [19:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_imm_packed; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_csr_addr; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_rob_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ldq_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_stq_idx; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_rxq_idx; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_pdst; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs1; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs2; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs3; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ppred; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs1_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs2_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs3_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ppred_busy; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_stale_pdst; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_exception; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_exc_cause; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_bypassable; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_mem_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_mem_size; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_mem_signed; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_fence; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_fencei; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_amo; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_uses_ldq; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_uses_stq; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_sys_pc2epc; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_unique; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_flush_on_commit; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ldst_is_rs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ldst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs2; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs3; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ldst_val; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_dst_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs1_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs2_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_frs3_en; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_fp_val; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_fp_single; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_pf_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_ae_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_ma_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_bp_debug_if; // @[tile.scala 159:20]
  wire  core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_bp_xcpt_if; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_debug_fsrc; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_debug_tsrc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_exe_0_fresp_bits_fflagdata_bits_fflag; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_valid; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_switch; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_switch_off; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_is_unicore; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_dis_uops_0_bits_shift; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_0_bits_lrs3_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_rflag; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_wflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_dis_uops_0_bits_prflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_dis_uops_0_bits_pwflag; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_pflag_busy; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_dis_uops_0_bits_stale_pflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_dis_uops_0_bits_op1_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_dis_uops_0_bits_op2_sel; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_dis_uops_0_bits_split_num; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_dis_uops_0_bits_self_index; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_dis_uops_0_bits_rob_inst_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_dis_uops_0_bits_address_num; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_dis_uops_0_bits_uopc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_dis_uops_0_bits_inst; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_dis_uops_0_bits_debug_inst; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_is_rvc; // @[tile.scala 159:20]
  wire [39:0] core_io_lsu_dis_uops_0_bits_debug_pc; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_dis_uops_0_bits_iq_type; // @[tile.scala 159:20]
  wire [9:0] core_io_lsu_dis_uops_0_bits_fu_code; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_dis_uops_0_bits_ctrl_br_type; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_0_bits_ctrl_op1_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_dis_uops_0_bits_ctrl_op2_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_dis_uops_0_bits_ctrl_imm_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_dis_uops_0_bits_ctrl_op_fcn; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_ctrl_fcn_dw; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_dis_uops_0_bits_ctrl_csr_cmd; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_ctrl_is_load; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_ctrl_is_sta; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_ctrl_is_std; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_0_bits_ctrl_op3_sel; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_0_bits_iw_state; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_iw_p1_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_iw_p2_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_is_br; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_is_jalr; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_is_jal; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_is_sfb; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_dis_uops_0_bits_br_mask; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_dis_uops_0_bits_br_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_dis_uops_0_bits_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_edge_inst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_dis_uops_0_bits_pc_lob; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_taken; // @[tile.scala 159:20]
  wire [19:0] core_io_lsu_dis_uops_0_bits_imm_packed; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_dis_uops_0_bits_csr_addr; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_dis_uops_0_bits_rob_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_dis_uops_0_bits_ldq_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_dis_uops_0_bits_stq_idx; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_0_bits_rxq_idx; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_dis_uops_0_bits_pdst; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_dis_uops_0_bits_prs1; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_dis_uops_0_bits_prs2; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_dis_uops_0_bits_prs3; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_dis_uops_0_bits_ppred; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_prs1_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_prs2_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_prs3_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_ppred_busy; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_dis_uops_0_bits_stale_pdst; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_exception; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_dis_uops_0_bits_exc_cause; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_bypassable; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_dis_uops_0_bits_mem_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_0_bits_mem_size; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_mem_signed; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_is_fence; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_is_fencei; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_is_amo; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_uses_ldq; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_uses_stq; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_is_sys_pc2epc; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_is_unique; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_flush_on_commit; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_ldst_is_rs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_dis_uops_0_bits_ldst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_dis_uops_0_bits_lrs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_dis_uops_0_bits_lrs2; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_dis_uops_0_bits_lrs3; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_ldst_val; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_0_bits_dst_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_0_bits_lrs1_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_0_bits_lrs2_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_frs3_en; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_fp_val; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_fp_single; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_xcpt_pf_if; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_xcpt_ae_if; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_xcpt_ma_if; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_bp_debug_if; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_0_bits_bp_xcpt_if; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_0_bits_debug_fsrc; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_0_bits_debug_tsrc; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_valid; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_switch; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_switch_off; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_is_unicore; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_dis_uops_1_bits_shift; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_1_bits_lrs3_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_rflag; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_wflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_dis_uops_1_bits_prflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_dis_uops_1_bits_pwflag; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_pflag_busy; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_dis_uops_1_bits_stale_pflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_dis_uops_1_bits_op1_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_dis_uops_1_bits_op2_sel; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_dis_uops_1_bits_split_num; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_dis_uops_1_bits_self_index; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_dis_uops_1_bits_rob_inst_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_dis_uops_1_bits_address_num; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_dis_uops_1_bits_uopc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_dis_uops_1_bits_inst; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_dis_uops_1_bits_debug_inst; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_is_rvc; // @[tile.scala 159:20]
  wire [39:0] core_io_lsu_dis_uops_1_bits_debug_pc; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_dis_uops_1_bits_iq_type; // @[tile.scala 159:20]
  wire [9:0] core_io_lsu_dis_uops_1_bits_fu_code; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_dis_uops_1_bits_ctrl_br_type; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_1_bits_ctrl_op1_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_dis_uops_1_bits_ctrl_op2_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_dis_uops_1_bits_ctrl_imm_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_dis_uops_1_bits_ctrl_op_fcn; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_ctrl_fcn_dw; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_dis_uops_1_bits_ctrl_csr_cmd; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_ctrl_is_load; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_ctrl_is_sta; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_ctrl_is_std; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_1_bits_ctrl_op3_sel; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_1_bits_iw_state; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_iw_p1_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_iw_p2_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_is_br; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_is_jalr; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_is_jal; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_is_sfb; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_dis_uops_1_bits_br_mask; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_dis_uops_1_bits_br_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_dis_uops_1_bits_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_edge_inst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_dis_uops_1_bits_pc_lob; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_taken; // @[tile.scala 159:20]
  wire [19:0] core_io_lsu_dis_uops_1_bits_imm_packed; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_dis_uops_1_bits_csr_addr; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_dis_uops_1_bits_rob_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_dis_uops_1_bits_ldq_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_dis_uops_1_bits_stq_idx; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_1_bits_rxq_idx; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_dis_uops_1_bits_pdst; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_dis_uops_1_bits_prs1; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_dis_uops_1_bits_prs2; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_dis_uops_1_bits_prs3; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_dis_uops_1_bits_ppred; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_prs1_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_prs2_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_prs3_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_ppred_busy; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_dis_uops_1_bits_stale_pdst; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_exception; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_dis_uops_1_bits_exc_cause; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_bypassable; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_dis_uops_1_bits_mem_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_1_bits_mem_size; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_mem_signed; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_is_fence; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_is_fencei; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_is_amo; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_uses_ldq; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_uses_stq; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_is_sys_pc2epc; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_is_unique; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_flush_on_commit; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_ldst_is_rs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_dis_uops_1_bits_ldst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_dis_uops_1_bits_lrs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_dis_uops_1_bits_lrs2; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_dis_uops_1_bits_lrs3; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_ldst_val; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_1_bits_dst_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_1_bits_lrs1_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_1_bits_lrs2_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_frs3_en; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_fp_val; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_fp_single; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_xcpt_pf_if; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_xcpt_ae_if; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_xcpt_ma_if; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_bp_debug_if; // @[tile.scala 159:20]
  wire  core_io_lsu_dis_uops_1_bits_bp_xcpt_if; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_1_bits_debug_fsrc; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_dis_uops_1_bits_debug_tsrc; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_dis_ldq_idx_0; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_dis_ldq_idx_1; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_dis_stq_idx_0; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_dis_stq_idx_1; // @[tile.scala 159:20]
  wire  core_io_lsu_ldq_full_0; // @[tile.scala 159:20]
  wire  core_io_lsu_ldq_full_1; // @[tile.scala 159:20]
  wire  core_io_lsu_stq_full_0; // @[tile.scala 159:20]
  wire  core_io_lsu_stq_full_1; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_ready; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_valid; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_switch; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_switch_off; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_is_unicore; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_fp_stdata_bits_uop_shift; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_uop_lrs3_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_rflag; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_wflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_uop_prflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_uop_pwflag; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_pflag_busy; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_uop_stale_pflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_uop_op1_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_uop_op2_sel; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_uop_split_num; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_uop_self_index; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_uop_rob_inst_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_uop_address_num; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_fp_stdata_bits_uop_uopc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_fp_stdata_bits_uop_inst; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_fp_stdata_bits_uop_debug_inst; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_is_rvc; // @[tile.scala 159:20]
  wire [39:0] core_io_lsu_fp_stdata_bits_uop_debug_pc; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_fp_stdata_bits_uop_iq_type; // @[tile.scala 159:20]
  wire [9:0] core_io_lsu_fp_stdata_bits_uop_fu_code; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_uop_ctrl_br_type; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_uop_ctrl_op1_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_fp_stdata_bits_uop_ctrl_op2_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_fp_stdata_bits_uop_ctrl_imm_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_uop_ctrl_op_fcn; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_ctrl_fcn_dw; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_fp_stdata_bits_uop_ctrl_csr_cmd; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_ctrl_is_load; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_ctrl_is_sta; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_ctrl_is_std; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_uop_ctrl_op3_sel; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_uop_iw_state; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_iw_p1_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_iw_p2_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_is_br; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_is_jalr; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_is_jal; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_is_sfb; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_fp_stdata_bits_uop_br_mask; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_uop_br_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_fp_stdata_bits_uop_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_edge_inst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_uop_pc_lob; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_taken; // @[tile.scala 159:20]
  wire [19:0] core_io_lsu_fp_stdata_bits_uop_imm_packed; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_fp_stdata_bits_uop_csr_addr; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_uop_rob_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_fp_stdata_bits_uop_ldq_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_fp_stdata_bits_uop_stq_idx; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_uop_rxq_idx; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_fp_stdata_bits_uop_pdst; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_fp_stdata_bits_uop_prs1; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_fp_stdata_bits_uop_prs2; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_fp_stdata_bits_uop_prs3; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_fp_stdata_bits_uop_ppred; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_prs1_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_prs2_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_prs3_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_ppred_busy; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_fp_stdata_bits_uop_stale_pdst; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_exception; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_fp_stdata_bits_uop_exc_cause; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_bypassable; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_fp_stdata_bits_uop_mem_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_uop_mem_size; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_mem_signed; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_is_fence; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_is_fencei; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_is_amo; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_uses_ldq; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_uses_stq; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_is_sys_pc2epc; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_is_unique; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_flush_on_commit; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_ldst_is_rs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_uop_ldst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_uop_lrs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_uop_lrs2; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_uop_lrs3; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_ldst_val; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_uop_dst_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_uop_lrs1_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_uop_lrs2_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_frs3_en; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_fp_val; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_fp_single; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_xcpt_pf_if; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_xcpt_ae_if; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_xcpt_ma_if; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_bp_debug_if; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_uop_bp_xcpt_if; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_uop_debug_fsrc; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_uop_debug_tsrc; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_fp_stdata_bits_data; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_predicated; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_valid; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_switch; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_switch_off; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_unicore; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_shift; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_lrs3_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_rflag; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_wflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_prflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_pwflag; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_pflag_busy; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_stale_pflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_op1_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_op2_sel; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_split_num; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_self_index; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_rob_inst_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_address_num; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_uopc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_inst; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_debug_inst; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_rvc; // @[tile.scala 159:20]
  wire [39:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_debug_pc; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_iq_type; // @[tile.scala 159:20]
  wire [9:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_fu_code; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_br_type; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_op1_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_op2_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_imm_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_op_fcn; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_fcn_dw; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_csr_cmd; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_is_load; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_is_sta; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_is_std; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_op3_sel; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_iw_state; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_iw_p1_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_iw_p2_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_br; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_jalr; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_jal; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_sfb; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_br_mask; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_br_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_edge_inst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_pc_lob; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_taken; // @[tile.scala 159:20]
  wire [19:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_imm_packed; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_csr_addr; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_rob_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_ldq_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_stq_idx; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_rxq_idx; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_pdst; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_prs1; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_prs2; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_prs3; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_ppred; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_prs1_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_prs2_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_prs3_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_ppred_busy; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_stale_pdst; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_exception; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_exc_cause; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_bypassable; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_mem_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_mem_size; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_mem_signed; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_fence; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_fencei; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_amo; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_uses_ldq; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_uses_stq; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_sys_pc2epc; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_unique; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_flush_on_commit; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_ldst_is_rs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_ldst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_lrs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_lrs2; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_lrs3; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_ldst_val; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_dst_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_lrs1_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_lrs2_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_frs3_en; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_fp_val; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_fp_single; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_xcpt_pf_if; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_xcpt_ae_if; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_xcpt_ma_if; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_bp_debug_if; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflags_bits_uop_bp_xcpt_if; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_debug_fsrc; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflags_bits_uop_debug_tsrc; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_fp_stdata_bits_fflags_bits_flags; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_flagdata; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_valid; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_switch; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_switch_off; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_unicore; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_shift; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs3_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_rflag; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_wflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_prflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_pwflag; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_pflag_busy; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_stale_pflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_op1_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_op2_sel; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_split_num; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_self_index; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_rob_inst_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_address_num; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_uopc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_inst; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_debug_inst; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_rvc; // @[tile.scala 159:20]
  wire [39:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_debug_pc; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_iq_type; // @[tile.scala 159:20]
  wire [9:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_fu_code; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_br_type; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_op1_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_op2_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_imm_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_op_fcn; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_fcn_dw; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_csr_cmd; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_load; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_sta; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_std; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_op3_sel; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_iw_state; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_iw_p1_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_iw_p2_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_br; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_jalr; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_jal; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_sfb; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_br_mask; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_br_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_edge_inst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_pc_lob; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_taken; // @[tile.scala 159:20]
  wire [19:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_imm_packed; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_csr_addr; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_rob_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ldq_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_stq_idx; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_rxq_idx; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_pdst; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs1; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs2; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs3; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ppred; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs1_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs2_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs3_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ppred_busy; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_stale_pdst; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_exception; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_exc_cause; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_bypassable; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_mem_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_mem_size; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_mem_signed; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_fence; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_fencei; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_amo; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_uses_ldq; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_uses_stq; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_sys_pc2epc; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_unique; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_flush_on_commit; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ldst_is_rs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ldst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs2; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs3; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ldst_val; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_dst_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs1_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs2_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_frs3_en; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_fp_val; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_fp_single; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_xcpt_pf_if; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_xcpt_ae_if; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_xcpt_ma_if; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_bp_debug_if; // @[tile.scala 159:20]
  wire  core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_bp_xcpt_if; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_debug_fsrc; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_debug_tsrc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_fp_stdata_bits_fflagdata_bits_fflag; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_valids_0; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_valids_1; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_arch_valids_0; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_arch_valids_1; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_switch; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_switch_off; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_is_unicore; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_commit_uops_0_shift; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_0_lrs3_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_rflag; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_wflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_commit_uops_0_prflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_commit_uops_0_pwflag; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_pflag_busy; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_commit_uops_0_stale_pflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_commit_uops_0_op1_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_commit_uops_0_op2_sel; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_commit_uops_0_split_num; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_commit_uops_0_self_index; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_commit_uops_0_rob_inst_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_commit_uops_0_address_num; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_commit_uops_0_uopc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_commit_uops_0_inst; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_commit_uops_0_debug_inst; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_is_rvc; // @[tile.scala 159:20]
  wire [39:0] core_io_lsu_commit_uops_0_debug_pc; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_commit_uops_0_iq_type; // @[tile.scala 159:20]
  wire [9:0] core_io_lsu_commit_uops_0_fu_code; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_commit_uops_0_ctrl_br_type; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_0_ctrl_op1_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_commit_uops_0_ctrl_op2_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_commit_uops_0_ctrl_imm_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_commit_uops_0_ctrl_op_fcn; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_ctrl_fcn_dw; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_commit_uops_0_ctrl_csr_cmd; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_ctrl_is_load; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_ctrl_is_sta; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_ctrl_is_std; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_0_ctrl_op3_sel; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_0_iw_state; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_iw_p1_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_iw_p2_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_is_br; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_is_jalr; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_is_jal; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_is_sfb; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_commit_uops_0_br_mask; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_commit_uops_0_br_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_commit_uops_0_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_edge_inst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_commit_uops_0_pc_lob; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_taken; // @[tile.scala 159:20]
  wire [19:0] core_io_lsu_commit_uops_0_imm_packed; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_commit_uops_0_csr_addr; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_commit_uops_0_rob_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_commit_uops_0_ldq_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_commit_uops_0_stq_idx; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_0_rxq_idx; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_commit_uops_0_pdst; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_commit_uops_0_prs1; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_commit_uops_0_prs2; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_commit_uops_0_prs3; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_commit_uops_0_ppred; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_prs1_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_prs2_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_prs3_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_ppred_busy; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_commit_uops_0_stale_pdst; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_exception; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_commit_uops_0_exc_cause; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_bypassable; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_commit_uops_0_mem_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_0_mem_size; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_mem_signed; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_is_fence; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_is_fencei; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_is_amo; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_uses_ldq; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_uses_stq; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_is_sys_pc2epc; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_is_unique; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_flush_on_commit; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_ldst_is_rs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_commit_uops_0_ldst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_commit_uops_0_lrs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_commit_uops_0_lrs2; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_commit_uops_0_lrs3; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_ldst_val; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_0_dst_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_0_lrs1_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_0_lrs2_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_frs3_en; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_fp_val; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_fp_single; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_xcpt_pf_if; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_xcpt_ae_if; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_xcpt_ma_if; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_bp_debug_if; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_0_bp_xcpt_if; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_0_debug_fsrc; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_0_debug_tsrc; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_switch; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_switch_off; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_is_unicore; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_commit_uops_1_shift; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_1_lrs3_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_rflag; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_wflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_commit_uops_1_prflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_commit_uops_1_pwflag; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_pflag_busy; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_commit_uops_1_stale_pflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_commit_uops_1_op1_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_commit_uops_1_op2_sel; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_commit_uops_1_split_num; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_commit_uops_1_self_index; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_commit_uops_1_rob_inst_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_commit_uops_1_address_num; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_commit_uops_1_uopc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_commit_uops_1_inst; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_commit_uops_1_debug_inst; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_is_rvc; // @[tile.scala 159:20]
  wire [39:0] core_io_lsu_commit_uops_1_debug_pc; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_commit_uops_1_iq_type; // @[tile.scala 159:20]
  wire [9:0] core_io_lsu_commit_uops_1_fu_code; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_commit_uops_1_ctrl_br_type; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_1_ctrl_op1_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_commit_uops_1_ctrl_op2_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_commit_uops_1_ctrl_imm_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_commit_uops_1_ctrl_op_fcn; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_ctrl_fcn_dw; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_commit_uops_1_ctrl_csr_cmd; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_ctrl_is_load; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_ctrl_is_sta; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_ctrl_is_std; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_1_ctrl_op3_sel; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_1_iw_state; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_iw_p1_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_iw_p2_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_is_br; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_is_jalr; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_is_jal; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_is_sfb; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_commit_uops_1_br_mask; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_commit_uops_1_br_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_commit_uops_1_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_edge_inst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_commit_uops_1_pc_lob; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_taken; // @[tile.scala 159:20]
  wire [19:0] core_io_lsu_commit_uops_1_imm_packed; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_commit_uops_1_csr_addr; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_commit_uops_1_rob_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_commit_uops_1_ldq_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_commit_uops_1_stq_idx; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_1_rxq_idx; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_commit_uops_1_pdst; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_commit_uops_1_prs1; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_commit_uops_1_prs2; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_commit_uops_1_prs3; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_commit_uops_1_ppred; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_prs1_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_prs2_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_prs3_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_ppred_busy; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_commit_uops_1_stale_pdst; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_exception; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_commit_uops_1_exc_cause; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_bypassable; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_commit_uops_1_mem_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_1_mem_size; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_mem_signed; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_is_fence; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_is_fencei; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_is_amo; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_uses_ldq; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_uses_stq; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_is_sys_pc2epc; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_is_unique; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_flush_on_commit; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_ldst_is_rs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_commit_uops_1_ldst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_commit_uops_1_lrs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_commit_uops_1_lrs2; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_commit_uops_1_lrs3; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_ldst_val; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_1_dst_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_1_lrs1_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_1_lrs2_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_frs3_en; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_fp_val; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_fp_single; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_xcpt_pf_if; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_xcpt_ae_if; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_xcpt_ma_if; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_bp_debug_if; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_uops_1_bp_xcpt_if; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_1_debug_fsrc; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_commit_uops_1_debug_tsrc; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_fflags_valid; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_commit_fflags_bits; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_fflag_exception_valid; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_commit_fflag_exception_bits; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_commit_debug_insts_0; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_commit_debug_insts_1; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_rbk_valids_0; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_rbk_valids_1; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_rollback; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_commit_debug_wdata_0; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_commit_debug_wdata_1; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_commit_debug_wflagdata_0; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_commit_debug_wflagdata_1; // @[tile.scala 159:20]
  wire  core_io_lsu_commit_load_at_rob_head; // @[tile.scala 159:20]
  wire  core_io_lsu_clr_bsy_0_valid; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_clr_bsy_0_bits; // @[tile.scala 159:20]
  wire  core_io_lsu_clr_bsy_1_valid; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_clr_bsy_1_bits; // @[tile.scala 159:20]
  wire  core_io_lsu_clr_unsafe_0_valid; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_clr_unsafe_0_bits; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_clr_bsy_first_idx_0; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_clr_bsy_first_idx_1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_clr_bsy_self_idx_0; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_clr_bsy_self_idx_1; // @[tile.scala 159:20]
  wire  core_io_lsu_fence_dmem; // @[tile.scala 159:20]
  wire  core_io_lsu_spec_ld_wakeup_0_valid; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_spec_ld_wakeup_0_bits; // @[tile.scala 159:20]
  wire  core_io_lsu_ld_miss; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_brupdate_b1_resolve_mask; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_brupdate_b1_mispredict_mask; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_switch; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_switch_off; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_is_unicore; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_brupdate_b2_uop_shift; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_brupdate_b2_uop_lrs3_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_rflag; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_wflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_brupdate_b2_uop_prflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_brupdate_b2_uop_pwflag; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_pflag_busy; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_brupdate_b2_uop_stale_pflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_brupdate_b2_uop_op1_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_brupdate_b2_uop_op2_sel; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_brupdate_b2_uop_split_num; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_brupdate_b2_uop_self_index; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_brupdate_b2_uop_rob_inst_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_brupdate_b2_uop_address_num; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_brupdate_b2_uop_uopc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_brupdate_b2_uop_inst; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_brupdate_b2_uop_debug_inst; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_is_rvc; // @[tile.scala 159:20]
  wire [39:0] core_io_lsu_brupdate_b2_uop_debug_pc; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_brupdate_b2_uop_iq_type; // @[tile.scala 159:20]
  wire [9:0] core_io_lsu_brupdate_b2_uop_fu_code; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_brupdate_b2_uop_ctrl_br_type; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_brupdate_b2_uop_ctrl_op1_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_brupdate_b2_uop_ctrl_op2_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_brupdate_b2_uop_ctrl_imm_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_brupdate_b2_uop_ctrl_op_fcn; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_ctrl_fcn_dw; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_brupdate_b2_uop_ctrl_csr_cmd; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_ctrl_is_load; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_ctrl_is_sta; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_ctrl_is_std; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_brupdate_b2_uop_ctrl_op3_sel; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_brupdate_b2_uop_iw_state; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_iw_p1_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_iw_p2_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_is_br; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_is_jalr; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_is_jal; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_is_sfb; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_brupdate_b2_uop_br_mask; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_brupdate_b2_uop_br_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_brupdate_b2_uop_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_edge_inst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_brupdate_b2_uop_pc_lob; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_taken; // @[tile.scala 159:20]
  wire [19:0] core_io_lsu_brupdate_b2_uop_imm_packed; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_brupdate_b2_uop_csr_addr; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_brupdate_b2_uop_rob_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_brupdate_b2_uop_ldq_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_brupdate_b2_uop_stq_idx; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_brupdate_b2_uop_rxq_idx; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_brupdate_b2_uop_pdst; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_brupdate_b2_uop_prs1; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_brupdate_b2_uop_prs2; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_brupdate_b2_uop_prs3; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_brupdate_b2_uop_ppred; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_prs1_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_prs2_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_prs3_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_ppred_busy; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_brupdate_b2_uop_stale_pdst; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_exception; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_brupdate_b2_uop_exc_cause; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_bypassable; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_brupdate_b2_uop_mem_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_brupdate_b2_uop_mem_size; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_mem_signed; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_is_fence; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_is_fencei; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_is_amo; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_uses_ldq; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_uses_stq; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_is_sys_pc2epc; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_is_unique; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_flush_on_commit; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_ldst_is_rs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_brupdate_b2_uop_ldst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_brupdate_b2_uop_lrs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_brupdate_b2_uop_lrs2; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_brupdate_b2_uop_lrs3; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_ldst_val; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_brupdate_b2_uop_dst_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_brupdate_b2_uop_lrs1_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_brupdate_b2_uop_lrs2_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_frs3_en; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_fp_val; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_fp_single; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_xcpt_pf_if; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_xcpt_ae_if; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_xcpt_ma_if; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_bp_debug_if; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_uop_bp_xcpt_if; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_brupdate_b2_uop_debug_fsrc; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_brupdate_b2_uop_debug_tsrc; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_valid; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_mispredict; // @[tile.scala 159:20]
  wire  core_io_lsu_brupdate_b2_taken; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_brupdate_b2_cfi_type; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_brupdate_b2_pc_sel; // @[tile.scala 159:20]
  wire [39:0] core_io_lsu_brupdate_b2_jalr_target; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_brupdate_b2_target_offset; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_rob_pnr_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_rob_head_idx; // @[tile.scala 159:20]
  wire  core_io_lsu_exception; // @[tile.scala 159:20]
  wire  core_io_lsu_fencei_rdy; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_valid; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_switch; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_switch_off; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_is_unicore; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_lxcpt_bits_uop_shift; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_lxcpt_bits_uop_lrs3_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_rflag; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_wflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_lxcpt_bits_uop_prflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_lxcpt_bits_uop_pwflag; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_pflag_busy; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_lxcpt_bits_uop_stale_pflag; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_lxcpt_bits_uop_op1_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_lxcpt_bits_uop_op2_sel; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_lxcpt_bits_uop_split_num; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_lxcpt_bits_uop_self_index; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_lxcpt_bits_uop_rob_inst_idx; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_lxcpt_bits_uop_address_num; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_lxcpt_bits_uop_uopc; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_lxcpt_bits_uop_inst; // @[tile.scala 159:20]
  wire [31:0] core_io_lsu_lxcpt_bits_uop_debug_inst; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_is_rvc; // @[tile.scala 159:20]
  wire [39:0] core_io_lsu_lxcpt_bits_uop_debug_pc; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_lxcpt_bits_uop_iq_type; // @[tile.scala 159:20]
  wire [9:0] core_io_lsu_lxcpt_bits_uop_fu_code; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_lxcpt_bits_uop_ctrl_br_type; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_lxcpt_bits_uop_ctrl_op1_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_lxcpt_bits_uop_ctrl_op2_sel; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_lxcpt_bits_uop_ctrl_imm_sel; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_lxcpt_bits_uop_ctrl_op_fcn; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_ctrl_fcn_dw; // @[tile.scala 159:20]
  wire [2:0] core_io_lsu_lxcpt_bits_uop_ctrl_csr_cmd; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_ctrl_is_load; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_ctrl_is_sta; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_ctrl_is_std; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_lxcpt_bits_uop_ctrl_op3_sel; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_lxcpt_bits_uop_iw_state; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_iw_p1_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_iw_p2_poisoned; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_is_br; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_is_jalr; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_is_jal; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_is_sfb; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_lxcpt_bits_uop_br_mask; // @[tile.scala 159:20]
  wire [3:0] core_io_lsu_lxcpt_bits_uop_br_tag; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_lxcpt_bits_uop_ftq_idx; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_edge_inst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_lxcpt_bits_uop_pc_lob; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_taken; // @[tile.scala 159:20]
  wire [19:0] core_io_lsu_lxcpt_bits_uop_imm_packed; // @[tile.scala 159:20]
  wire [11:0] core_io_lsu_lxcpt_bits_uop_csr_addr; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_lxcpt_bits_uop_rob_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_lxcpt_bits_uop_ldq_idx; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_lxcpt_bits_uop_stq_idx; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_lxcpt_bits_uop_rxq_idx; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_lxcpt_bits_uop_pdst; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_lxcpt_bits_uop_prs1; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_lxcpt_bits_uop_prs2; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_lxcpt_bits_uop_prs3; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_lxcpt_bits_uop_ppred; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_prs1_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_prs2_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_prs3_busy; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_ppred_busy; // @[tile.scala 159:20]
  wire [6:0] core_io_lsu_lxcpt_bits_uop_stale_pdst; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_exception; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_lxcpt_bits_uop_exc_cause; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_bypassable; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_lxcpt_bits_uop_mem_cmd; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_lxcpt_bits_uop_mem_size; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_mem_signed; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_is_fence; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_is_fencei; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_is_amo; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_uses_ldq; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_uses_stq; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_is_sys_pc2epc; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_is_unique; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_flush_on_commit; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_ldst_is_rs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_lxcpt_bits_uop_ldst; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_lxcpt_bits_uop_lrs1; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_lxcpt_bits_uop_lrs2; // @[tile.scala 159:20]
  wire [5:0] core_io_lsu_lxcpt_bits_uop_lrs3; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_ldst_val; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_lxcpt_bits_uop_dst_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_lxcpt_bits_uop_lrs1_rtype; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_lxcpt_bits_uop_lrs2_rtype; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_frs3_en; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_fp_val; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_fp_single; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_xcpt_pf_if; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_xcpt_ae_if; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_xcpt_ma_if; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_bp_debug_if; // @[tile.scala 159:20]
  wire  core_io_lsu_lxcpt_bits_uop_bp_xcpt_if; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_lxcpt_bits_uop_debug_fsrc; // @[tile.scala 159:20]
  wire [1:0] core_io_lsu_lxcpt_bits_uop_debug_tsrc; // @[tile.scala 159:20]
  wire [4:0] core_io_lsu_lxcpt_bits_cause; // @[tile.scala 159:20]
  wire [39:0] core_io_lsu_lxcpt_bits_badvaddr; // @[tile.scala 159:20]
  wire [63:0] core_io_lsu_tsc_reg; // @[tile.scala 159:20]
  wire  core_io_lsu_perf_acquire; // @[tile.scala 159:20]
  wire  core_io_lsu_perf_release; // @[tile.scala 159:20]
  wire  core_io_lsu_perf_tlbMiss; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_req_ready; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_req_valid; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_req_bits_valid; // @[tile.scala 159:20]
  wire [26:0] core_io_ptw_tlb_req_bits_bits_addr; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_resp_valid; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_resp_bits_ae; // @[tile.scala 159:20]
  wire [53:0] core_io_ptw_tlb_resp_bits_pte_ppn; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_resp_bits_pte_reserved_for_software; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_resp_bits_pte_d; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_resp_bits_pte_a; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_resp_bits_pte_g; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_resp_bits_pte_u; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_resp_bits_pte_x; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_resp_bits_pte_w; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_resp_bits_pte_r; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_resp_bits_pte_v; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_resp_bits_level; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_resp_bits_fragmented_superpage; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_resp_bits_homogeneous; // @[tile.scala 159:20]
  wire [3:0] core_io_ptw_tlb_ptbr_mode; // @[tile.scala 159:20]
  wire [15:0] core_io_ptw_tlb_ptbr_asid; // @[tile.scala 159:20]
  wire [43:0] core_io_ptw_tlb_ptbr_ppn; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_status_debug; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_status_cease; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_status_wfi; // @[tile.scala 159:20]
  wire [31:0] core_io_ptw_tlb_status_isa; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_status_dprv; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_status_prv; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_status_sd; // @[tile.scala 159:20]
  wire [26:0] core_io_ptw_tlb_status_zero2; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_status_sxl; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_status_uxl; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_status_sd_rv32; // @[tile.scala 159:20]
  wire [7:0] core_io_ptw_tlb_status_zero1; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_status_tsr; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_status_tw; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_status_tvm; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_status_mxr; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_status_sum; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_status_mprv; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_status_xs; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_status_fs; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_status_mpp; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_status_vs; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_status_spp; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_status_mpie; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_status_hpie; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_status_spie; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_status_upie; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_status_mie; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_status_hie; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_status_sie; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_status_uie; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_0_cfg_l; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_pmp_0_cfg_res; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_pmp_0_cfg_a; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_0_cfg_x; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_0_cfg_w; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_0_cfg_r; // @[tile.scala 159:20]
  wire [29:0] core_io_ptw_tlb_pmp_0_addr; // @[tile.scala 159:20]
  wire [31:0] core_io_ptw_tlb_pmp_0_mask; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_1_cfg_l; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_pmp_1_cfg_res; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_pmp_1_cfg_a; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_1_cfg_x; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_1_cfg_w; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_1_cfg_r; // @[tile.scala 159:20]
  wire [29:0] core_io_ptw_tlb_pmp_1_addr; // @[tile.scala 159:20]
  wire [31:0] core_io_ptw_tlb_pmp_1_mask; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_2_cfg_l; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_pmp_2_cfg_res; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_pmp_2_cfg_a; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_2_cfg_x; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_2_cfg_w; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_2_cfg_r; // @[tile.scala 159:20]
  wire [29:0] core_io_ptw_tlb_pmp_2_addr; // @[tile.scala 159:20]
  wire [31:0] core_io_ptw_tlb_pmp_2_mask; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_3_cfg_l; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_pmp_3_cfg_res; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_pmp_3_cfg_a; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_3_cfg_x; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_3_cfg_w; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_3_cfg_r; // @[tile.scala 159:20]
  wire [29:0] core_io_ptw_tlb_pmp_3_addr; // @[tile.scala 159:20]
  wire [31:0] core_io_ptw_tlb_pmp_3_mask; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_4_cfg_l; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_pmp_4_cfg_res; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_pmp_4_cfg_a; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_4_cfg_x; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_4_cfg_w; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_4_cfg_r; // @[tile.scala 159:20]
  wire [29:0] core_io_ptw_tlb_pmp_4_addr; // @[tile.scala 159:20]
  wire [31:0] core_io_ptw_tlb_pmp_4_mask; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_5_cfg_l; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_pmp_5_cfg_res; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_pmp_5_cfg_a; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_5_cfg_x; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_5_cfg_w; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_5_cfg_r; // @[tile.scala 159:20]
  wire [29:0] core_io_ptw_tlb_pmp_5_addr; // @[tile.scala 159:20]
  wire [31:0] core_io_ptw_tlb_pmp_5_mask; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_6_cfg_l; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_pmp_6_cfg_res; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_pmp_6_cfg_a; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_6_cfg_x; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_6_cfg_w; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_6_cfg_r; // @[tile.scala 159:20]
  wire [29:0] core_io_ptw_tlb_pmp_6_addr; // @[tile.scala 159:20]
  wire [31:0] core_io_ptw_tlb_pmp_6_mask; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_7_cfg_l; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_pmp_7_cfg_res; // @[tile.scala 159:20]
  wire [1:0] core_io_ptw_tlb_pmp_7_cfg_a; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_7_cfg_x; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_7_cfg_w; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_pmp_7_cfg_r; // @[tile.scala 159:20]
  wire [29:0] core_io_ptw_tlb_pmp_7_addr; // @[tile.scala 159:20]
  wire [31:0] core_io_ptw_tlb_pmp_7_mask; // @[tile.scala 159:20]
  wire  core_io_ptw_tlb_customCSRs_csrs_0_wen; // @[tile.scala 159:20]
  wire [63:0] core_io_ptw_tlb_customCSRs_csrs_0_wdata; // @[tile.scala 159:20]
  wire [63:0] core_io_ptw_tlb_customCSRs_csrs_0_value; // @[tile.scala 159:20]
  wire  core_io_trace_0_valid; // @[tile.scala 159:20]
  wire [39:0] core_io_trace_0_iaddr; // @[tile.scala 159:20]
  wire [31:0] core_io_trace_0_insn; // @[tile.scala 159:20]
  wire [2:0] core_io_trace_0_priv; // @[tile.scala 159:20]
  wire  core_io_trace_0_exception; // @[tile.scala 159:20]
  wire  core_io_trace_0_interrupt; // @[tile.scala 159:20]
  wire [63:0] core_io_trace_0_cause; // @[tile.scala 159:20]
  wire [39:0] core_io_trace_0_tval; // @[tile.scala 159:20]
  wire [63:0] core_io_trace_0_wdata; // @[tile.scala 159:20]
  wire  core_io_trace_1_valid; // @[tile.scala 159:20]
  wire [39:0] core_io_trace_1_iaddr; // @[tile.scala 159:20]
  wire [31:0] core_io_trace_1_insn; // @[tile.scala 159:20]
  wire [2:0] core_io_trace_1_priv; // @[tile.scala 159:20]
  wire  core_io_trace_1_exception; // @[tile.scala 159:20]
  wire  core_io_trace_1_interrupt; // @[tile.scala 159:20]
  wire [63:0] core_io_trace_1_cause; // @[tile.scala 159:20]
  wire [39:0] core_io_trace_1_tval; // @[tile.scala 159:20]
  wire [63:0] core_io_trace_1_wdata; // @[tile.scala 159:20]
  wire [2:0] core_io_fcsr_rm; // @[tile.scala 159:20]
  wire  lsu_clock; // @[tile.scala 160:20]
  wire  lsu_reset; // @[tile.scala 160:20]
  wire  lsu_io_ptw_req_ready; // @[tile.scala 160:20]
  wire  lsu_io_ptw_req_valid; // @[tile.scala 160:20]
  wire  lsu_io_ptw_req_bits_valid; // @[tile.scala 160:20]
  wire [26:0] lsu_io_ptw_req_bits_bits_addr; // @[tile.scala 160:20]
  wire  lsu_io_ptw_resp_valid; // @[tile.scala 160:20]
  wire  lsu_io_ptw_resp_bits_ae; // @[tile.scala 160:20]
  wire [53:0] lsu_io_ptw_resp_bits_pte_ppn; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_resp_bits_pte_reserved_for_software; // @[tile.scala 160:20]
  wire  lsu_io_ptw_resp_bits_pte_d; // @[tile.scala 160:20]
  wire  lsu_io_ptw_resp_bits_pte_a; // @[tile.scala 160:20]
  wire  lsu_io_ptw_resp_bits_pte_g; // @[tile.scala 160:20]
  wire  lsu_io_ptw_resp_bits_pte_u; // @[tile.scala 160:20]
  wire  lsu_io_ptw_resp_bits_pte_x; // @[tile.scala 160:20]
  wire  lsu_io_ptw_resp_bits_pte_w; // @[tile.scala 160:20]
  wire  lsu_io_ptw_resp_bits_pte_r; // @[tile.scala 160:20]
  wire  lsu_io_ptw_resp_bits_pte_v; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_resp_bits_level; // @[tile.scala 160:20]
  wire  lsu_io_ptw_resp_bits_fragmented_superpage; // @[tile.scala 160:20]
  wire  lsu_io_ptw_resp_bits_homogeneous; // @[tile.scala 160:20]
  wire [3:0] lsu_io_ptw_ptbr_mode; // @[tile.scala 160:20]
  wire [15:0] lsu_io_ptw_ptbr_asid; // @[tile.scala 160:20]
  wire [43:0] lsu_io_ptw_ptbr_ppn; // @[tile.scala 160:20]
  wire  lsu_io_ptw_status_debug; // @[tile.scala 160:20]
  wire  lsu_io_ptw_status_cease; // @[tile.scala 160:20]
  wire  lsu_io_ptw_status_wfi; // @[tile.scala 160:20]
  wire [31:0] lsu_io_ptw_status_isa; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_status_dprv; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_status_prv; // @[tile.scala 160:20]
  wire  lsu_io_ptw_status_sd; // @[tile.scala 160:20]
  wire [26:0] lsu_io_ptw_status_zero2; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_status_sxl; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_status_uxl; // @[tile.scala 160:20]
  wire  lsu_io_ptw_status_sd_rv32; // @[tile.scala 160:20]
  wire [7:0] lsu_io_ptw_status_zero1; // @[tile.scala 160:20]
  wire  lsu_io_ptw_status_tsr; // @[tile.scala 160:20]
  wire  lsu_io_ptw_status_tw; // @[tile.scala 160:20]
  wire  lsu_io_ptw_status_tvm; // @[tile.scala 160:20]
  wire  lsu_io_ptw_status_mxr; // @[tile.scala 160:20]
  wire  lsu_io_ptw_status_sum; // @[tile.scala 160:20]
  wire  lsu_io_ptw_status_mprv; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_status_xs; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_status_fs; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_status_mpp; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_status_vs; // @[tile.scala 160:20]
  wire  lsu_io_ptw_status_spp; // @[tile.scala 160:20]
  wire  lsu_io_ptw_status_mpie; // @[tile.scala 160:20]
  wire  lsu_io_ptw_status_hpie; // @[tile.scala 160:20]
  wire  lsu_io_ptw_status_spie; // @[tile.scala 160:20]
  wire  lsu_io_ptw_status_upie; // @[tile.scala 160:20]
  wire  lsu_io_ptw_status_mie; // @[tile.scala 160:20]
  wire  lsu_io_ptw_status_hie; // @[tile.scala 160:20]
  wire  lsu_io_ptw_status_sie; // @[tile.scala 160:20]
  wire  lsu_io_ptw_status_uie; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_0_cfg_l; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_pmp_0_cfg_res; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_pmp_0_cfg_a; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_0_cfg_x; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_0_cfg_w; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_0_cfg_r; // @[tile.scala 160:20]
  wire [29:0] lsu_io_ptw_pmp_0_addr; // @[tile.scala 160:20]
  wire [31:0] lsu_io_ptw_pmp_0_mask; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_1_cfg_l; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_pmp_1_cfg_res; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_pmp_1_cfg_a; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_1_cfg_x; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_1_cfg_w; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_1_cfg_r; // @[tile.scala 160:20]
  wire [29:0] lsu_io_ptw_pmp_1_addr; // @[tile.scala 160:20]
  wire [31:0] lsu_io_ptw_pmp_1_mask; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_2_cfg_l; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_pmp_2_cfg_res; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_pmp_2_cfg_a; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_2_cfg_x; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_2_cfg_w; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_2_cfg_r; // @[tile.scala 160:20]
  wire [29:0] lsu_io_ptw_pmp_2_addr; // @[tile.scala 160:20]
  wire [31:0] lsu_io_ptw_pmp_2_mask; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_3_cfg_l; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_pmp_3_cfg_res; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_pmp_3_cfg_a; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_3_cfg_x; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_3_cfg_w; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_3_cfg_r; // @[tile.scala 160:20]
  wire [29:0] lsu_io_ptw_pmp_3_addr; // @[tile.scala 160:20]
  wire [31:0] lsu_io_ptw_pmp_3_mask; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_4_cfg_l; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_pmp_4_cfg_res; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_pmp_4_cfg_a; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_4_cfg_x; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_4_cfg_w; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_4_cfg_r; // @[tile.scala 160:20]
  wire [29:0] lsu_io_ptw_pmp_4_addr; // @[tile.scala 160:20]
  wire [31:0] lsu_io_ptw_pmp_4_mask; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_5_cfg_l; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_pmp_5_cfg_res; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_pmp_5_cfg_a; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_5_cfg_x; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_5_cfg_w; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_5_cfg_r; // @[tile.scala 160:20]
  wire [29:0] lsu_io_ptw_pmp_5_addr; // @[tile.scala 160:20]
  wire [31:0] lsu_io_ptw_pmp_5_mask; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_6_cfg_l; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_pmp_6_cfg_res; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_pmp_6_cfg_a; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_6_cfg_x; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_6_cfg_w; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_6_cfg_r; // @[tile.scala 160:20]
  wire [29:0] lsu_io_ptw_pmp_6_addr; // @[tile.scala 160:20]
  wire [31:0] lsu_io_ptw_pmp_6_mask; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_7_cfg_l; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_pmp_7_cfg_res; // @[tile.scala 160:20]
  wire [1:0] lsu_io_ptw_pmp_7_cfg_a; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_7_cfg_x; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_7_cfg_w; // @[tile.scala 160:20]
  wire  lsu_io_ptw_pmp_7_cfg_r; // @[tile.scala 160:20]
  wire [29:0] lsu_io_ptw_pmp_7_addr; // @[tile.scala 160:20]
  wire [31:0] lsu_io_ptw_pmp_7_mask; // @[tile.scala 160:20]
  wire  lsu_io_ptw_customCSRs_csrs_0_wen; // @[tile.scala 160:20]
  wire [63:0] lsu_io_ptw_customCSRs_csrs_0_wdata; // @[tile.scala 160:20]
  wire [63:0] lsu_io_ptw_customCSRs_csrs_0_value; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_valid; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_switch; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_req_bits_uop_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_uop_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_rflag; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_uop_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_uop_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_uop_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_uop_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_uop_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_uop_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_uop_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_uop_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_uop_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_req_bits_uop_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_exe_0_req_bits_uop_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_exe_0_req_bits_uop_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_core_exe_0_req_bits_uop_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_req_bits_uop_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_core_exe_0_req_bits_uop_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_uop_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_uop_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_req_bits_uop_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_req_bits_uop_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_uop_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_req_bits_uop_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_uop_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_uop_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_is_br; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_exe_0_req_bits_uop_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_uop_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_req_bits_uop_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_uop_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_core_exe_0_req_bits_uop_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_exe_0_req_bits_uop_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_uop_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_req_bits_uop_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_req_bits_uop_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_uop_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_req_bits_uop_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_req_bits_uop_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_req_bits_uop_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_req_bits_uop_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_req_bits_uop_ppred; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_req_bits_uop_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_exe_0_req_bits_uop_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_req_bits_uop_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_uop_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_uop_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_uop_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_uop_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_uop_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_uop_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_uop_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_uop_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_uop_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_uop_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_uop_debug_tsrc; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_predicated; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_exe_0_req_bits_data; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_valid; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_switch; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_rflag; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_br; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_ppred; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflags_bits_uop_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflags_bits_uop_debug_tsrc; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_req_bits_fflags_bits_flags; // @[tile.scala 160:20]
  wire [39:0] lsu_io_core_exe_0_req_bits_addr; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_mxcpt_valid; // @[tile.scala 160:20]
  wire [16:0] lsu_io_core_exe_0_req_bits_mxcpt_bits; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_sfence_valid; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_sfence_bits_rs1; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_sfence_bits_rs2; // @[tile.scala 160:20]
  wire [38:0] lsu_io_core_exe_0_req_bits_sfence_bits_addr; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_sfence_bits_asid; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_flagdata; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_valid; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_switch; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_rflag; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_br; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ppred; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_debug_tsrc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_exe_0_req_bits_fflagdata_bits_fflag; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_ready; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_valid; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_switch; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_iresp_bits_uop_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_uop_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_rflag; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_uop_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_uop_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_uop_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_uop_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_uop_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_uop_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_uop_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_uop_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_uop_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_iresp_bits_uop_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_exe_0_iresp_bits_uop_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_exe_0_iresp_bits_uop_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_core_exe_0_iresp_bits_uop_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_iresp_bits_uop_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_core_exe_0_iresp_bits_uop_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_uop_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_uop_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_iresp_bits_uop_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_iresp_bits_uop_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_uop_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_iresp_bits_uop_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_uop_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_uop_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_is_br; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_exe_0_iresp_bits_uop_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_uop_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_iresp_bits_uop_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_uop_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_core_exe_0_iresp_bits_uop_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_exe_0_iresp_bits_uop_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_uop_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_iresp_bits_uop_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_iresp_bits_uop_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_uop_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_iresp_bits_uop_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_iresp_bits_uop_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_iresp_bits_uop_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_iresp_bits_uop_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_iresp_bits_uop_ppred; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_iresp_bits_uop_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_exe_0_iresp_bits_uop_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_iresp_bits_uop_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_uop_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_uop_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_uop_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_uop_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_uop_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_uop_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_uop_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_uop_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_uop_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_uop_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_uop_debug_tsrc; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_exe_0_iresp_bits_data; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_predicated; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_valid; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_switch; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_rflag; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_br; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ppred; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_debug_tsrc; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_iresp_bits_fflags_bits_flags; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_flagdata; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_valid; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_switch; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_rflag; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_br; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ppred; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_debug_tsrc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_exe_0_iresp_bits_fflagdata_bits_fflag; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_ready; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_valid; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_switch; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_fresp_bits_uop_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_uop_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_rflag; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_uop_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_uop_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_uop_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_uop_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_uop_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_uop_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_uop_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_uop_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_uop_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_fresp_bits_uop_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_exe_0_fresp_bits_uop_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_exe_0_fresp_bits_uop_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_core_exe_0_fresp_bits_uop_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_fresp_bits_uop_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_core_exe_0_fresp_bits_uop_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_uop_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_uop_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_fresp_bits_uop_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_fresp_bits_uop_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_uop_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_fresp_bits_uop_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_uop_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_uop_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_is_br; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_exe_0_fresp_bits_uop_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_uop_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_fresp_bits_uop_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_uop_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_core_exe_0_fresp_bits_uop_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_exe_0_fresp_bits_uop_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_uop_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_fresp_bits_uop_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_fresp_bits_uop_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_uop_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_fresp_bits_uop_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_fresp_bits_uop_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_fresp_bits_uop_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_fresp_bits_uop_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_fresp_bits_uop_ppred; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_fresp_bits_uop_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_exe_0_fresp_bits_uop_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_fresp_bits_uop_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_uop_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_uop_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_uop_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_uop_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_uop_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_uop_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_uop_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_uop_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_uop_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_uop_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_uop_debug_tsrc; // @[tile.scala 160:20]
  wire [64:0] lsu_io_core_exe_0_fresp_bits_data; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_predicated; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_valid; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_switch; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_rflag; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_br; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ppred; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_debug_tsrc; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_fresp_bits_fflags_bits_flags; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_flagdata; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_valid; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_switch; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_rflag; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_br; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ppred; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_debug_tsrc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_exe_0_fresp_bits_fflagdata_bits_fflag; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_valid; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_switch; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_dis_uops_0_bits_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_0_bits_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_rflag; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_dis_uops_0_bits_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_dis_uops_0_bits_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_dis_uops_0_bits_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_dis_uops_0_bits_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_dis_uops_0_bits_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_dis_uops_0_bits_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_dis_uops_0_bits_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_dis_uops_0_bits_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_dis_uops_0_bits_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_dis_uops_0_bits_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_dis_uops_0_bits_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_dis_uops_0_bits_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_core_dis_uops_0_bits_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_dis_uops_0_bits_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_core_dis_uops_0_bits_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_dis_uops_0_bits_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_0_bits_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_dis_uops_0_bits_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_dis_uops_0_bits_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_dis_uops_0_bits_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_dis_uops_0_bits_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_0_bits_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_0_bits_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_is_br; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_dis_uops_0_bits_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_dis_uops_0_bits_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_dis_uops_0_bits_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_dis_uops_0_bits_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_core_dis_uops_0_bits_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_dis_uops_0_bits_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_dis_uops_0_bits_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_dis_uops_0_bits_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_dis_uops_0_bits_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_0_bits_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_dis_uops_0_bits_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_dis_uops_0_bits_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_dis_uops_0_bits_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_dis_uops_0_bits_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_dis_uops_0_bits_ppred; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_dis_uops_0_bits_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_dis_uops_0_bits_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_dis_uops_0_bits_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_0_bits_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_dis_uops_0_bits_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_dis_uops_0_bits_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_dis_uops_0_bits_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_dis_uops_0_bits_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_0_bits_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_0_bits_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_0_bits_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_0_bits_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_0_bits_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_0_bits_debug_tsrc; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_valid; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_switch; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_dis_uops_1_bits_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_1_bits_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_rflag; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_dis_uops_1_bits_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_dis_uops_1_bits_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_dis_uops_1_bits_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_dis_uops_1_bits_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_dis_uops_1_bits_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_dis_uops_1_bits_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_dis_uops_1_bits_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_dis_uops_1_bits_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_dis_uops_1_bits_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_dis_uops_1_bits_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_dis_uops_1_bits_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_dis_uops_1_bits_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_core_dis_uops_1_bits_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_dis_uops_1_bits_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_core_dis_uops_1_bits_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_dis_uops_1_bits_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_1_bits_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_dis_uops_1_bits_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_dis_uops_1_bits_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_dis_uops_1_bits_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_dis_uops_1_bits_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_1_bits_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_1_bits_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_is_br; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_dis_uops_1_bits_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_dis_uops_1_bits_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_dis_uops_1_bits_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_dis_uops_1_bits_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_core_dis_uops_1_bits_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_dis_uops_1_bits_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_dis_uops_1_bits_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_dis_uops_1_bits_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_dis_uops_1_bits_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_1_bits_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_dis_uops_1_bits_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_dis_uops_1_bits_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_dis_uops_1_bits_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_dis_uops_1_bits_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_dis_uops_1_bits_ppred; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_dis_uops_1_bits_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_dis_uops_1_bits_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_dis_uops_1_bits_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_1_bits_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_dis_uops_1_bits_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_dis_uops_1_bits_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_dis_uops_1_bits_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_dis_uops_1_bits_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_1_bits_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_1_bits_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_1_bits_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_core_dis_uops_1_bits_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_1_bits_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_dis_uops_1_bits_debug_tsrc; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_dis_ldq_idx_0; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_dis_ldq_idx_1; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_dis_stq_idx_0; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_dis_stq_idx_1; // @[tile.scala 160:20]
  wire  lsu_io_core_ldq_full_0; // @[tile.scala 160:20]
  wire  lsu_io_core_ldq_full_1; // @[tile.scala 160:20]
  wire  lsu_io_core_stq_full_0; // @[tile.scala 160:20]
  wire  lsu_io_core_stq_full_1; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_ready; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_valid; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_switch; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_fp_stdata_bits_uop_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_uop_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_rflag; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_uop_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_uop_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_uop_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_uop_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_uop_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_uop_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_uop_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_uop_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_uop_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_fp_stdata_bits_uop_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_fp_stdata_bits_uop_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_fp_stdata_bits_uop_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_core_fp_stdata_bits_uop_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_fp_stdata_bits_uop_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_core_fp_stdata_bits_uop_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_uop_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_uop_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_fp_stdata_bits_uop_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_fp_stdata_bits_uop_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_uop_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_fp_stdata_bits_uop_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_uop_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_uop_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_is_br; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_fp_stdata_bits_uop_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_uop_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_fp_stdata_bits_uop_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_uop_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_core_fp_stdata_bits_uop_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_fp_stdata_bits_uop_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_uop_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_fp_stdata_bits_uop_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_fp_stdata_bits_uop_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_uop_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_fp_stdata_bits_uop_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_fp_stdata_bits_uop_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_fp_stdata_bits_uop_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_fp_stdata_bits_uop_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_fp_stdata_bits_uop_ppred; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_fp_stdata_bits_uop_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_fp_stdata_bits_uop_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_fp_stdata_bits_uop_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_uop_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_uop_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_uop_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_uop_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_uop_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_uop_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_uop_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_uop_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_uop_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_uop_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_uop_debug_tsrc; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_fp_stdata_bits_data; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_predicated; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_valid; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_switch; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_rflag; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_br; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_ppred; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflags_bits_uop_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflags_bits_uop_debug_tsrc; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_fp_stdata_bits_fflags_bits_flags; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_flagdata; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_valid; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_switch; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_rflag; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_br; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ppred; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_debug_tsrc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_fp_stdata_bits_fflagdata_bits_fflag; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_valids_0; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_valids_1; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_arch_valids_0; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_arch_valids_1; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_switch; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_commit_uops_0_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_0_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_rflag; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_commit_uops_0_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_commit_uops_0_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_commit_uops_0_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_commit_uops_0_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_commit_uops_0_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_commit_uops_0_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_commit_uops_0_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_commit_uops_0_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_commit_uops_0_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_commit_uops_0_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_commit_uops_0_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_commit_uops_0_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_core_commit_uops_0_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_commit_uops_0_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_core_commit_uops_0_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_commit_uops_0_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_0_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_commit_uops_0_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_commit_uops_0_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_commit_uops_0_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_commit_uops_0_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_0_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_0_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_is_br; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_commit_uops_0_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_commit_uops_0_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_commit_uops_0_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_commit_uops_0_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_core_commit_uops_0_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_commit_uops_0_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_commit_uops_0_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_commit_uops_0_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_commit_uops_0_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_0_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_commit_uops_0_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_commit_uops_0_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_commit_uops_0_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_commit_uops_0_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_commit_uops_0_ppred; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_commit_uops_0_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_commit_uops_0_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_commit_uops_0_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_0_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_commit_uops_0_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_commit_uops_0_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_commit_uops_0_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_commit_uops_0_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_0_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_0_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_0_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_0_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_0_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_0_debug_tsrc; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_switch; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_commit_uops_1_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_1_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_rflag; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_commit_uops_1_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_commit_uops_1_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_commit_uops_1_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_commit_uops_1_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_commit_uops_1_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_commit_uops_1_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_commit_uops_1_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_commit_uops_1_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_commit_uops_1_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_commit_uops_1_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_commit_uops_1_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_commit_uops_1_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_core_commit_uops_1_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_commit_uops_1_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_core_commit_uops_1_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_commit_uops_1_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_1_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_commit_uops_1_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_commit_uops_1_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_commit_uops_1_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_commit_uops_1_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_1_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_1_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_is_br; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_commit_uops_1_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_commit_uops_1_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_commit_uops_1_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_commit_uops_1_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_core_commit_uops_1_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_commit_uops_1_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_commit_uops_1_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_commit_uops_1_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_commit_uops_1_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_1_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_commit_uops_1_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_commit_uops_1_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_commit_uops_1_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_commit_uops_1_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_commit_uops_1_ppred; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_commit_uops_1_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_commit_uops_1_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_commit_uops_1_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_1_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_commit_uops_1_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_commit_uops_1_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_commit_uops_1_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_commit_uops_1_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_1_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_1_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_1_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_uops_1_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_1_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_commit_uops_1_debug_tsrc; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_fflags_valid; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_commit_fflags_bits; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_fflag_exception_valid; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_commit_fflag_exception_bits; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_commit_debug_insts_0; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_commit_debug_insts_1; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_rbk_valids_0; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_rbk_valids_1; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_rollback; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_commit_debug_wdata_0; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_commit_debug_wdata_1; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_commit_debug_wflagdata_0; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_commit_debug_wflagdata_1; // @[tile.scala 160:20]
  wire  lsu_io_core_commit_load_at_rob_head; // @[tile.scala 160:20]
  wire  lsu_io_core_clr_bsy_0_valid; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_clr_bsy_0_bits; // @[tile.scala 160:20]
  wire  lsu_io_core_clr_bsy_1_valid; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_clr_bsy_1_bits; // @[tile.scala 160:20]
  wire  lsu_io_core_clr_unsafe_0_valid; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_clr_unsafe_0_bits; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_clr_bsy_first_idx_0; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_clr_bsy_first_idx_1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_clr_bsy_self_idx_0; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_clr_bsy_self_idx_1; // @[tile.scala 160:20]
  wire  lsu_io_core_fence_dmem; // @[tile.scala 160:20]
  wire  lsu_io_core_spec_ld_wakeup_0_valid; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_spec_ld_wakeup_0_bits; // @[tile.scala 160:20]
  wire  lsu_io_core_ld_miss; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_brupdate_b1_resolve_mask; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_brupdate_b1_mispredict_mask; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_switch; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_brupdate_b2_uop_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_brupdate_b2_uop_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_rflag; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_brupdate_b2_uop_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_brupdate_b2_uop_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_brupdate_b2_uop_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_brupdate_b2_uop_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_brupdate_b2_uop_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_brupdate_b2_uop_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_brupdate_b2_uop_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_brupdate_b2_uop_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_brupdate_b2_uop_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_brupdate_b2_uop_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_brupdate_b2_uop_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_brupdate_b2_uop_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_core_brupdate_b2_uop_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_brupdate_b2_uop_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_core_brupdate_b2_uop_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_brupdate_b2_uop_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_brupdate_b2_uop_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_brupdate_b2_uop_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_brupdate_b2_uop_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_brupdate_b2_uop_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_brupdate_b2_uop_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_brupdate_b2_uop_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_brupdate_b2_uop_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_is_br; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_brupdate_b2_uop_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_brupdate_b2_uop_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_brupdate_b2_uop_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_brupdate_b2_uop_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_core_brupdate_b2_uop_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_brupdate_b2_uop_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_brupdate_b2_uop_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_brupdate_b2_uop_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_brupdate_b2_uop_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_brupdate_b2_uop_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_brupdate_b2_uop_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_brupdate_b2_uop_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_brupdate_b2_uop_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_brupdate_b2_uop_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_brupdate_b2_uop_ppred; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_brupdate_b2_uop_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_brupdate_b2_uop_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_brupdate_b2_uop_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_brupdate_b2_uop_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_brupdate_b2_uop_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_brupdate_b2_uop_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_brupdate_b2_uop_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_brupdate_b2_uop_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_brupdate_b2_uop_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_brupdate_b2_uop_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_brupdate_b2_uop_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_uop_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_brupdate_b2_uop_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_brupdate_b2_uop_debug_tsrc; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_valid; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_mispredict; // @[tile.scala 160:20]
  wire  lsu_io_core_brupdate_b2_taken; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_brupdate_b2_cfi_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_brupdate_b2_pc_sel; // @[tile.scala 160:20]
  wire [39:0] lsu_io_core_brupdate_b2_jalr_target; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_brupdate_b2_target_offset; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_rob_pnr_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_rob_head_idx; // @[tile.scala 160:20]
  wire  lsu_io_core_exception; // @[tile.scala 160:20]
  wire  lsu_io_core_fencei_rdy; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_valid; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_switch; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_lxcpt_bits_uop_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_lxcpt_bits_uop_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_rflag; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_lxcpt_bits_uop_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_lxcpt_bits_uop_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_lxcpt_bits_uop_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_lxcpt_bits_uop_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_lxcpt_bits_uop_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_lxcpt_bits_uop_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_lxcpt_bits_uop_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_lxcpt_bits_uop_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_lxcpt_bits_uop_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_lxcpt_bits_uop_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_lxcpt_bits_uop_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_core_lxcpt_bits_uop_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_core_lxcpt_bits_uop_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_lxcpt_bits_uop_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_core_lxcpt_bits_uop_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_lxcpt_bits_uop_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_lxcpt_bits_uop_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_lxcpt_bits_uop_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_lxcpt_bits_uop_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_lxcpt_bits_uop_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_core_lxcpt_bits_uop_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_lxcpt_bits_uop_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_lxcpt_bits_uop_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_is_br; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_lxcpt_bits_uop_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_core_lxcpt_bits_uop_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_lxcpt_bits_uop_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_lxcpt_bits_uop_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_core_lxcpt_bits_uop_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_core_lxcpt_bits_uop_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_lxcpt_bits_uop_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_lxcpt_bits_uop_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_lxcpt_bits_uop_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_lxcpt_bits_uop_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_lxcpt_bits_uop_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_lxcpt_bits_uop_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_lxcpt_bits_uop_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_lxcpt_bits_uop_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_lxcpt_bits_uop_ppred; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_core_lxcpt_bits_uop_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_lxcpt_bits_uop_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_lxcpt_bits_uop_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_lxcpt_bits_uop_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_lxcpt_bits_uop_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_lxcpt_bits_uop_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_lxcpt_bits_uop_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_core_lxcpt_bits_uop_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_lxcpt_bits_uop_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_lxcpt_bits_uop_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_lxcpt_bits_uop_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_core_lxcpt_bits_uop_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_lxcpt_bits_uop_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_core_lxcpt_bits_uop_debug_tsrc; // @[tile.scala 160:20]
  wire [4:0] lsu_io_core_lxcpt_bits_cause; // @[tile.scala 160:20]
  wire [39:0] lsu_io_core_lxcpt_bits_badvaddr; // @[tile.scala 160:20]
  wire [63:0] lsu_io_core_tsc_reg; // @[tile.scala 160:20]
  wire  lsu_io_core_perf_acquire; // @[tile.scala 160:20]
  wire  lsu_io_core_perf_release; // @[tile.scala 160:20]
  wire  lsu_io_core_perf_tlbMiss; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_ready; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_valid; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_valid; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_switch; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_req_bits_0_bits_uop_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_req_bits_0_bits_uop_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_rflag; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_req_bits_0_bits_uop_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_req_bits_0_bits_uop_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_req_bits_0_bits_uop_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_req_bits_0_bits_uop_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_req_bits_0_bits_uop_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_req_bits_0_bits_uop_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_req_bits_0_bits_uop_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_req_bits_0_bits_uop_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_req_bits_0_bits_uop_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_req_bits_0_bits_uop_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_dmem_req_bits_0_bits_uop_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_dmem_req_bits_0_bits_uop_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_dmem_req_bits_0_bits_uop_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_req_bits_0_bits_uop_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_dmem_req_bits_0_bits_uop_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_req_bits_0_bits_uop_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_req_bits_0_bits_uop_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_req_bits_0_bits_uop_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_req_bits_0_bits_uop_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_req_bits_0_bits_uop_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_req_bits_0_bits_uop_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_req_bits_0_bits_uop_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_req_bits_0_bits_uop_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_is_br; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_dmem_req_bits_0_bits_uop_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_req_bits_0_bits_uop_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_dmem_req_bits_0_bits_uop_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_req_bits_0_bits_uop_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_dmem_req_bits_0_bits_uop_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_dmem_req_bits_0_bits_uop_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_req_bits_0_bits_uop_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_dmem_req_bits_0_bits_uop_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_dmem_req_bits_0_bits_uop_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_req_bits_0_bits_uop_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_req_bits_0_bits_uop_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_req_bits_0_bits_uop_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_req_bits_0_bits_uop_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_req_bits_0_bits_uop_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_dmem_req_bits_0_bits_uop_ppred; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_req_bits_0_bits_uop_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_dmem_req_bits_0_bits_uop_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_dmem_req_bits_0_bits_uop_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_req_bits_0_bits_uop_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_req_bits_0_bits_uop_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_req_bits_0_bits_uop_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_req_bits_0_bits_uop_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_req_bits_0_bits_uop_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_req_bits_0_bits_uop_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_req_bits_0_bits_uop_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_req_bits_0_bits_uop_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_uop_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_req_bits_0_bits_uop_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_req_bits_0_bits_uop_debug_tsrc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_dmem_req_bits_0_bits_addr; // @[tile.scala 160:20]
  wire [63:0] lsu_io_dmem_req_bits_0_bits_data; // @[tile.scala 160:20]
  wire  lsu_io_dmem_req_bits_0_bits_is_hella; // @[tile.scala 160:20]
  wire  lsu_io_dmem_s1_kill_0; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_valid; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_switch; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_resp_0_bits_uop_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_resp_0_bits_uop_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_rflag; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_resp_0_bits_uop_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_resp_0_bits_uop_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_resp_0_bits_uop_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_resp_0_bits_uop_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_resp_0_bits_uop_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_resp_0_bits_uop_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_resp_0_bits_uop_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_resp_0_bits_uop_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_resp_0_bits_uop_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_resp_0_bits_uop_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_dmem_resp_0_bits_uop_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_dmem_resp_0_bits_uop_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_dmem_resp_0_bits_uop_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_resp_0_bits_uop_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_dmem_resp_0_bits_uop_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_resp_0_bits_uop_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_resp_0_bits_uop_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_resp_0_bits_uop_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_resp_0_bits_uop_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_resp_0_bits_uop_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_resp_0_bits_uop_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_resp_0_bits_uop_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_resp_0_bits_uop_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_is_br; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_dmem_resp_0_bits_uop_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_resp_0_bits_uop_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_dmem_resp_0_bits_uop_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_resp_0_bits_uop_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_dmem_resp_0_bits_uop_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_dmem_resp_0_bits_uop_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_resp_0_bits_uop_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_dmem_resp_0_bits_uop_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_dmem_resp_0_bits_uop_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_resp_0_bits_uop_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_resp_0_bits_uop_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_resp_0_bits_uop_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_resp_0_bits_uop_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_resp_0_bits_uop_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_dmem_resp_0_bits_uop_ppred; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_resp_0_bits_uop_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_dmem_resp_0_bits_uop_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_dmem_resp_0_bits_uop_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_resp_0_bits_uop_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_resp_0_bits_uop_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_resp_0_bits_uop_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_resp_0_bits_uop_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_resp_0_bits_uop_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_resp_0_bits_uop_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_resp_0_bits_uop_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_resp_0_bits_uop_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_uop_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_resp_0_bits_uop_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_resp_0_bits_uop_debug_tsrc; // @[tile.scala 160:20]
  wire [63:0] lsu_io_dmem_resp_0_bits_data; // @[tile.scala 160:20]
  wire  lsu_io_dmem_resp_0_bits_is_hella; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_valid; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_switch; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_nack_0_bits_uop_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_nack_0_bits_uop_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_rflag; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_nack_0_bits_uop_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_nack_0_bits_uop_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_nack_0_bits_uop_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_nack_0_bits_uop_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_nack_0_bits_uop_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_nack_0_bits_uop_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_nack_0_bits_uop_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_nack_0_bits_uop_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_nack_0_bits_uop_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_nack_0_bits_uop_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_dmem_nack_0_bits_uop_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_dmem_nack_0_bits_uop_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_dmem_nack_0_bits_uop_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_nack_0_bits_uop_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_dmem_nack_0_bits_uop_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_nack_0_bits_uop_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_nack_0_bits_uop_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_nack_0_bits_uop_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_nack_0_bits_uop_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_nack_0_bits_uop_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_nack_0_bits_uop_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_nack_0_bits_uop_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_nack_0_bits_uop_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_is_br; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_dmem_nack_0_bits_uop_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_nack_0_bits_uop_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_dmem_nack_0_bits_uop_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_nack_0_bits_uop_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_dmem_nack_0_bits_uop_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_dmem_nack_0_bits_uop_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_nack_0_bits_uop_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_dmem_nack_0_bits_uop_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_dmem_nack_0_bits_uop_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_nack_0_bits_uop_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_nack_0_bits_uop_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_nack_0_bits_uop_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_nack_0_bits_uop_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_nack_0_bits_uop_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_dmem_nack_0_bits_uop_ppred; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_nack_0_bits_uop_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_dmem_nack_0_bits_uop_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_dmem_nack_0_bits_uop_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_nack_0_bits_uop_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_nack_0_bits_uop_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_nack_0_bits_uop_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_nack_0_bits_uop_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_nack_0_bits_uop_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_nack_0_bits_uop_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_nack_0_bits_uop_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_nack_0_bits_uop_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_uop_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_nack_0_bits_uop_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_nack_0_bits_uop_debug_tsrc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_dmem_nack_0_bits_addr; // @[tile.scala 160:20]
  wire [63:0] lsu_io_dmem_nack_0_bits_data; // @[tile.scala 160:20]
  wire  lsu_io_dmem_nack_0_bits_is_hella; // @[tile.scala 160:20]
  wire [11:0] lsu_io_dmem_brupdate_b1_resolve_mask; // @[tile.scala 160:20]
  wire [11:0] lsu_io_dmem_brupdate_b1_mispredict_mask; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_switch; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_switch_off; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_is_unicore; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_brupdate_b2_uop_shift; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_brupdate_b2_uop_lrs3_rtype; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_rflag; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_wflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_brupdate_b2_uop_prflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_brupdate_b2_uop_pwflag; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_pflag_busy; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_brupdate_b2_uop_stale_pflag; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_brupdate_b2_uop_op1_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_brupdate_b2_uop_op2_sel; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_brupdate_b2_uop_split_num; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_brupdate_b2_uop_self_index; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_brupdate_b2_uop_rob_inst_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_brupdate_b2_uop_address_num; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_brupdate_b2_uop_uopc; // @[tile.scala 160:20]
  wire [31:0] lsu_io_dmem_brupdate_b2_uop_inst; // @[tile.scala 160:20]
  wire [31:0] lsu_io_dmem_brupdate_b2_uop_debug_inst; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_is_rvc; // @[tile.scala 160:20]
  wire [39:0] lsu_io_dmem_brupdate_b2_uop_debug_pc; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_brupdate_b2_uop_iq_type; // @[tile.scala 160:20]
  wire [9:0] lsu_io_dmem_brupdate_b2_uop_fu_code; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_brupdate_b2_uop_ctrl_br_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_brupdate_b2_uop_ctrl_op1_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_brupdate_b2_uop_ctrl_op2_sel; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_brupdate_b2_uop_ctrl_imm_sel; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_brupdate_b2_uop_ctrl_op_fcn; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_ctrl_fcn_dw; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_brupdate_b2_uop_ctrl_csr_cmd; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_ctrl_is_load; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_ctrl_is_sta; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_ctrl_is_std; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_brupdate_b2_uop_ctrl_op3_sel; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_brupdate_b2_uop_iw_state; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_iw_p1_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_iw_p2_poisoned; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_is_br; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_is_jalr; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_is_jal; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_is_sfb; // @[tile.scala 160:20]
  wire [11:0] lsu_io_dmem_brupdate_b2_uop_br_mask; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_brupdate_b2_uop_br_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_dmem_brupdate_b2_uop_ftq_idx; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_edge_inst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_brupdate_b2_uop_pc_lob; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_taken; // @[tile.scala 160:20]
  wire [19:0] lsu_io_dmem_brupdate_b2_uop_imm_packed; // @[tile.scala 160:20]
  wire [11:0] lsu_io_dmem_brupdate_b2_uop_csr_addr; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_brupdate_b2_uop_rob_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_dmem_brupdate_b2_uop_ldq_idx; // @[tile.scala 160:20]
  wire [4:0] lsu_io_dmem_brupdate_b2_uop_stq_idx; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_brupdate_b2_uop_rxq_idx; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_brupdate_b2_uop_pdst; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_brupdate_b2_uop_prs1; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_brupdate_b2_uop_prs2; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_brupdate_b2_uop_prs3; // @[tile.scala 160:20]
  wire [4:0] lsu_io_dmem_brupdate_b2_uop_ppred; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_prs1_busy; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_prs2_busy; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_prs3_busy; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_ppred_busy; // @[tile.scala 160:20]
  wire [6:0] lsu_io_dmem_brupdate_b2_uop_stale_pdst; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_exception; // @[tile.scala 160:20]
  wire [63:0] lsu_io_dmem_brupdate_b2_uop_exc_cause; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_bypassable; // @[tile.scala 160:20]
  wire [4:0] lsu_io_dmem_brupdate_b2_uop_mem_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_brupdate_b2_uop_mem_size; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_mem_signed; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_is_fence; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_is_fencei; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_is_amo; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_uses_ldq; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_uses_stq; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_is_sys_pc2epc; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_is_unique; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_flush_on_commit; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_ldst_is_rs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_brupdate_b2_uop_ldst; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_brupdate_b2_uop_lrs1; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_brupdate_b2_uop_lrs2; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_brupdate_b2_uop_lrs3; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_ldst_val; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_brupdate_b2_uop_dst_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_brupdate_b2_uop_lrs1_rtype; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_brupdate_b2_uop_lrs2_rtype; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_frs3_en; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_fp_val; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_fp_single; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_xcpt_pf_if; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_xcpt_ae_if; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_xcpt_ma_if; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_bp_debug_if; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_uop_bp_xcpt_if; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_brupdate_b2_uop_debug_fsrc; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_brupdate_b2_uop_debug_tsrc; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_valid; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_mispredict; // @[tile.scala 160:20]
  wire  lsu_io_dmem_brupdate_b2_taken; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_brupdate_b2_cfi_type; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_brupdate_b2_pc_sel; // @[tile.scala 160:20]
  wire [39:0] lsu_io_dmem_brupdate_b2_jalr_target; // @[tile.scala 160:20]
  wire [31:0] lsu_io_dmem_brupdate_b2_target_offset; // @[tile.scala 160:20]
  wire  lsu_io_dmem_exception; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_rob_pnr_idx; // @[tile.scala 160:20]
  wire [5:0] lsu_io_dmem_rob_head_idx; // @[tile.scala 160:20]
  wire  lsu_io_dmem_release_ready; // @[tile.scala 160:20]
  wire  lsu_io_dmem_release_valid; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_release_bits_opcode; // @[tile.scala 160:20]
  wire [2:0] lsu_io_dmem_release_bits_param; // @[tile.scala 160:20]
  wire [3:0] lsu_io_dmem_release_bits_size; // @[tile.scala 160:20]
  wire [1:0] lsu_io_dmem_release_bits_source; // @[tile.scala 160:20]
  wire [31:0] lsu_io_dmem_release_bits_address; // @[tile.scala 160:20]
  wire [63:0] lsu_io_dmem_release_bits_data; // @[tile.scala 160:20]
  wire  lsu_io_dmem_release_bits_corrupt; // @[tile.scala 160:20]
  wire  lsu_io_dmem_force_order; // @[tile.scala 160:20]
  wire  lsu_io_dmem_ordered; // @[tile.scala 160:20]
  wire  lsu_io_dmem_perf_acquire; // @[tile.scala 160:20]
  wire  lsu_io_dmem_perf_release; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_req_ready; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_req_valid; // @[tile.scala 160:20]
  wire [39:0] lsu_io_hellacache_req_bits_addr; // @[tile.scala 160:20]
  wire [6:0] lsu_io_hellacache_req_bits_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_hellacache_req_bits_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_hellacache_req_bits_size; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_req_bits_signed; // @[tile.scala 160:20]
  wire [1:0] lsu_io_hellacache_req_bits_dprv; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_req_bits_phys; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_req_bits_no_alloc; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_req_bits_no_xcpt; // @[tile.scala 160:20]
  wire [63:0] lsu_io_hellacache_req_bits_data; // @[tile.scala 160:20]
  wire [7:0] lsu_io_hellacache_req_bits_mask; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_s1_kill; // @[tile.scala 160:20]
  wire [63:0] lsu_io_hellacache_s1_data_data; // @[tile.scala 160:20]
  wire [7:0] lsu_io_hellacache_s1_data_mask; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_s2_nack; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_s2_nack_cause_raw; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_s2_kill; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_s2_uncached; // @[tile.scala 160:20]
  wire [31:0] lsu_io_hellacache_s2_paddr; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_resp_valid; // @[tile.scala 160:20]
  wire [39:0] lsu_io_hellacache_resp_bits_addr; // @[tile.scala 160:20]
  wire [6:0] lsu_io_hellacache_resp_bits_tag; // @[tile.scala 160:20]
  wire [4:0] lsu_io_hellacache_resp_bits_cmd; // @[tile.scala 160:20]
  wire [1:0] lsu_io_hellacache_resp_bits_size; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_resp_bits_signed; // @[tile.scala 160:20]
  wire [1:0] lsu_io_hellacache_resp_bits_dprv; // @[tile.scala 160:20]
  wire [63:0] lsu_io_hellacache_resp_bits_data; // @[tile.scala 160:20]
  wire [7:0] lsu_io_hellacache_resp_bits_mask; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_resp_bits_replay; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_resp_bits_has_data; // @[tile.scala 160:20]
  wire [63:0] lsu_io_hellacache_resp_bits_data_word_bypass; // @[tile.scala 160:20]
  wire [63:0] lsu_io_hellacache_resp_bits_data_raw; // @[tile.scala 160:20]
  wire [63:0] lsu_io_hellacache_resp_bits_store_data; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_replay_next; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_s2_xcpt_ma_ld; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_s2_xcpt_ma_st; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_s2_xcpt_pf_ld; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_s2_xcpt_pf_st; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_s2_xcpt_ae_ld; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_s2_xcpt_ae_st; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_ordered; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_perf_acquire; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_perf_release; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_perf_grant; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_perf_tlbMiss; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_perf_blocked; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_perf_canAcceptStoreThenLoad; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_perf_canAcceptStoreThenRMW; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_perf_canAcceptLoadThenLoad; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_perf_storeBufferEmptyAfterLoad; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_perf_storeBufferEmptyAfterStore; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_keep_clock_enabled; // @[tile.scala 160:20]
  wire  lsu_io_hellacache_clock_enabled; // @[tile.scala 160:20]
  wire  ptw_clock; // @[tile.scala 230:20]
  wire  ptw_reset; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_req_ready; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_req_valid; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_req_bits_valid; // @[tile.scala 230:20]
  wire [26:0] ptw_io_requestor_0_req_bits_bits_addr; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_resp_valid; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_resp_bits_ae; // @[tile.scala 230:20]
  wire [53:0] ptw_io_requestor_0_resp_bits_pte_ppn; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_resp_bits_pte_reserved_for_software; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_resp_bits_pte_d; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_resp_bits_pte_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_resp_bits_pte_g; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_resp_bits_pte_u; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_resp_bits_pte_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_resp_bits_pte_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_resp_bits_pte_r; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_resp_bits_pte_v; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_resp_bits_level; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_resp_bits_fragmented_superpage; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_resp_bits_homogeneous; // @[tile.scala 230:20]
  wire [3:0] ptw_io_requestor_0_ptbr_mode; // @[tile.scala 230:20]
  wire [15:0] ptw_io_requestor_0_ptbr_asid; // @[tile.scala 230:20]
  wire [43:0] ptw_io_requestor_0_ptbr_ppn; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_status_debug; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_status_cease; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_status_wfi; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_0_status_isa; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_status_dprv; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_status_prv; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_status_sd; // @[tile.scala 230:20]
  wire [26:0] ptw_io_requestor_0_status_zero2; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_status_sxl; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_status_uxl; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_status_sd_rv32; // @[tile.scala 230:20]
  wire [7:0] ptw_io_requestor_0_status_zero1; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_status_tsr; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_status_tw; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_status_tvm; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_status_mxr; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_status_sum; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_status_mprv; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_status_xs; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_status_fs; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_status_mpp; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_status_vs; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_status_spp; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_status_mpie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_status_hpie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_status_spie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_status_upie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_status_mie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_status_hie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_status_sie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_status_uie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_0_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_pmp_0_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_pmp_0_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_0_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_0_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_0_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_0_pmp_0_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_0_pmp_0_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_1_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_pmp_1_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_pmp_1_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_1_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_1_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_1_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_0_pmp_1_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_0_pmp_1_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_2_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_pmp_2_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_pmp_2_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_2_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_2_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_2_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_0_pmp_2_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_0_pmp_2_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_3_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_pmp_3_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_pmp_3_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_3_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_3_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_3_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_0_pmp_3_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_0_pmp_3_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_4_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_pmp_4_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_pmp_4_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_4_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_4_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_4_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_0_pmp_4_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_0_pmp_4_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_5_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_pmp_5_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_pmp_5_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_5_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_5_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_5_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_0_pmp_5_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_0_pmp_5_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_6_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_pmp_6_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_pmp_6_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_6_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_6_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_6_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_0_pmp_6_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_0_pmp_6_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_7_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_pmp_7_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_0_pmp_7_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_7_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_7_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_pmp_7_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_0_pmp_7_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_0_pmp_7_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_0_customCSRs_csrs_0_wen; // @[tile.scala 230:20]
  wire [63:0] ptw_io_requestor_0_customCSRs_csrs_0_wdata; // @[tile.scala 230:20]
  wire [63:0] ptw_io_requestor_0_customCSRs_csrs_0_value; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_req_ready; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_req_valid; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_req_bits_valid; // @[tile.scala 230:20]
  wire [26:0] ptw_io_requestor_1_req_bits_bits_addr; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_resp_valid; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_resp_bits_ae; // @[tile.scala 230:20]
  wire [53:0] ptw_io_requestor_1_resp_bits_pte_ppn; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_resp_bits_pte_reserved_for_software; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_resp_bits_pte_d; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_resp_bits_pte_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_resp_bits_pte_g; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_resp_bits_pte_u; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_resp_bits_pte_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_resp_bits_pte_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_resp_bits_pte_r; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_resp_bits_pte_v; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_resp_bits_level; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_resp_bits_fragmented_superpage; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_resp_bits_homogeneous; // @[tile.scala 230:20]
  wire [3:0] ptw_io_requestor_1_ptbr_mode; // @[tile.scala 230:20]
  wire [15:0] ptw_io_requestor_1_ptbr_asid; // @[tile.scala 230:20]
  wire [43:0] ptw_io_requestor_1_ptbr_ppn; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_status_debug; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_status_cease; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_status_wfi; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_1_status_isa; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_status_dprv; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_status_prv; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_status_sd; // @[tile.scala 230:20]
  wire [26:0] ptw_io_requestor_1_status_zero2; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_status_sxl; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_status_uxl; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_status_sd_rv32; // @[tile.scala 230:20]
  wire [7:0] ptw_io_requestor_1_status_zero1; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_status_tsr; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_status_tw; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_status_tvm; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_status_mxr; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_status_sum; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_status_mprv; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_status_xs; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_status_fs; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_status_mpp; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_status_vs; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_status_spp; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_status_mpie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_status_hpie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_status_spie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_status_upie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_status_mie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_status_hie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_status_sie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_status_uie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_0_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_pmp_0_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_pmp_0_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_0_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_0_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_0_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_1_pmp_0_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_1_pmp_0_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_1_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_pmp_1_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_pmp_1_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_1_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_1_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_1_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_1_pmp_1_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_1_pmp_1_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_2_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_pmp_2_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_pmp_2_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_2_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_2_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_2_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_1_pmp_2_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_1_pmp_2_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_3_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_pmp_3_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_pmp_3_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_3_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_3_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_3_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_1_pmp_3_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_1_pmp_3_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_4_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_pmp_4_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_pmp_4_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_4_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_4_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_4_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_1_pmp_4_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_1_pmp_4_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_5_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_pmp_5_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_pmp_5_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_5_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_5_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_5_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_1_pmp_5_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_1_pmp_5_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_6_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_pmp_6_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_pmp_6_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_6_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_6_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_6_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_1_pmp_6_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_1_pmp_6_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_7_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_pmp_7_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_1_pmp_7_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_7_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_7_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_pmp_7_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_1_pmp_7_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_1_pmp_7_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_1_customCSRs_csrs_0_wen; // @[tile.scala 230:20]
  wire [63:0] ptw_io_requestor_1_customCSRs_csrs_0_wdata; // @[tile.scala 230:20]
  wire [63:0] ptw_io_requestor_1_customCSRs_csrs_0_value; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_req_ready; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_req_valid; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_req_bits_valid; // @[tile.scala 230:20]
  wire [26:0] ptw_io_requestor_2_req_bits_bits_addr; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_resp_valid; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_resp_bits_ae; // @[tile.scala 230:20]
  wire [53:0] ptw_io_requestor_2_resp_bits_pte_ppn; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_resp_bits_pte_reserved_for_software; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_resp_bits_pte_d; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_resp_bits_pte_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_resp_bits_pte_g; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_resp_bits_pte_u; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_resp_bits_pte_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_resp_bits_pte_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_resp_bits_pte_r; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_resp_bits_pte_v; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_resp_bits_level; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_resp_bits_fragmented_superpage; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_resp_bits_homogeneous; // @[tile.scala 230:20]
  wire [3:0] ptw_io_requestor_2_ptbr_mode; // @[tile.scala 230:20]
  wire [15:0] ptw_io_requestor_2_ptbr_asid; // @[tile.scala 230:20]
  wire [43:0] ptw_io_requestor_2_ptbr_ppn; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_status_debug; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_status_cease; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_status_wfi; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_2_status_isa; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_status_dprv; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_status_prv; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_status_sd; // @[tile.scala 230:20]
  wire [26:0] ptw_io_requestor_2_status_zero2; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_status_sxl; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_status_uxl; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_status_sd_rv32; // @[tile.scala 230:20]
  wire [7:0] ptw_io_requestor_2_status_zero1; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_status_tsr; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_status_tw; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_status_tvm; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_status_mxr; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_status_sum; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_status_mprv; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_status_xs; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_status_fs; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_status_mpp; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_status_vs; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_status_spp; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_status_mpie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_status_hpie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_status_spie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_status_upie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_status_mie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_status_hie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_status_sie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_status_uie; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_0_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_pmp_0_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_pmp_0_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_0_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_0_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_0_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_2_pmp_0_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_2_pmp_0_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_1_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_pmp_1_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_pmp_1_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_1_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_1_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_1_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_2_pmp_1_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_2_pmp_1_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_2_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_pmp_2_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_pmp_2_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_2_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_2_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_2_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_2_pmp_2_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_2_pmp_2_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_3_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_pmp_3_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_pmp_3_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_3_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_3_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_3_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_2_pmp_3_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_2_pmp_3_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_4_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_pmp_4_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_pmp_4_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_4_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_4_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_4_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_2_pmp_4_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_2_pmp_4_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_5_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_pmp_5_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_pmp_5_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_5_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_5_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_5_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_2_pmp_5_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_2_pmp_5_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_6_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_pmp_6_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_pmp_6_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_6_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_6_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_6_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_2_pmp_6_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_2_pmp_6_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_7_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_pmp_7_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_requestor_2_pmp_7_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_7_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_7_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_pmp_7_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_requestor_2_pmp_7_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_requestor_2_pmp_7_mask; // @[tile.scala 230:20]
  wire  ptw_io_requestor_2_customCSRs_csrs_0_wen; // @[tile.scala 230:20]
  wire [63:0] ptw_io_requestor_2_customCSRs_csrs_0_wdata; // @[tile.scala 230:20]
  wire [63:0] ptw_io_requestor_2_customCSRs_csrs_0_value; // @[tile.scala 230:20]
  wire  ptw_io_mem_req_ready; // @[tile.scala 230:20]
  wire  ptw_io_mem_req_valid; // @[tile.scala 230:20]
  wire [39:0] ptw_io_mem_req_bits_addr; // @[tile.scala 230:20]
  wire [6:0] ptw_io_mem_req_bits_tag; // @[tile.scala 230:20]
  wire [4:0] ptw_io_mem_req_bits_cmd; // @[tile.scala 230:20]
  wire [1:0] ptw_io_mem_req_bits_size; // @[tile.scala 230:20]
  wire  ptw_io_mem_req_bits_signed; // @[tile.scala 230:20]
  wire [1:0] ptw_io_mem_req_bits_dprv; // @[tile.scala 230:20]
  wire  ptw_io_mem_req_bits_phys; // @[tile.scala 230:20]
  wire  ptw_io_mem_req_bits_no_alloc; // @[tile.scala 230:20]
  wire  ptw_io_mem_req_bits_no_xcpt; // @[tile.scala 230:20]
  wire [63:0] ptw_io_mem_req_bits_data; // @[tile.scala 230:20]
  wire [7:0] ptw_io_mem_req_bits_mask; // @[tile.scala 230:20]
  wire  ptw_io_mem_s1_kill; // @[tile.scala 230:20]
  wire [63:0] ptw_io_mem_s1_data_data; // @[tile.scala 230:20]
  wire [7:0] ptw_io_mem_s1_data_mask; // @[tile.scala 230:20]
  wire  ptw_io_mem_s2_nack; // @[tile.scala 230:20]
  wire  ptw_io_mem_s2_nack_cause_raw; // @[tile.scala 230:20]
  wire  ptw_io_mem_s2_kill; // @[tile.scala 230:20]
  wire  ptw_io_mem_s2_uncached; // @[tile.scala 230:20]
  wire [31:0] ptw_io_mem_s2_paddr; // @[tile.scala 230:20]
  wire  ptw_io_mem_resp_valid; // @[tile.scala 230:20]
  wire [39:0] ptw_io_mem_resp_bits_addr; // @[tile.scala 230:20]
  wire [6:0] ptw_io_mem_resp_bits_tag; // @[tile.scala 230:20]
  wire [4:0] ptw_io_mem_resp_bits_cmd; // @[tile.scala 230:20]
  wire [1:0] ptw_io_mem_resp_bits_size; // @[tile.scala 230:20]
  wire  ptw_io_mem_resp_bits_signed; // @[tile.scala 230:20]
  wire [1:0] ptw_io_mem_resp_bits_dprv; // @[tile.scala 230:20]
  wire [63:0] ptw_io_mem_resp_bits_data; // @[tile.scala 230:20]
  wire [7:0] ptw_io_mem_resp_bits_mask; // @[tile.scala 230:20]
  wire  ptw_io_mem_resp_bits_replay; // @[tile.scala 230:20]
  wire  ptw_io_mem_resp_bits_has_data; // @[tile.scala 230:20]
  wire [63:0] ptw_io_mem_resp_bits_data_word_bypass; // @[tile.scala 230:20]
  wire [63:0] ptw_io_mem_resp_bits_data_raw; // @[tile.scala 230:20]
  wire [63:0] ptw_io_mem_resp_bits_store_data; // @[tile.scala 230:20]
  wire  ptw_io_mem_replay_next; // @[tile.scala 230:20]
  wire  ptw_io_mem_s2_xcpt_ma_ld; // @[tile.scala 230:20]
  wire  ptw_io_mem_s2_xcpt_ma_st; // @[tile.scala 230:20]
  wire  ptw_io_mem_s2_xcpt_pf_ld; // @[tile.scala 230:20]
  wire  ptw_io_mem_s2_xcpt_pf_st; // @[tile.scala 230:20]
  wire  ptw_io_mem_s2_xcpt_ae_ld; // @[tile.scala 230:20]
  wire  ptw_io_mem_s2_xcpt_ae_st; // @[tile.scala 230:20]
  wire  ptw_io_mem_ordered; // @[tile.scala 230:20]
  wire  ptw_io_mem_perf_acquire; // @[tile.scala 230:20]
  wire  ptw_io_mem_perf_release; // @[tile.scala 230:20]
  wire  ptw_io_mem_perf_grant; // @[tile.scala 230:20]
  wire  ptw_io_mem_perf_tlbMiss; // @[tile.scala 230:20]
  wire  ptw_io_mem_perf_blocked; // @[tile.scala 230:20]
  wire  ptw_io_mem_perf_canAcceptStoreThenLoad; // @[tile.scala 230:20]
  wire  ptw_io_mem_perf_canAcceptStoreThenRMW; // @[tile.scala 230:20]
  wire  ptw_io_mem_perf_canAcceptLoadThenLoad; // @[tile.scala 230:20]
  wire  ptw_io_mem_perf_storeBufferEmptyAfterLoad; // @[tile.scala 230:20]
  wire  ptw_io_mem_perf_storeBufferEmptyAfterStore; // @[tile.scala 230:20]
  wire  ptw_io_mem_keep_clock_enabled; // @[tile.scala 230:20]
  wire  ptw_io_mem_clock_enabled; // @[tile.scala 230:20]
  wire [3:0] ptw_io_dpath_ptbr_mode; // @[tile.scala 230:20]
  wire [15:0] ptw_io_dpath_ptbr_asid; // @[tile.scala 230:20]
  wire [43:0] ptw_io_dpath_ptbr_ppn; // @[tile.scala 230:20]
  wire  ptw_io_dpath_sfence_valid; // @[tile.scala 230:20]
  wire  ptw_io_dpath_sfence_bits_rs1; // @[tile.scala 230:20]
  wire  ptw_io_dpath_sfence_bits_rs2; // @[tile.scala 230:20]
  wire [38:0] ptw_io_dpath_sfence_bits_addr; // @[tile.scala 230:20]
  wire  ptw_io_dpath_sfence_bits_asid; // @[tile.scala 230:20]
  wire  ptw_io_dpath_status_debug; // @[tile.scala 230:20]
  wire  ptw_io_dpath_status_cease; // @[tile.scala 230:20]
  wire  ptw_io_dpath_status_wfi; // @[tile.scala 230:20]
  wire [31:0] ptw_io_dpath_status_isa; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_status_dprv; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_status_prv; // @[tile.scala 230:20]
  wire  ptw_io_dpath_status_sd; // @[tile.scala 230:20]
  wire [26:0] ptw_io_dpath_status_zero2; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_status_sxl; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_status_uxl; // @[tile.scala 230:20]
  wire  ptw_io_dpath_status_sd_rv32; // @[tile.scala 230:20]
  wire [7:0] ptw_io_dpath_status_zero1; // @[tile.scala 230:20]
  wire  ptw_io_dpath_status_tsr; // @[tile.scala 230:20]
  wire  ptw_io_dpath_status_tw; // @[tile.scala 230:20]
  wire  ptw_io_dpath_status_tvm; // @[tile.scala 230:20]
  wire  ptw_io_dpath_status_mxr; // @[tile.scala 230:20]
  wire  ptw_io_dpath_status_sum; // @[tile.scala 230:20]
  wire  ptw_io_dpath_status_mprv; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_status_xs; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_status_fs; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_status_mpp; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_status_vs; // @[tile.scala 230:20]
  wire  ptw_io_dpath_status_spp; // @[tile.scala 230:20]
  wire  ptw_io_dpath_status_mpie; // @[tile.scala 230:20]
  wire  ptw_io_dpath_status_hpie; // @[tile.scala 230:20]
  wire  ptw_io_dpath_status_spie; // @[tile.scala 230:20]
  wire  ptw_io_dpath_status_upie; // @[tile.scala 230:20]
  wire  ptw_io_dpath_status_mie; // @[tile.scala 230:20]
  wire  ptw_io_dpath_status_hie; // @[tile.scala 230:20]
  wire  ptw_io_dpath_status_sie; // @[tile.scala 230:20]
  wire  ptw_io_dpath_status_uie; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_0_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_pmp_0_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_pmp_0_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_0_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_0_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_0_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_dpath_pmp_0_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_dpath_pmp_0_mask; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_1_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_pmp_1_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_pmp_1_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_1_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_1_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_1_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_dpath_pmp_1_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_dpath_pmp_1_mask; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_2_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_pmp_2_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_pmp_2_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_2_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_2_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_2_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_dpath_pmp_2_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_dpath_pmp_2_mask; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_3_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_pmp_3_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_pmp_3_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_3_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_3_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_3_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_dpath_pmp_3_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_dpath_pmp_3_mask; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_4_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_pmp_4_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_pmp_4_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_4_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_4_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_4_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_dpath_pmp_4_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_dpath_pmp_4_mask; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_5_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_pmp_5_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_pmp_5_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_5_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_5_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_5_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_dpath_pmp_5_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_dpath_pmp_5_mask; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_6_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_pmp_6_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_pmp_6_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_6_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_6_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_6_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_dpath_pmp_6_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_dpath_pmp_6_mask; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_7_cfg_l; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_pmp_7_cfg_res; // @[tile.scala 230:20]
  wire [1:0] ptw_io_dpath_pmp_7_cfg_a; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_7_cfg_x; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_7_cfg_w; // @[tile.scala 230:20]
  wire  ptw_io_dpath_pmp_7_cfg_r; // @[tile.scala 230:20]
  wire [29:0] ptw_io_dpath_pmp_7_addr; // @[tile.scala 230:20]
  wire [31:0] ptw_io_dpath_pmp_7_mask; // @[tile.scala 230:20]
  wire  ptw_io_dpath_perf_l2miss; // @[tile.scala 230:20]
  wire  ptw_io_dpath_perf_l2hit; // @[tile.scala 230:20]
  wire  ptw_io_dpath_perf_pte_miss; // @[tile.scala 230:20]
  wire  ptw_io_dpath_perf_pte_hit; // @[tile.scala 230:20]
  wire  ptw_io_dpath_customCSRs_csrs_0_wen; // @[tile.scala 230:20]
  wire [63:0] ptw_io_dpath_customCSRs_csrs_0_wdata; // @[tile.scala 230:20]
  wire [63:0] ptw_io_dpath_customCSRs_csrs_0_value; // @[tile.scala 230:20]
  wire  ptw_io_dpath_clock_enabled; // @[tile.scala 230:20]
  wire  hellaCacheArb_clock; // @[tile.scala 236:29]
  wire  hellaCacheArb_reset; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_req_ready; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_req_valid; // @[tile.scala 236:29]
  wire [39:0] hellaCacheArb_io_requestor_0_req_bits_addr; // @[tile.scala 236:29]
  wire [6:0] hellaCacheArb_io_requestor_0_req_bits_tag; // @[tile.scala 236:29]
  wire [4:0] hellaCacheArb_io_requestor_0_req_bits_cmd; // @[tile.scala 236:29]
  wire [1:0] hellaCacheArb_io_requestor_0_req_bits_size; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_req_bits_signed; // @[tile.scala 236:29]
  wire [1:0] hellaCacheArb_io_requestor_0_req_bits_dprv; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_req_bits_phys; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_req_bits_no_alloc; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_req_bits_no_xcpt; // @[tile.scala 236:29]
  wire [63:0] hellaCacheArb_io_requestor_0_req_bits_data; // @[tile.scala 236:29]
  wire [7:0] hellaCacheArb_io_requestor_0_req_bits_mask; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_s1_kill; // @[tile.scala 236:29]
  wire [63:0] hellaCacheArb_io_requestor_0_s1_data_data; // @[tile.scala 236:29]
  wire [7:0] hellaCacheArb_io_requestor_0_s1_data_mask; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_s2_nack; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_s2_nack_cause_raw; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_s2_kill; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_s2_uncached; // @[tile.scala 236:29]
  wire [31:0] hellaCacheArb_io_requestor_0_s2_paddr; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_resp_valid; // @[tile.scala 236:29]
  wire [39:0] hellaCacheArb_io_requestor_0_resp_bits_addr; // @[tile.scala 236:29]
  wire [6:0] hellaCacheArb_io_requestor_0_resp_bits_tag; // @[tile.scala 236:29]
  wire [4:0] hellaCacheArb_io_requestor_0_resp_bits_cmd; // @[tile.scala 236:29]
  wire [1:0] hellaCacheArb_io_requestor_0_resp_bits_size; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_resp_bits_signed; // @[tile.scala 236:29]
  wire [1:0] hellaCacheArb_io_requestor_0_resp_bits_dprv; // @[tile.scala 236:29]
  wire [63:0] hellaCacheArb_io_requestor_0_resp_bits_data; // @[tile.scala 236:29]
  wire [7:0] hellaCacheArb_io_requestor_0_resp_bits_mask; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_resp_bits_replay; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_resp_bits_has_data; // @[tile.scala 236:29]
  wire [63:0] hellaCacheArb_io_requestor_0_resp_bits_data_word_bypass; // @[tile.scala 236:29]
  wire [63:0] hellaCacheArb_io_requestor_0_resp_bits_data_raw; // @[tile.scala 236:29]
  wire [63:0] hellaCacheArb_io_requestor_0_resp_bits_store_data; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_replay_next; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_s2_xcpt_ma_ld; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_s2_xcpt_ma_st; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_s2_xcpt_pf_ld; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_s2_xcpt_pf_st; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_s2_xcpt_ae_ld; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_s2_xcpt_ae_st; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_ordered; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_perf_acquire; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_perf_release; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_perf_grant; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_perf_tlbMiss; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_perf_blocked; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_perf_canAcceptStoreThenLoad; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_perf_canAcceptStoreThenRMW; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_perf_canAcceptLoadThenLoad; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_perf_storeBufferEmptyAfterLoad; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_perf_storeBufferEmptyAfterStore; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_keep_clock_enabled; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_requestor_0_clock_enabled; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_req_ready; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_req_valid; // @[tile.scala 236:29]
  wire [39:0] hellaCacheArb_io_mem_req_bits_addr; // @[tile.scala 236:29]
  wire [6:0] hellaCacheArb_io_mem_req_bits_tag; // @[tile.scala 236:29]
  wire [4:0] hellaCacheArb_io_mem_req_bits_cmd; // @[tile.scala 236:29]
  wire [1:0] hellaCacheArb_io_mem_req_bits_size; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_req_bits_signed; // @[tile.scala 236:29]
  wire [1:0] hellaCacheArb_io_mem_req_bits_dprv; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_req_bits_phys; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_req_bits_no_alloc; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_req_bits_no_xcpt; // @[tile.scala 236:29]
  wire [63:0] hellaCacheArb_io_mem_req_bits_data; // @[tile.scala 236:29]
  wire [7:0] hellaCacheArb_io_mem_req_bits_mask; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_s1_kill; // @[tile.scala 236:29]
  wire [63:0] hellaCacheArb_io_mem_s1_data_data; // @[tile.scala 236:29]
  wire [7:0] hellaCacheArb_io_mem_s1_data_mask; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_s2_nack; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_s2_nack_cause_raw; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_s2_kill; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_s2_uncached; // @[tile.scala 236:29]
  wire [31:0] hellaCacheArb_io_mem_s2_paddr; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_resp_valid; // @[tile.scala 236:29]
  wire [39:0] hellaCacheArb_io_mem_resp_bits_addr; // @[tile.scala 236:29]
  wire [6:0] hellaCacheArb_io_mem_resp_bits_tag; // @[tile.scala 236:29]
  wire [4:0] hellaCacheArb_io_mem_resp_bits_cmd; // @[tile.scala 236:29]
  wire [1:0] hellaCacheArb_io_mem_resp_bits_size; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_resp_bits_signed; // @[tile.scala 236:29]
  wire [1:0] hellaCacheArb_io_mem_resp_bits_dprv; // @[tile.scala 236:29]
  wire [63:0] hellaCacheArb_io_mem_resp_bits_data; // @[tile.scala 236:29]
  wire [7:0] hellaCacheArb_io_mem_resp_bits_mask; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_resp_bits_replay; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_resp_bits_has_data; // @[tile.scala 236:29]
  wire [63:0] hellaCacheArb_io_mem_resp_bits_data_word_bypass; // @[tile.scala 236:29]
  wire [63:0] hellaCacheArb_io_mem_resp_bits_data_raw; // @[tile.scala 236:29]
  wire [63:0] hellaCacheArb_io_mem_resp_bits_store_data; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_replay_next; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_s2_xcpt_ma_ld; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_s2_xcpt_ma_st; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_s2_xcpt_pf_ld; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_s2_xcpt_pf_st; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_s2_xcpt_ae_ld; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_s2_xcpt_ae_st; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_ordered; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_perf_acquire; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_perf_release; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_perf_grant; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_perf_tlbMiss; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_perf_blocked; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_perf_canAcceptStoreThenLoad; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_perf_canAcceptStoreThenRMW; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_perf_canAcceptLoadThenLoad; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_perf_storeBufferEmptyAfterLoad; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_perf_storeBufferEmptyAfterStore; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_keep_clock_enabled; // @[tile.scala 236:29]
  wire  hellaCacheArb_io_mem_clock_enabled; // @[tile.scala 236:29]
  TLXbar_7 tlMasterXbar ( // @[BaseTile.scala 195:42]
    .clock(tlMasterXbar_clock),
    .reset(tlMasterXbar_reset),
    .auto_in_1_a_ready(tlMasterXbar_auto_in_1_a_ready),
    .auto_in_1_a_valid(tlMasterXbar_auto_in_1_a_valid),
    .auto_in_1_a_bits_opcode(tlMasterXbar_auto_in_1_a_bits_opcode),
    .auto_in_1_a_bits_param(tlMasterXbar_auto_in_1_a_bits_param),
    .auto_in_1_a_bits_size(tlMasterXbar_auto_in_1_a_bits_size),
    .auto_in_1_a_bits_source(tlMasterXbar_auto_in_1_a_bits_source),
    .auto_in_1_a_bits_address(tlMasterXbar_auto_in_1_a_bits_address),
    .auto_in_1_a_bits_mask(tlMasterXbar_auto_in_1_a_bits_mask),
    .auto_in_1_a_bits_data(tlMasterXbar_auto_in_1_a_bits_data),
    .auto_in_1_a_bits_corrupt(tlMasterXbar_auto_in_1_a_bits_corrupt),
    .auto_in_1_d_ready(tlMasterXbar_auto_in_1_d_ready),
    .auto_in_1_d_valid(tlMasterXbar_auto_in_1_d_valid),
    .auto_in_1_d_bits_opcode(tlMasterXbar_auto_in_1_d_bits_opcode),
    .auto_in_1_d_bits_param(tlMasterXbar_auto_in_1_d_bits_param),
    .auto_in_1_d_bits_size(tlMasterXbar_auto_in_1_d_bits_size),
    .auto_in_1_d_bits_source(tlMasterXbar_auto_in_1_d_bits_source),
    .auto_in_1_d_bits_sink(tlMasterXbar_auto_in_1_d_bits_sink),
    .auto_in_1_d_bits_denied(tlMasterXbar_auto_in_1_d_bits_denied),
    .auto_in_1_d_bits_data(tlMasterXbar_auto_in_1_d_bits_data),
    .auto_in_1_d_bits_corrupt(tlMasterXbar_auto_in_1_d_bits_corrupt),
    .auto_in_0_a_ready(tlMasterXbar_auto_in_0_a_ready),
    .auto_in_0_a_valid(tlMasterXbar_auto_in_0_a_valid),
    .auto_in_0_a_bits_opcode(tlMasterXbar_auto_in_0_a_bits_opcode),
    .auto_in_0_a_bits_param(tlMasterXbar_auto_in_0_a_bits_param),
    .auto_in_0_a_bits_size(tlMasterXbar_auto_in_0_a_bits_size),
    .auto_in_0_a_bits_source(tlMasterXbar_auto_in_0_a_bits_source),
    .auto_in_0_a_bits_address(tlMasterXbar_auto_in_0_a_bits_address),
    .auto_in_0_a_bits_mask(tlMasterXbar_auto_in_0_a_bits_mask),
    .auto_in_0_a_bits_data(tlMasterXbar_auto_in_0_a_bits_data),
    .auto_in_0_a_bits_corrupt(tlMasterXbar_auto_in_0_a_bits_corrupt),
    .auto_in_0_b_ready(tlMasterXbar_auto_in_0_b_ready),
    .auto_in_0_b_valid(tlMasterXbar_auto_in_0_b_valid),
    .auto_in_0_b_bits_opcode(tlMasterXbar_auto_in_0_b_bits_opcode),
    .auto_in_0_b_bits_param(tlMasterXbar_auto_in_0_b_bits_param),
    .auto_in_0_b_bits_size(tlMasterXbar_auto_in_0_b_bits_size),
    .auto_in_0_b_bits_source(tlMasterXbar_auto_in_0_b_bits_source),
    .auto_in_0_b_bits_address(tlMasterXbar_auto_in_0_b_bits_address),
    .auto_in_0_b_bits_mask(tlMasterXbar_auto_in_0_b_bits_mask),
    .auto_in_0_b_bits_data(tlMasterXbar_auto_in_0_b_bits_data),
    .auto_in_0_b_bits_corrupt(tlMasterXbar_auto_in_0_b_bits_corrupt),
    .auto_in_0_c_ready(tlMasterXbar_auto_in_0_c_ready),
    .auto_in_0_c_valid(tlMasterXbar_auto_in_0_c_valid),
    .auto_in_0_c_bits_opcode(tlMasterXbar_auto_in_0_c_bits_opcode),
    .auto_in_0_c_bits_param(tlMasterXbar_auto_in_0_c_bits_param),
    .auto_in_0_c_bits_size(tlMasterXbar_auto_in_0_c_bits_size),
    .auto_in_0_c_bits_source(tlMasterXbar_auto_in_0_c_bits_source),
    .auto_in_0_c_bits_address(tlMasterXbar_auto_in_0_c_bits_address),
    .auto_in_0_c_bits_data(tlMasterXbar_auto_in_0_c_bits_data),
    .auto_in_0_c_bits_corrupt(tlMasterXbar_auto_in_0_c_bits_corrupt),
    .auto_in_0_d_ready(tlMasterXbar_auto_in_0_d_ready),
    .auto_in_0_d_valid(tlMasterXbar_auto_in_0_d_valid),
    .auto_in_0_d_bits_opcode(tlMasterXbar_auto_in_0_d_bits_opcode),
    .auto_in_0_d_bits_param(tlMasterXbar_auto_in_0_d_bits_param),
    .auto_in_0_d_bits_size(tlMasterXbar_auto_in_0_d_bits_size),
    .auto_in_0_d_bits_source(tlMasterXbar_auto_in_0_d_bits_source),
    .auto_in_0_d_bits_sink(tlMasterXbar_auto_in_0_d_bits_sink),
    .auto_in_0_d_bits_denied(tlMasterXbar_auto_in_0_d_bits_denied),
    .auto_in_0_d_bits_data(tlMasterXbar_auto_in_0_d_bits_data),
    .auto_in_0_d_bits_corrupt(tlMasterXbar_auto_in_0_d_bits_corrupt),
    .auto_in_0_e_ready(tlMasterXbar_auto_in_0_e_ready),
    .auto_in_0_e_valid(tlMasterXbar_auto_in_0_e_valid),
    .auto_in_0_e_bits_sink(tlMasterXbar_auto_in_0_e_bits_sink),
    .auto_out_a_ready(tlMasterXbar_auto_out_a_ready),
    .auto_out_a_valid(tlMasterXbar_auto_out_a_valid),
    .auto_out_a_bits_opcode(tlMasterXbar_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(tlMasterXbar_auto_out_a_bits_param),
    .auto_out_a_bits_size(tlMasterXbar_auto_out_a_bits_size),
    .auto_out_a_bits_source(tlMasterXbar_auto_out_a_bits_source),
    .auto_out_a_bits_address(tlMasterXbar_auto_out_a_bits_address),
    .auto_out_a_bits_mask(tlMasterXbar_auto_out_a_bits_mask),
    .auto_out_a_bits_data(tlMasterXbar_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(tlMasterXbar_auto_out_a_bits_corrupt),
    .auto_out_b_ready(tlMasterXbar_auto_out_b_ready),
    .auto_out_b_valid(tlMasterXbar_auto_out_b_valid),
    .auto_out_b_bits_opcode(tlMasterXbar_auto_out_b_bits_opcode),
    .auto_out_b_bits_param(tlMasterXbar_auto_out_b_bits_param),
    .auto_out_b_bits_size(tlMasterXbar_auto_out_b_bits_size),
    .auto_out_b_bits_source(tlMasterXbar_auto_out_b_bits_source),
    .auto_out_b_bits_address(tlMasterXbar_auto_out_b_bits_address),
    .auto_out_b_bits_mask(tlMasterXbar_auto_out_b_bits_mask),
    .auto_out_b_bits_data(tlMasterXbar_auto_out_b_bits_data),
    .auto_out_b_bits_corrupt(tlMasterXbar_auto_out_b_bits_corrupt),
    .auto_out_c_ready(tlMasterXbar_auto_out_c_ready),
    .auto_out_c_valid(tlMasterXbar_auto_out_c_valid),
    .auto_out_c_bits_opcode(tlMasterXbar_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(tlMasterXbar_auto_out_c_bits_param),
    .auto_out_c_bits_size(tlMasterXbar_auto_out_c_bits_size),
    .auto_out_c_bits_source(tlMasterXbar_auto_out_c_bits_source),
    .auto_out_c_bits_address(tlMasterXbar_auto_out_c_bits_address),
    .auto_out_c_bits_data(tlMasterXbar_auto_out_c_bits_data),
    .auto_out_c_bits_corrupt(tlMasterXbar_auto_out_c_bits_corrupt),
    .auto_out_d_ready(tlMasterXbar_auto_out_d_ready),
    .auto_out_d_valid(tlMasterXbar_auto_out_d_valid),
    .auto_out_d_bits_opcode(tlMasterXbar_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(tlMasterXbar_auto_out_d_bits_param),
    .auto_out_d_bits_size(tlMasterXbar_auto_out_d_bits_size),
    .auto_out_d_bits_source(tlMasterXbar_auto_out_d_bits_source),
    .auto_out_d_bits_sink(tlMasterXbar_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(tlMasterXbar_auto_out_d_bits_denied),
    .auto_out_d_bits_data(tlMasterXbar_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(tlMasterXbar_auto_out_d_bits_corrupt),
    .auto_out_e_ready(tlMasterXbar_auto_out_e_ready),
    .auto_out_e_valid(tlMasterXbar_auto_out_e_valid),
    .auto_out_e_bits_sink(tlMasterXbar_auto_out_e_bits_sink)
  );
  TLXbar_8 tlSlaveXbar ( // @[BaseTile.scala 196:41]
    .clock(tlSlaveXbar_clock),
    .reset(tlSlaveXbar_reset)
  );
  IntXbar_1 intXbar ( // @[BaseTile.scala 197:37]
    .clock(intXbar_clock),
    .reset(intXbar_reset),
    .auto_int_in_3_0(intXbar_auto_int_in_3_0),
    .auto_int_in_2_0(intXbar_auto_int_in_2_0),
    .auto_int_in_1_0(intXbar_auto_int_in_1_0),
    .auto_int_in_1_1(intXbar_auto_int_in_1_1),
    .auto_int_in_0_0(intXbar_auto_int_in_0_0),
    .auto_int_out_0(intXbar_auto_int_out_0),
    .auto_int_out_1(intXbar_auto_int_out_1),
    .auto_int_out_2(intXbar_auto_int_out_2),
    .auto_int_out_3(intXbar_auto_int_out_3),
    .auto_int_out_4(intXbar_auto_int_out_4)
  );
  BundleBridgeNexus_6 broadcast ( // @[BundleBridge.scala 196:31]
    .clock(broadcast_clock),
    .reset(broadcast_reset),
    .auto_in(broadcast_auto_in),
    .auto_out(broadcast_auto_out)
  );
  BundleBridgeNexus_7 broadcast_1 ( // @[BundleBridge.scala 196:31]
    .clock(broadcast_1_clock),
    .reset(broadcast_1_reset),
    .auto_in(broadcast_1_auto_in),
    .auto_out_1(broadcast_1_auto_out_1),
    .auto_out_0(broadcast_1_auto_out_0)
  );
  BundleBridgeNexus_8 broadcast_2 ( // @[BundleBridge.scala 196:31]
    .clock(broadcast_2_clock),
    .reset(broadcast_2_reset),
    .auto_in_rnmi(broadcast_2_auto_in_rnmi),
    .auto_in_rnmi_interrupt_vector(broadcast_2_auto_in_rnmi_interrupt_vector),
    .auto_in_rnmi_exception_vector(broadcast_2_auto_in_rnmi_exception_vector),
    .auto_in_unmi(broadcast_2_auto_in_unmi),
    .auto_in_unmi_interrupt_vector(broadcast_2_auto_in_unmi_interrupt_vector),
    .auto_in_unmi_exception_vector(broadcast_2_auto_in_unmi_exception_vector),
    .auto_out_rnmi(broadcast_2_auto_out_rnmi),
    .auto_out_rnmi_interrupt_vector(broadcast_2_auto_out_rnmi_interrupt_vector),
    .auto_out_rnmi_exception_vector(broadcast_2_auto_out_rnmi_exception_vector),
    .auto_out_unmi(broadcast_2_auto_out_unmi),
    .auto_out_unmi_interrupt_vector(broadcast_2_auto_out_unmi_interrupt_vector),
    .auto_out_unmi_exception_vector(broadcast_2_auto_out_unmi_exception_vector)
  );
  BundleBridgeNexus nexus ( // @[BundleBridge.scala 183:27]
    .clock(nexus_clock),
    .reset(nexus_reset)
  );
  BundleBridgeNexus_10 broadcast_3 ( // @[BundleBridge.scala 196:31]
    .clock(broadcast_3_clock),
    .reset(broadcast_3_reset),
    .auto_in_0_valid(broadcast_3_auto_in_0_valid),
    .auto_in_0_iaddr(broadcast_3_auto_in_0_iaddr),
    .auto_in_0_insn(broadcast_3_auto_in_0_insn),
    .auto_in_0_priv(broadcast_3_auto_in_0_priv),
    .auto_in_0_exception(broadcast_3_auto_in_0_exception),
    .auto_in_0_interrupt(broadcast_3_auto_in_0_interrupt),
    .auto_in_0_cause(broadcast_3_auto_in_0_cause),
    .auto_in_0_tval(broadcast_3_auto_in_0_tval),
    .auto_in_1_valid(broadcast_3_auto_in_1_valid),
    .auto_in_1_iaddr(broadcast_3_auto_in_1_iaddr),
    .auto_in_1_insn(broadcast_3_auto_in_1_insn),
    .auto_in_1_priv(broadcast_3_auto_in_1_priv),
    .auto_in_1_exception(broadcast_3_auto_in_1_exception),
    .auto_in_1_interrupt(broadcast_3_auto_in_1_interrupt),
    .auto_in_1_cause(broadcast_3_auto_in_1_cause),
    .auto_in_1_tval(broadcast_3_auto_in_1_tval),
    .auto_out_0_valid(broadcast_3_auto_out_0_valid),
    .auto_out_0_iaddr(broadcast_3_auto_out_0_iaddr),
    .auto_out_0_insn(broadcast_3_auto_out_0_insn),
    .auto_out_0_priv(broadcast_3_auto_out_0_priv),
    .auto_out_0_exception(broadcast_3_auto_out_0_exception),
    .auto_out_0_interrupt(broadcast_3_auto_out_0_interrupt),
    .auto_out_0_cause(broadcast_3_auto_out_0_cause),
    .auto_out_0_tval(broadcast_3_auto_out_0_tval),
    .auto_out_1_valid(broadcast_3_auto_out_1_valid),
    .auto_out_1_iaddr(broadcast_3_auto_out_1_iaddr),
    .auto_out_1_insn(broadcast_3_auto_out_1_insn),
    .auto_out_1_priv(broadcast_3_auto_out_1_priv),
    .auto_out_1_exception(broadcast_3_auto_out_1_exception),
    .auto_out_1_interrupt(broadcast_3_auto_out_1_interrupt),
    .auto_out_1_cause(broadcast_3_auto_out_1_cause),
    .auto_out_1_tval(broadcast_3_auto_out_1_tval)
  );
  BundleBridgeNexus_11 nexus_1 ( // @[BundleBridge.scala 183:27]
    .clock(nexus_1_clock),
    .reset(nexus_1_reset),
    .auto_out_enable(nexus_1_auto_out_enable),
    .auto_out_stall(nexus_1_auto_out_stall)
  );
  BundleBridgeNexus_12 broadcast_4 ( // @[BundleBridge.scala 196:31]
    .clock(broadcast_4_clock),
    .reset(broadcast_4_reset)
  );
  BundleBridgeNexus_13 trace ( // @[BundleBridge.scala 196:31]
    .clock(trace_clock),
    .reset(trace_reset),
    .auto_in_0_valid(trace_auto_in_0_valid),
    .auto_in_0_iaddr(trace_auto_in_0_iaddr),
    .auto_in_0_insn(trace_auto_in_0_insn),
    .auto_in_0_priv(trace_auto_in_0_priv),
    .auto_in_0_exception(trace_auto_in_0_exception),
    .auto_in_0_interrupt(trace_auto_in_0_interrupt),
    .auto_in_0_cause(trace_auto_in_0_cause),
    .auto_in_0_tval(trace_auto_in_0_tval),
    .auto_in_0_wdata(trace_auto_in_0_wdata),
    .auto_in_1_valid(trace_auto_in_1_valid),
    .auto_in_1_iaddr(trace_auto_in_1_iaddr),
    .auto_in_1_insn(trace_auto_in_1_insn),
    .auto_in_1_priv(trace_auto_in_1_priv),
    .auto_in_1_exception(trace_auto_in_1_exception),
    .auto_in_1_interrupt(trace_auto_in_1_interrupt),
    .auto_in_1_cause(trace_auto_in_1_cause),
    .auto_in_1_tval(trace_auto_in_1_tval),
    .auto_in_1_wdata(trace_auto_in_1_wdata),
    .auto_out_0_valid(trace_auto_out_0_valid),
    .auto_out_0_iaddr(trace_auto_out_0_iaddr),
    .auto_out_0_insn(trace_auto_out_0_insn),
    .auto_out_0_priv(trace_auto_out_0_priv),
    .auto_out_0_exception(trace_auto_out_0_exception),
    .auto_out_0_interrupt(trace_auto_out_0_interrupt),
    .auto_out_0_cause(trace_auto_out_0_cause),
    .auto_out_0_tval(trace_auto_out_0_tval),
    .auto_out_0_wdata(trace_auto_out_0_wdata),
    .auto_out_1_valid(trace_auto_out_1_valid),
    .auto_out_1_iaddr(trace_auto_out_1_iaddr),
    .auto_out_1_insn(trace_auto_out_1_insn),
    .auto_out_1_priv(trace_auto_out_1_priv),
    .auto_out_1_exception(trace_auto_out_1_exception),
    .auto_out_1_interrupt(trace_auto_out_1_interrupt),
    .auto_out_1_cause(trace_auto_out_1_cause),
    .auto_out_1_tval(trace_auto_out_1_tval),
    .auto_out_1_wdata(trace_auto_out_1_wdata)
  );
  BoomNonBlockingDCache dcache ( // @[tile.scala 134:54]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .auto_out_a_ready(dcache_auto_out_a_ready),
    .auto_out_a_valid(dcache_auto_out_a_valid),
    .auto_out_a_bits_opcode(dcache_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(dcache_auto_out_a_bits_param),
    .auto_out_a_bits_size(dcache_auto_out_a_bits_size),
    .auto_out_a_bits_source(dcache_auto_out_a_bits_source),
    .auto_out_a_bits_address(dcache_auto_out_a_bits_address),
    .auto_out_a_bits_mask(dcache_auto_out_a_bits_mask),
    .auto_out_a_bits_data(dcache_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(dcache_auto_out_a_bits_corrupt),
    .auto_out_b_ready(dcache_auto_out_b_ready),
    .auto_out_b_valid(dcache_auto_out_b_valid),
    .auto_out_b_bits_opcode(dcache_auto_out_b_bits_opcode),
    .auto_out_b_bits_param(dcache_auto_out_b_bits_param),
    .auto_out_b_bits_size(dcache_auto_out_b_bits_size),
    .auto_out_b_bits_source(dcache_auto_out_b_bits_source),
    .auto_out_b_bits_address(dcache_auto_out_b_bits_address),
    .auto_out_b_bits_mask(dcache_auto_out_b_bits_mask),
    .auto_out_b_bits_data(dcache_auto_out_b_bits_data),
    .auto_out_b_bits_corrupt(dcache_auto_out_b_bits_corrupt),
    .auto_out_c_ready(dcache_auto_out_c_ready),
    .auto_out_c_valid(dcache_auto_out_c_valid),
    .auto_out_c_bits_opcode(dcache_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(dcache_auto_out_c_bits_param),
    .auto_out_c_bits_size(dcache_auto_out_c_bits_size),
    .auto_out_c_bits_source(dcache_auto_out_c_bits_source),
    .auto_out_c_bits_address(dcache_auto_out_c_bits_address),
    .auto_out_c_bits_data(dcache_auto_out_c_bits_data),
    .auto_out_c_bits_corrupt(dcache_auto_out_c_bits_corrupt),
    .auto_out_d_ready(dcache_auto_out_d_ready),
    .auto_out_d_valid(dcache_auto_out_d_valid),
    .auto_out_d_bits_opcode(dcache_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(dcache_auto_out_d_bits_param),
    .auto_out_d_bits_size(dcache_auto_out_d_bits_size),
    .auto_out_d_bits_source(dcache_auto_out_d_bits_source),
    .auto_out_d_bits_sink(dcache_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(dcache_auto_out_d_bits_denied),
    .auto_out_d_bits_data(dcache_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(dcache_auto_out_d_bits_corrupt),
    .auto_out_e_ready(dcache_auto_out_e_ready),
    .auto_out_e_valid(dcache_auto_out_e_valid),
    .auto_out_e_bits_sink(dcache_auto_out_e_bits_sink),
    .io_errors_bus_valid(dcache_io_errors_bus_valid),
    .io_errors_bus_bits(dcache_io_errors_bus_bits),
    .io_lsu_req_ready(dcache_io_lsu_req_ready),
    .io_lsu_req_valid(dcache_io_lsu_req_valid),
    .io_lsu_req_bits_0_valid(dcache_io_lsu_req_bits_0_valid),
    .io_lsu_req_bits_0_bits_uop_switch(dcache_io_lsu_req_bits_0_bits_uop_switch),
    .io_lsu_req_bits_0_bits_uop_switch_off(dcache_io_lsu_req_bits_0_bits_uop_switch_off),
    .io_lsu_req_bits_0_bits_uop_is_unicore(dcache_io_lsu_req_bits_0_bits_uop_is_unicore),
    .io_lsu_req_bits_0_bits_uop_shift(dcache_io_lsu_req_bits_0_bits_uop_shift),
    .io_lsu_req_bits_0_bits_uop_lrs3_rtype(dcache_io_lsu_req_bits_0_bits_uop_lrs3_rtype),
    .io_lsu_req_bits_0_bits_uop_rflag(dcache_io_lsu_req_bits_0_bits_uop_rflag),
    .io_lsu_req_bits_0_bits_uop_wflag(dcache_io_lsu_req_bits_0_bits_uop_wflag),
    .io_lsu_req_bits_0_bits_uop_prflag(dcache_io_lsu_req_bits_0_bits_uop_prflag),
    .io_lsu_req_bits_0_bits_uop_pwflag(dcache_io_lsu_req_bits_0_bits_uop_pwflag),
    .io_lsu_req_bits_0_bits_uop_pflag_busy(dcache_io_lsu_req_bits_0_bits_uop_pflag_busy),
    .io_lsu_req_bits_0_bits_uop_stale_pflag(dcache_io_lsu_req_bits_0_bits_uop_stale_pflag),
    .io_lsu_req_bits_0_bits_uop_op1_sel(dcache_io_lsu_req_bits_0_bits_uop_op1_sel),
    .io_lsu_req_bits_0_bits_uop_op2_sel(dcache_io_lsu_req_bits_0_bits_uop_op2_sel),
    .io_lsu_req_bits_0_bits_uop_split_num(dcache_io_lsu_req_bits_0_bits_uop_split_num),
    .io_lsu_req_bits_0_bits_uop_self_index(dcache_io_lsu_req_bits_0_bits_uop_self_index),
    .io_lsu_req_bits_0_bits_uop_rob_inst_idx(dcache_io_lsu_req_bits_0_bits_uop_rob_inst_idx),
    .io_lsu_req_bits_0_bits_uop_address_num(dcache_io_lsu_req_bits_0_bits_uop_address_num),
    .io_lsu_req_bits_0_bits_uop_uopc(dcache_io_lsu_req_bits_0_bits_uop_uopc),
    .io_lsu_req_bits_0_bits_uop_inst(dcache_io_lsu_req_bits_0_bits_uop_inst),
    .io_lsu_req_bits_0_bits_uop_debug_inst(dcache_io_lsu_req_bits_0_bits_uop_debug_inst),
    .io_lsu_req_bits_0_bits_uop_is_rvc(dcache_io_lsu_req_bits_0_bits_uop_is_rvc),
    .io_lsu_req_bits_0_bits_uop_debug_pc(dcache_io_lsu_req_bits_0_bits_uop_debug_pc),
    .io_lsu_req_bits_0_bits_uop_iq_type(dcache_io_lsu_req_bits_0_bits_uop_iq_type),
    .io_lsu_req_bits_0_bits_uop_fu_code(dcache_io_lsu_req_bits_0_bits_uop_fu_code),
    .io_lsu_req_bits_0_bits_uop_ctrl_br_type(dcache_io_lsu_req_bits_0_bits_uop_ctrl_br_type),
    .io_lsu_req_bits_0_bits_uop_ctrl_op1_sel(dcache_io_lsu_req_bits_0_bits_uop_ctrl_op1_sel),
    .io_lsu_req_bits_0_bits_uop_ctrl_op2_sel(dcache_io_lsu_req_bits_0_bits_uop_ctrl_op2_sel),
    .io_lsu_req_bits_0_bits_uop_ctrl_imm_sel(dcache_io_lsu_req_bits_0_bits_uop_ctrl_imm_sel),
    .io_lsu_req_bits_0_bits_uop_ctrl_op_fcn(dcache_io_lsu_req_bits_0_bits_uop_ctrl_op_fcn),
    .io_lsu_req_bits_0_bits_uop_ctrl_fcn_dw(dcache_io_lsu_req_bits_0_bits_uop_ctrl_fcn_dw),
    .io_lsu_req_bits_0_bits_uop_ctrl_csr_cmd(dcache_io_lsu_req_bits_0_bits_uop_ctrl_csr_cmd),
    .io_lsu_req_bits_0_bits_uop_ctrl_is_load(dcache_io_lsu_req_bits_0_bits_uop_ctrl_is_load),
    .io_lsu_req_bits_0_bits_uop_ctrl_is_sta(dcache_io_lsu_req_bits_0_bits_uop_ctrl_is_sta),
    .io_lsu_req_bits_0_bits_uop_ctrl_is_std(dcache_io_lsu_req_bits_0_bits_uop_ctrl_is_std),
    .io_lsu_req_bits_0_bits_uop_ctrl_op3_sel(dcache_io_lsu_req_bits_0_bits_uop_ctrl_op3_sel),
    .io_lsu_req_bits_0_bits_uop_iw_state(dcache_io_lsu_req_bits_0_bits_uop_iw_state),
    .io_lsu_req_bits_0_bits_uop_iw_p1_poisoned(dcache_io_lsu_req_bits_0_bits_uop_iw_p1_poisoned),
    .io_lsu_req_bits_0_bits_uop_iw_p2_poisoned(dcache_io_lsu_req_bits_0_bits_uop_iw_p2_poisoned),
    .io_lsu_req_bits_0_bits_uop_is_br(dcache_io_lsu_req_bits_0_bits_uop_is_br),
    .io_lsu_req_bits_0_bits_uop_is_jalr(dcache_io_lsu_req_bits_0_bits_uop_is_jalr),
    .io_lsu_req_bits_0_bits_uop_is_jal(dcache_io_lsu_req_bits_0_bits_uop_is_jal),
    .io_lsu_req_bits_0_bits_uop_is_sfb(dcache_io_lsu_req_bits_0_bits_uop_is_sfb),
    .io_lsu_req_bits_0_bits_uop_br_mask(dcache_io_lsu_req_bits_0_bits_uop_br_mask),
    .io_lsu_req_bits_0_bits_uop_br_tag(dcache_io_lsu_req_bits_0_bits_uop_br_tag),
    .io_lsu_req_bits_0_bits_uop_ftq_idx(dcache_io_lsu_req_bits_0_bits_uop_ftq_idx),
    .io_lsu_req_bits_0_bits_uop_edge_inst(dcache_io_lsu_req_bits_0_bits_uop_edge_inst),
    .io_lsu_req_bits_0_bits_uop_pc_lob(dcache_io_lsu_req_bits_0_bits_uop_pc_lob),
    .io_lsu_req_bits_0_bits_uop_taken(dcache_io_lsu_req_bits_0_bits_uop_taken),
    .io_lsu_req_bits_0_bits_uop_imm_packed(dcache_io_lsu_req_bits_0_bits_uop_imm_packed),
    .io_lsu_req_bits_0_bits_uop_csr_addr(dcache_io_lsu_req_bits_0_bits_uop_csr_addr),
    .io_lsu_req_bits_0_bits_uop_rob_idx(dcache_io_lsu_req_bits_0_bits_uop_rob_idx),
    .io_lsu_req_bits_0_bits_uop_ldq_idx(dcache_io_lsu_req_bits_0_bits_uop_ldq_idx),
    .io_lsu_req_bits_0_bits_uop_stq_idx(dcache_io_lsu_req_bits_0_bits_uop_stq_idx),
    .io_lsu_req_bits_0_bits_uop_rxq_idx(dcache_io_lsu_req_bits_0_bits_uop_rxq_idx),
    .io_lsu_req_bits_0_bits_uop_pdst(dcache_io_lsu_req_bits_0_bits_uop_pdst),
    .io_lsu_req_bits_0_bits_uop_prs1(dcache_io_lsu_req_bits_0_bits_uop_prs1),
    .io_lsu_req_bits_0_bits_uop_prs2(dcache_io_lsu_req_bits_0_bits_uop_prs2),
    .io_lsu_req_bits_0_bits_uop_prs3(dcache_io_lsu_req_bits_0_bits_uop_prs3),
    .io_lsu_req_bits_0_bits_uop_ppred(dcache_io_lsu_req_bits_0_bits_uop_ppred),
    .io_lsu_req_bits_0_bits_uop_prs1_busy(dcache_io_lsu_req_bits_0_bits_uop_prs1_busy),
    .io_lsu_req_bits_0_bits_uop_prs2_busy(dcache_io_lsu_req_bits_0_bits_uop_prs2_busy),
    .io_lsu_req_bits_0_bits_uop_prs3_busy(dcache_io_lsu_req_bits_0_bits_uop_prs3_busy),
    .io_lsu_req_bits_0_bits_uop_ppred_busy(dcache_io_lsu_req_bits_0_bits_uop_ppred_busy),
    .io_lsu_req_bits_0_bits_uop_stale_pdst(dcache_io_lsu_req_bits_0_bits_uop_stale_pdst),
    .io_lsu_req_bits_0_bits_uop_exception(dcache_io_lsu_req_bits_0_bits_uop_exception),
    .io_lsu_req_bits_0_bits_uop_exc_cause(dcache_io_lsu_req_bits_0_bits_uop_exc_cause),
    .io_lsu_req_bits_0_bits_uop_bypassable(dcache_io_lsu_req_bits_0_bits_uop_bypassable),
    .io_lsu_req_bits_0_bits_uop_mem_cmd(dcache_io_lsu_req_bits_0_bits_uop_mem_cmd),
    .io_lsu_req_bits_0_bits_uop_mem_size(dcache_io_lsu_req_bits_0_bits_uop_mem_size),
    .io_lsu_req_bits_0_bits_uop_mem_signed(dcache_io_lsu_req_bits_0_bits_uop_mem_signed),
    .io_lsu_req_bits_0_bits_uop_is_fence(dcache_io_lsu_req_bits_0_bits_uop_is_fence),
    .io_lsu_req_bits_0_bits_uop_is_fencei(dcache_io_lsu_req_bits_0_bits_uop_is_fencei),
    .io_lsu_req_bits_0_bits_uop_is_amo(dcache_io_lsu_req_bits_0_bits_uop_is_amo),
    .io_lsu_req_bits_0_bits_uop_uses_ldq(dcache_io_lsu_req_bits_0_bits_uop_uses_ldq),
    .io_lsu_req_bits_0_bits_uop_uses_stq(dcache_io_lsu_req_bits_0_bits_uop_uses_stq),
    .io_lsu_req_bits_0_bits_uop_is_sys_pc2epc(dcache_io_lsu_req_bits_0_bits_uop_is_sys_pc2epc),
    .io_lsu_req_bits_0_bits_uop_is_unique(dcache_io_lsu_req_bits_0_bits_uop_is_unique),
    .io_lsu_req_bits_0_bits_uop_flush_on_commit(dcache_io_lsu_req_bits_0_bits_uop_flush_on_commit),
    .io_lsu_req_bits_0_bits_uop_ldst_is_rs1(dcache_io_lsu_req_bits_0_bits_uop_ldst_is_rs1),
    .io_lsu_req_bits_0_bits_uop_ldst(dcache_io_lsu_req_bits_0_bits_uop_ldst),
    .io_lsu_req_bits_0_bits_uop_lrs1(dcache_io_lsu_req_bits_0_bits_uop_lrs1),
    .io_lsu_req_bits_0_bits_uop_lrs2(dcache_io_lsu_req_bits_0_bits_uop_lrs2),
    .io_lsu_req_bits_0_bits_uop_lrs3(dcache_io_lsu_req_bits_0_bits_uop_lrs3),
    .io_lsu_req_bits_0_bits_uop_ldst_val(dcache_io_lsu_req_bits_0_bits_uop_ldst_val),
    .io_lsu_req_bits_0_bits_uop_dst_rtype(dcache_io_lsu_req_bits_0_bits_uop_dst_rtype),
    .io_lsu_req_bits_0_bits_uop_lrs1_rtype(dcache_io_lsu_req_bits_0_bits_uop_lrs1_rtype),
    .io_lsu_req_bits_0_bits_uop_lrs2_rtype(dcache_io_lsu_req_bits_0_bits_uop_lrs2_rtype),
    .io_lsu_req_bits_0_bits_uop_frs3_en(dcache_io_lsu_req_bits_0_bits_uop_frs3_en),
    .io_lsu_req_bits_0_bits_uop_fp_val(dcache_io_lsu_req_bits_0_bits_uop_fp_val),
    .io_lsu_req_bits_0_bits_uop_fp_single(dcache_io_lsu_req_bits_0_bits_uop_fp_single),
    .io_lsu_req_bits_0_bits_uop_xcpt_pf_if(dcache_io_lsu_req_bits_0_bits_uop_xcpt_pf_if),
    .io_lsu_req_bits_0_bits_uop_xcpt_ae_if(dcache_io_lsu_req_bits_0_bits_uop_xcpt_ae_if),
    .io_lsu_req_bits_0_bits_uop_xcpt_ma_if(dcache_io_lsu_req_bits_0_bits_uop_xcpt_ma_if),
    .io_lsu_req_bits_0_bits_uop_bp_debug_if(dcache_io_lsu_req_bits_0_bits_uop_bp_debug_if),
    .io_lsu_req_bits_0_bits_uop_bp_xcpt_if(dcache_io_lsu_req_bits_0_bits_uop_bp_xcpt_if),
    .io_lsu_req_bits_0_bits_uop_debug_fsrc(dcache_io_lsu_req_bits_0_bits_uop_debug_fsrc),
    .io_lsu_req_bits_0_bits_uop_debug_tsrc(dcache_io_lsu_req_bits_0_bits_uop_debug_tsrc),
    .io_lsu_req_bits_0_bits_addr(dcache_io_lsu_req_bits_0_bits_addr),
    .io_lsu_req_bits_0_bits_data(dcache_io_lsu_req_bits_0_bits_data),
    .io_lsu_req_bits_0_bits_is_hella(dcache_io_lsu_req_bits_0_bits_is_hella),
    .io_lsu_s1_kill_0(dcache_io_lsu_s1_kill_0),
    .io_lsu_resp_0_valid(dcache_io_lsu_resp_0_valid),
    .io_lsu_resp_0_bits_uop_switch(dcache_io_lsu_resp_0_bits_uop_switch),
    .io_lsu_resp_0_bits_uop_switch_off(dcache_io_lsu_resp_0_bits_uop_switch_off),
    .io_lsu_resp_0_bits_uop_is_unicore(dcache_io_lsu_resp_0_bits_uop_is_unicore),
    .io_lsu_resp_0_bits_uop_shift(dcache_io_lsu_resp_0_bits_uop_shift),
    .io_lsu_resp_0_bits_uop_lrs3_rtype(dcache_io_lsu_resp_0_bits_uop_lrs3_rtype),
    .io_lsu_resp_0_bits_uop_rflag(dcache_io_lsu_resp_0_bits_uop_rflag),
    .io_lsu_resp_0_bits_uop_wflag(dcache_io_lsu_resp_0_bits_uop_wflag),
    .io_lsu_resp_0_bits_uop_prflag(dcache_io_lsu_resp_0_bits_uop_prflag),
    .io_lsu_resp_0_bits_uop_pwflag(dcache_io_lsu_resp_0_bits_uop_pwflag),
    .io_lsu_resp_0_bits_uop_pflag_busy(dcache_io_lsu_resp_0_bits_uop_pflag_busy),
    .io_lsu_resp_0_bits_uop_stale_pflag(dcache_io_lsu_resp_0_bits_uop_stale_pflag),
    .io_lsu_resp_0_bits_uop_op1_sel(dcache_io_lsu_resp_0_bits_uop_op1_sel),
    .io_lsu_resp_0_bits_uop_op2_sel(dcache_io_lsu_resp_0_bits_uop_op2_sel),
    .io_lsu_resp_0_bits_uop_split_num(dcache_io_lsu_resp_0_bits_uop_split_num),
    .io_lsu_resp_0_bits_uop_self_index(dcache_io_lsu_resp_0_bits_uop_self_index),
    .io_lsu_resp_0_bits_uop_rob_inst_idx(dcache_io_lsu_resp_0_bits_uop_rob_inst_idx),
    .io_lsu_resp_0_bits_uop_address_num(dcache_io_lsu_resp_0_bits_uop_address_num),
    .io_lsu_resp_0_bits_uop_uopc(dcache_io_lsu_resp_0_bits_uop_uopc),
    .io_lsu_resp_0_bits_uop_inst(dcache_io_lsu_resp_0_bits_uop_inst),
    .io_lsu_resp_0_bits_uop_debug_inst(dcache_io_lsu_resp_0_bits_uop_debug_inst),
    .io_lsu_resp_0_bits_uop_is_rvc(dcache_io_lsu_resp_0_bits_uop_is_rvc),
    .io_lsu_resp_0_bits_uop_debug_pc(dcache_io_lsu_resp_0_bits_uop_debug_pc),
    .io_lsu_resp_0_bits_uop_iq_type(dcache_io_lsu_resp_0_bits_uop_iq_type),
    .io_lsu_resp_0_bits_uop_fu_code(dcache_io_lsu_resp_0_bits_uop_fu_code),
    .io_lsu_resp_0_bits_uop_ctrl_br_type(dcache_io_lsu_resp_0_bits_uop_ctrl_br_type),
    .io_lsu_resp_0_bits_uop_ctrl_op1_sel(dcache_io_lsu_resp_0_bits_uop_ctrl_op1_sel),
    .io_lsu_resp_0_bits_uop_ctrl_op2_sel(dcache_io_lsu_resp_0_bits_uop_ctrl_op2_sel),
    .io_lsu_resp_0_bits_uop_ctrl_imm_sel(dcache_io_lsu_resp_0_bits_uop_ctrl_imm_sel),
    .io_lsu_resp_0_bits_uop_ctrl_op_fcn(dcache_io_lsu_resp_0_bits_uop_ctrl_op_fcn),
    .io_lsu_resp_0_bits_uop_ctrl_fcn_dw(dcache_io_lsu_resp_0_bits_uop_ctrl_fcn_dw),
    .io_lsu_resp_0_bits_uop_ctrl_csr_cmd(dcache_io_lsu_resp_0_bits_uop_ctrl_csr_cmd),
    .io_lsu_resp_0_bits_uop_ctrl_is_load(dcache_io_lsu_resp_0_bits_uop_ctrl_is_load),
    .io_lsu_resp_0_bits_uop_ctrl_is_sta(dcache_io_lsu_resp_0_bits_uop_ctrl_is_sta),
    .io_lsu_resp_0_bits_uop_ctrl_is_std(dcache_io_lsu_resp_0_bits_uop_ctrl_is_std),
    .io_lsu_resp_0_bits_uop_ctrl_op3_sel(dcache_io_lsu_resp_0_bits_uop_ctrl_op3_sel),
    .io_lsu_resp_0_bits_uop_iw_state(dcache_io_lsu_resp_0_bits_uop_iw_state),
    .io_lsu_resp_0_bits_uop_iw_p1_poisoned(dcache_io_lsu_resp_0_bits_uop_iw_p1_poisoned),
    .io_lsu_resp_0_bits_uop_iw_p2_poisoned(dcache_io_lsu_resp_0_bits_uop_iw_p2_poisoned),
    .io_lsu_resp_0_bits_uop_is_br(dcache_io_lsu_resp_0_bits_uop_is_br),
    .io_lsu_resp_0_bits_uop_is_jalr(dcache_io_lsu_resp_0_bits_uop_is_jalr),
    .io_lsu_resp_0_bits_uop_is_jal(dcache_io_lsu_resp_0_bits_uop_is_jal),
    .io_lsu_resp_0_bits_uop_is_sfb(dcache_io_lsu_resp_0_bits_uop_is_sfb),
    .io_lsu_resp_0_bits_uop_br_mask(dcache_io_lsu_resp_0_bits_uop_br_mask),
    .io_lsu_resp_0_bits_uop_br_tag(dcache_io_lsu_resp_0_bits_uop_br_tag),
    .io_lsu_resp_0_bits_uop_ftq_idx(dcache_io_lsu_resp_0_bits_uop_ftq_idx),
    .io_lsu_resp_0_bits_uop_edge_inst(dcache_io_lsu_resp_0_bits_uop_edge_inst),
    .io_lsu_resp_0_bits_uop_pc_lob(dcache_io_lsu_resp_0_bits_uop_pc_lob),
    .io_lsu_resp_0_bits_uop_taken(dcache_io_lsu_resp_0_bits_uop_taken),
    .io_lsu_resp_0_bits_uop_imm_packed(dcache_io_lsu_resp_0_bits_uop_imm_packed),
    .io_lsu_resp_0_bits_uop_csr_addr(dcache_io_lsu_resp_0_bits_uop_csr_addr),
    .io_lsu_resp_0_bits_uop_rob_idx(dcache_io_lsu_resp_0_bits_uop_rob_idx),
    .io_lsu_resp_0_bits_uop_ldq_idx(dcache_io_lsu_resp_0_bits_uop_ldq_idx),
    .io_lsu_resp_0_bits_uop_stq_idx(dcache_io_lsu_resp_0_bits_uop_stq_idx),
    .io_lsu_resp_0_bits_uop_rxq_idx(dcache_io_lsu_resp_0_bits_uop_rxq_idx),
    .io_lsu_resp_0_bits_uop_pdst(dcache_io_lsu_resp_0_bits_uop_pdst),
    .io_lsu_resp_0_bits_uop_prs1(dcache_io_lsu_resp_0_bits_uop_prs1),
    .io_lsu_resp_0_bits_uop_prs2(dcache_io_lsu_resp_0_bits_uop_prs2),
    .io_lsu_resp_0_bits_uop_prs3(dcache_io_lsu_resp_0_bits_uop_prs3),
    .io_lsu_resp_0_bits_uop_ppred(dcache_io_lsu_resp_0_bits_uop_ppred),
    .io_lsu_resp_0_bits_uop_prs1_busy(dcache_io_lsu_resp_0_bits_uop_prs1_busy),
    .io_lsu_resp_0_bits_uop_prs2_busy(dcache_io_lsu_resp_0_bits_uop_prs2_busy),
    .io_lsu_resp_0_bits_uop_prs3_busy(dcache_io_lsu_resp_0_bits_uop_prs3_busy),
    .io_lsu_resp_0_bits_uop_ppred_busy(dcache_io_lsu_resp_0_bits_uop_ppred_busy),
    .io_lsu_resp_0_bits_uop_stale_pdst(dcache_io_lsu_resp_0_bits_uop_stale_pdst),
    .io_lsu_resp_0_bits_uop_exception(dcache_io_lsu_resp_0_bits_uop_exception),
    .io_lsu_resp_0_bits_uop_exc_cause(dcache_io_lsu_resp_0_bits_uop_exc_cause),
    .io_lsu_resp_0_bits_uop_bypassable(dcache_io_lsu_resp_0_bits_uop_bypassable),
    .io_lsu_resp_0_bits_uop_mem_cmd(dcache_io_lsu_resp_0_bits_uop_mem_cmd),
    .io_lsu_resp_0_bits_uop_mem_size(dcache_io_lsu_resp_0_bits_uop_mem_size),
    .io_lsu_resp_0_bits_uop_mem_signed(dcache_io_lsu_resp_0_bits_uop_mem_signed),
    .io_lsu_resp_0_bits_uop_is_fence(dcache_io_lsu_resp_0_bits_uop_is_fence),
    .io_lsu_resp_0_bits_uop_is_fencei(dcache_io_lsu_resp_0_bits_uop_is_fencei),
    .io_lsu_resp_0_bits_uop_is_amo(dcache_io_lsu_resp_0_bits_uop_is_amo),
    .io_lsu_resp_0_bits_uop_uses_ldq(dcache_io_lsu_resp_0_bits_uop_uses_ldq),
    .io_lsu_resp_0_bits_uop_uses_stq(dcache_io_lsu_resp_0_bits_uop_uses_stq),
    .io_lsu_resp_0_bits_uop_is_sys_pc2epc(dcache_io_lsu_resp_0_bits_uop_is_sys_pc2epc),
    .io_lsu_resp_0_bits_uop_is_unique(dcache_io_lsu_resp_0_bits_uop_is_unique),
    .io_lsu_resp_0_bits_uop_flush_on_commit(dcache_io_lsu_resp_0_bits_uop_flush_on_commit),
    .io_lsu_resp_0_bits_uop_ldst_is_rs1(dcache_io_lsu_resp_0_bits_uop_ldst_is_rs1),
    .io_lsu_resp_0_bits_uop_ldst(dcache_io_lsu_resp_0_bits_uop_ldst),
    .io_lsu_resp_0_bits_uop_lrs1(dcache_io_lsu_resp_0_bits_uop_lrs1),
    .io_lsu_resp_0_bits_uop_lrs2(dcache_io_lsu_resp_0_bits_uop_lrs2),
    .io_lsu_resp_0_bits_uop_lrs3(dcache_io_lsu_resp_0_bits_uop_lrs3),
    .io_lsu_resp_0_bits_uop_ldst_val(dcache_io_lsu_resp_0_bits_uop_ldst_val),
    .io_lsu_resp_0_bits_uop_dst_rtype(dcache_io_lsu_resp_0_bits_uop_dst_rtype),
    .io_lsu_resp_0_bits_uop_lrs1_rtype(dcache_io_lsu_resp_0_bits_uop_lrs1_rtype),
    .io_lsu_resp_0_bits_uop_lrs2_rtype(dcache_io_lsu_resp_0_bits_uop_lrs2_rtype),
    .io_lsu_resp_0_bits_uop_frs3_en(dcache_io_lsu_resp_0_bits_uop_frs3_en),
    .io_lsu_resp_0_bits_uop_fp_val(dcache_io_lsu_resp_0_bits_uop_fp_val),
    .io_lsu_resp_0_bits_uop_fp_single(dcache_io_lsu_resp_0_bits_uop_fp_single),
    .io_lsu_resp_0_bits_uop_xcpt_pf_if(dcache_io_lsu_resp_0_bits_uop_xcpt_pf_if),
    .io_lsu_resp_0_bits_uop_xcpt_ae_if(dcache_io_lsu_resp_0_bits_uop_xcpt_ae_if),
    .io_lsu_resp_0_bits_uop_xcpt_ma_if(dcache_io_lsu_resp_0_bits_uop_xcpt_ma_if),
    .io_lsu_resp_0_bits_uop_bp_debug_if(dcache_io_lsu_resp_0_bits_uop_bp_debug_if),
    .io_lsu_resp_0_bits_uop_bp_xcpt_if(dcache_io_lsu_resp_0_bits_uop_bp_xcpt_if),
    .io_lsu_resp_0_bits_uop_debug_fsrc(dcache_io_lsu_resp_0_bits_uop_debug_fsrc),
    .io_lsu_resp_0_bits_uop_debug_tsrc(dcache_io_lsu_resp_0_bits_uop_debug_tsrc),
    .io_lsu_resp_0_bits_data(dcache_io_lsu_resp_0_bits_data),
    .io_lsu_resp_0_bits_is_hella(dcache_io_lsu_resp_0_bits_is_hella),
    .io_lsu_nack_0_valid(dcache_io_lsu_nack_0_valid),
    .io_lsu_nack_0_bits_uop_switch(dcache_io_lsu_nack_0_bits_uop_switch),
    .io_lsu_nack_0_bits_uop_switch_off(dcache_io_lsu_nack_0_bits_uop_switch_off),
    .io_lsu_nack_0_bits_uop_is_unicore(dcache_io_lsu_nack_0_bits_uop_is_unicore),
    .io_lsu_nack_0_bits_uop_shift(dcache_io_lsu_nack_0_bits_uop_shift),
    .io_lsu_nack_0_bits_uop_lrs3_rtype(dcache_io_lsu_nack_0_bits_uop_lrs3_rtype),
    .io_lsu_nack_0_bits_uop_rflag(dcache_io_lsu_nack_0_bits_uop_rflag),
    .io_lsu_nack_0_bits_uop_wflag(dcache_io_lsu_nack_0_bits_uop_wflag),
    .io_lsu_nack_0_bits_uop_prflag(dcache_io_lsu_nack_0_bits_uop_prflag),
    .io_lsu_nack_0_bits_uop_pwflag(dcache_io_lsu_nack_0_bits_uop_pwflag),
    .io_lsu_nack_0_bits_uop_pflag_busy(dcache_io_lsu_nack_0_bits_uop_pflag_busy),
    .io_lsu_nack_0_bits_uop_stale_pflag(dcache_io_lsu_nack_0_bits_uop_stale_pflag),
    .io_lsu_nack_0_bits_uop_op1_sel(dcache_io_lsu_nack_0_bits_uop_op1_sel),
    .io_lsu_nack_0_bits_uop_op2_sel(dcache_io_lsu_nack_0_bits_uop_op2_sel),
    .io_lsu_nack_0_bits_uop_split_num(dcache_io_lsu_nack_0_bits_uop_split_num),
    .io_lsu_nack_0_bits_uop_self_index(dcache_io_lsu_nack_0_bits_uop_self_index),
    .io_lsu_nack_0_bits_uop_rob_inst_idx(dcache_io_lsu_nack_0_bits_uop_rob_inst_idx),
    .io_lsu_nack_0_bits_uop_address_num(dcache_io_lsu_nack_0_bits_uop_address_num),
    .io_lsu_nack_0_bits_uop_uopc(dcache_io_lsu_nack_0_bits_uop_uopc),
    .io_lsu_nack_0_bits_uop_inst(dcache_io_lsu_nack_0_bits_uop_inst),
    .io_lsu_nack_0_bits_uop_debug_inst(dcache_io_lsu_nack_0_bits_uop_debug_inst),
    .io_lsu_nack_0_bits_uop_is_rvc(dcache_io_lsu_nack_0_bits_uop_is_rvc),
    .io_lsu_nack_0_bits_uop_debug_pc(dcache_io_lsu_nack_0_bits_uop_debug_pc),
    .io_lsu_nack_0_bits_uop_iq_type(dcache_io_lsu_nack_0_bits_uop_iq_type),
    .io_lsu_nack_0_bits_uop_fu_code(dcache_io_lsu_nack_0_bits_uop_fu_code),
    .io_lsu_nack_0_bits_uop_ctrl_br_type(dcache_io_lsu_nack_0_bits_uop_ctrl_br_type),
    .io_lsu_nack_0_bits_uop_ctrl_op1_sel(dcache_io_lsu_nack_0_bits_uop_ctrl_op1_sel),
    .io_lsu_nack_0_bits_uop_ctrl_op2_sel(dcache_io_lsu_nack_0_bits_uop_ctrl_op2_sel),
    .io_lsu_nack_0_bits_uop_ctrl_imm_sel(dcache_io_lsu_nack_0_bits_uop_ctrl_imm_sel),
    .io_lsu_nack_0_bits_uop_ctrl_op_fcn(dcache_io_lsu_nack_0_bits_uop_ctrl_op_fcn),
    .io_lsu_nack_0_bits_uop_ctrl_fcn_dw(dcache_io_lsu_nack_0_bits_uop_ctrl_fcn_dw),
    .io_lsu_nack_0_bits_uop_ctrl_csr_cmd(dcache_io_lsu_nack_0_bits_uop_ctrl_csr_cmd),
    .io_lsu_nack_0_bits_uop_ctrl_is_load(dcache_io_lsu_nack_0_bits_uop_ctrl_is_load),
    .io_lsu_nack_0_bits_uop_ctrl_is_sta(dcache_io_lsu_nack_0_bits_uop_ctrl_is_sta),
    .io_lsu_nack_0_bits_uop_ctrl_is_std(dcache_io_lsu_nack_0_bits_uop_ctrl_is_std),
    .io_lsu_nack_0_bits_uop_ctrl_op3_sel(dcache_io_lsu_nack_0_bits_uop_ctrl_op3_sel),
    .io_lsu_nack_0_bits_uop_iw_state(dcache_io_lsu_nack_0_bits_uop_iw_state),
    .io_lsu_nack_0_bits_uop_iw_p1_poisoned(dcache_io_lsu_nack_0_bits_uop_iw_p1_poisoned),
    .io_lsu_nack_0_bits_uop_iw_p2_poisoned(dcache_io_lsu_nack_0_bits_uop_iw_p2_poisoned),
    .io_lsu_nack_0_bits_uop_is_br(dcache_io_lsu_nack_0_bits_uop_is_br),
    .io_lsu_nack_0_bits_uop_is_jalr(dcache_io_lsu_nack_0_bits_uop_is_jalr),
    .io_lsu_nack_0_bits_uop_is_jal(dcache_io_lsu_nack_0_bits_uop_is_jal),
    .io_lsu_nack_0_bits_uop_is_sfb(dcache_io_lsu_nack_0_bits_uop_is_sfb),
    .io_lsu_nack_0_bits_uop_br_mask(dcache_io_lsu_nack_0_bits_uop_br_mask),
    .io_lsu_nack_0_bits_uop_br_tag(dcache_io_lsu_nack_0_bits_uop_br_tag),
    .io_lsu_nack_0_bits_uop_ftq_idx(dcache_io_lsu_nack_0_bits_uop_ftq_idx),
    .io_lsu_nack_0_bits_uop_edge_inst(dcache_io_lsu_nack_0_bits_uop_edge_inst),
    .io_lsu_nack_0_bits_uop_pc_lob(dcache_io_lsu_nack_0_bits_uop_pc_lob),
    .io_lsu_nack_0_bits_uop_taken(dcache_io_lsu_nack_0_bits_uop_taken),
    .io_lsu_nack_0_bits_uop_imm_packed(dcache_io_lsu_nack_0_bits_uop_imm_packed),
    .io_lsu_nack_0_bits_uop_csr_addr(dcache_io_lsu_nack_0_bits_uop_csr_addr),
    .io_lsu_nack_0_bits_uop_rob_idx(dcache_io_lsu_nack_0_bits_uop_rob_idx),
    .io_lsu_nack_0_bits_uop_ldq_idx(dcache_io_lsu_nack_0_bits_uop_ldq_idx),
    .io_lsu_nack_0_bits_uop_stq_idx(dcache_io_lsu_nack_0_bits_uop_stq_idx),
    .io_lsu_nack_0_bits_uop_rxq_idx(dcache_io_lsu_nack_0_bits_uop_rxq_idx),
    .io_lsu_nack_0_bits_uop_pdst(dcache_io_lsu_nack_0_bits_uop_pdst),
    .io_lsu_nack_0_bits_uop_prs1(dcache_io_lsu_nack_0_bits_uop_prs1),
    .io_lsu_nack_0_bits_uop_prs2(dcache_io_lsu_nack_0_bits_uop_prs2),
    .io_lsu_nack_0_bits_uop_prs3(dcache_io_lsu_nack_0_bits_uop_prs3),
    .io_lsu_nack_0_bits_uop_ppred(dcache_io_lsu_nack_0_bits_uop_ppred),
    .io_lsu_nack_0_bits_uop_prs1_busy(dcache_io_lsu_nack_0_bits_uop_prs1_busy),
    .io_lsu_nack_0_bits_uop_prs2_busy(dcache_io_lsu_nack_0_bits_uop_prs2_busy),
    .io_lsu_nack_0_bits_uop_prs3_busy(dcache_io_lsu_nack_0_bits_uop_prs3_busy),
    .io_lsu_nack_0_bits_uop_ppred_busy(dcache_io_lsu_nack_0_bits_uop_ppred_busy),
    .io_lsu_nack_0_bits_uop_stale_pdst(dcache_io_lsu_nack_0_bits_uop_stale_pdst),
    .io_lsu_nack_0_bits_uop_exception(dcache_io_lsu_nack_0_bits_uop_exception),
    .io_lsu_nack_0_bits_uop_exc_cause(dcache_io_lsu_nack_0_bits_uop_exc_cause),
    .io_lsu_nack_0_bits_uop_bypassable(dcache_io_lsu_nack_0_bits_uop_bypassable),
    .io_lsu_nack_0_bits_uop_mem_cmd(dcache_io_lsu_nack_0_bits_uop_mem_cmd),
    .io_lsu_nack_0_bits_uop_mem_size(dcache_io_lsu_nack_0_bits_uop_mem_size),
    .io_lsu_nack_0_bits_uop_mem_signed(dcache_io_lsu_nack_0_bits_uop_mem_signed),
    .io_lsu_nack_0_bits_uop_is_fence(dcache_io_lsu_nack_0_bits_uop_is_fence),
    .io_lsu_nack_0_bits_uop_is_fencei(dcache_io_lsu_nack_0_bits_uop_is_fencei),
    .io_lsu_nack_0_bits_uop_is_amo(dcache_io_lsu_nack_0_bits_uop_is_amo),
    .io_lsu_nack_0_bits_uop_uses_ldq(dcache_io_lsu_nack_0_bits_uop_uses_ldq),
    .io_lsu_nack_0_bits_uop_uses_stq(dcache_io_lsu_nack_0_bits_uop_uses_stq),
    .io_lsu_nack_0_bits_uop_is_sys_pc2epc(dcache_io_lsu_nack_0_bits_uop_is_sys_pc2epc),
    .io_lsu_nack_0_bits_uop_is_unique(dcache_io_lsu_nack_0_bits_uop_is_unique),
    .io_lsu_nack_0_bits_uop_flush_on_commit(dcache_io_lsu_nack_0_bits_uop_flush_on_commit),
    .io_lsu_nack_0_bits_uop_ldst_is_rs1(dcache_io_lsu_nack_0_bits_uop_ldst_is_rs1),
    .io_lsu_nack_0_bits_uop_ldst(dcache_io_lsu_nack_0_bits_uop_ldst),
    .io_lsu_nack_0_bits_uop_lrs1(dcache_io_lsu_nack_0_bits_uop_lrs1),
    .io_lsu_nack_0_bits_uop_lrs2(dcache_io_lsu_nack_0_bits_uop_lrs2),
    .io_lsu_nack_0_bits_uop_lrs3(dcache_io_lsu_nack_0_bits_uop_lrs3),
    .io_lsu_nack_0_bits_uop_ldst_val(dcache_io_lsu_nack_0_bits_uop_ldst_val),
    .io_lsu_nack_0_bits_uop_dst_rtype(dcache_io_lsu_nack_0_bits_uop_dst_rtype),
    .io_lsu_nack_0_bits_uop_lrs1_rtype(dcache_io_lsu_nack_0_bits_uop_lrs1_rtype),
    .io_lsu_nack_0_bits_uop_lrs2_rtype(dcache_io_lsu_nack_0_bits_uop_lrs2_rtype),
    .io_lsu_nack_0_bits_uop_frs3_en(dcache_io_lsu_nack_0_bits_uop_frs3_en),
    .io_lsu_nack_0_bits_uop_fp_val(dcache_io_lsu_nack_0_bits_uop_fp_val),
    .io_lsu_nack_0_bits_uop_fp_single(dcache_io_lsu_nack_0_bits_uop_fp_single),
    .io_lsu_nack_0_bits_uop_xcpt_pf_if(dcache_io_lsu_nack_0_bits_uop_xcpt_pf_if),
    .io_lsu_nack_0_bits_uop_xcpt_ae_if(dcache_io_lsu_nack_0_bits_uop_xcpt_ae_if),
    .io_lsu_nack_0_bits_uop_xcpt_ma_if(dcache_io_lsu_nack_0_bits_uop_xcpt_ma_if),
    .io_lsu_nack_0_bits_uop_bp_debug_if(dcache_io_lsu_nack_0_bits_uop_bp_debug_if),
    .io_lsu_nack_0_bits_uop_bp_xcpt_if(dcache_io_lsu_nack_0_bits_uop_bp_xcpt_if),
    .io_lsu_nack_0_bits_uop_debug_fsrc(dcache_io_lsu_nack_0_bits_uop_debug_fsrc),
    .io_lsu_nack_0_bits_uop_debug_tsrc(dcache_io_lsu_nack_0_bits_uop_debug_tsrc),
    .io_lsu_nack_0_bits_addr(dcache_io_lsu_nack_0_bits_addr),
    .io_lsu_nack_0_bits_data(dcache_io_lsu_nack_0_bits_data),
    .io_lsu_nack_0_bits_is_hella(dcache_io_lsu_nack_0_bits_is_hella),
    .io_lsu_brupdate_b1_resolve_mask(dcache_io_lsu_brupdate_b1_resolve_mask),
    .io_lsu_brupdate_b1_mispredict_mask(dcache_io_lsu_brupdate_b1_mispredict_mask),
    .io_lsu_brupdate_b2_uop_switch(dcache_io_lsu_brupdate_b2_uop_switch),
    .io_lsu_brupdate_b2_uop_switch_off(dcache_io_lsu_brupdate_b2_uop_switch_off),
    .io_lsu_brupdate_b2_uop_is_unicore(dcache_io_lsu_brupdate_b2_uop_is_unicore),
    .io_lsu_brupdate_b2_uop_shift(dcache_io_lsu_brupdate_b2_uop_shift),
    .io_lsu_brupdate_b2_uop_lrs3_rtype(dcache_io_lsu_brupdate_b2_uop_lrs3_rtype),
    .io_lsu_brupdate_b2_uop_rflag(dcache_io_lsu_brupdate_b2_uop_rflag),
    .io_lsu_brupdate_b2_uop_wflag(dcache_io_lsu_brupdate_b2_uop_wflag),
    .io_lsu_brupdate_b2_uop_prflag(dcache_io_lsu_brupdate_b2_uop_prflag),
    .io_lsu_brupdate_b2_uop_pwflag(dcache_io_lsu_brupdate_b2_uop_pwflag),
    .io_lsu_brupdate_b2_uop_pflag_busy(dcache_io_lsu_brupdate_b2_uop_pflag_busy),
    .io_lsu_brupdate_b2_uop_stale_pflag(dcache_io_lsu_brupdate_b2_uop_stale_pflag),
    .io_lsu_brupdate_b2_uop_op1_sel(dcache_io_lsu_brupdate_b2_uop_op1_sel),
    .io_lsu_brupdate_b2_uop_op2_sel(dcache_io_lsu_brupdate_b2_uop_op2_sel),
    .io_lsu_brupdate_b2_uop_split_num(dcache_io_lsu_brupdate_b2_uop_split_num),
    .io_lsu_brupdate_b2_uop_self_index(dcache_io_lsu_brupdate_b2_uop_self_index),
    .io_lsu_brupdate_b2_uop_rob_inst_idx(dcache_io_lsu_brupdate_b2_uop_rob_inst_idx),
    .io_lsu_brupdate_b2_uop_address_num(dcache_io_lsu_brupdate_b2_uop_address_num),
    .io_lsu_brupdate_b2_uop_uopc(dcache_io_lsu_brupdate_b2_uop_uopc),
    .io_lsu_brupdate_b2_uop_inst(dcache_io_lsu_brupdate_b2_uop_inst),
    .io_lsu_brupdate_b2_uop_debug_inst(dcache_io_lsu_brupdate_b2_uop_debug_inst),
    .io_lsu_brupdate_b2_uop_is_rvc(dcache_io_lsu_brupdate_b2_uop_is_rvc),
    .io_lsu_brupdate_b2_uop_debug_pc(dcache_io_lsu_brupdate_b2_uop_debug_pc),
    .io_lsu_brupdate_b2_uop_iq_type(dcache_io_lsu_brupdate_b2_uop_iq_type),
    .io_lsu_brupdate_b2_uop_fu_code(dcache_io_lsu_brupdate_b2_uop_fu_code),
    .io_lsu_brupdate_b2_uop_ctrl_br_type(dcache_io_lsu_brupdate_b2_uop_ctrl_br_type),
    .io_lsu_brupdate_b2_uop_ctrl_op1_sel(dcache_io_lsu_brupdate_b2_uop_ctrl_op1_sel),
    .io_lsu_brupdate_b2_uop_ctrl_op2_sel(dcache_io_lsu_brupdate_b2_uop_ctrl_op2_sel),
    .io_lsu_brupdate_b2_uop_ctrl_imm_sel(dcache_io_lsu_brupdate_b2_uop_ctrl_imm_sel),
    .io_lsu_brupdate_b2_uop_ctrl_op_fcn(dcache_io_lsu_brupdate_b2_uop_ctrl_op_fcn),
    .io_lsu_brupdate_b2_uop_ctrl_fcn_dw(dcache_io_lsu_brupdate_b2_uop_ctrl_fcn_dw),
    .io_lsu_brupdate_b2_uop_ctrl_csr_cmd(dcache_io_lsu_brupdate_b2_uop_ctrl_csr_cmd),
    .io_lsu_brupdate_b2_uop_ctrl_is_load(dcache_io_lsu_brupdate_b2_uop_ctrl_is_load),
    .io_lsu_brupdate_b2_uop_ctrl_is_sta(dcache_io_lsu_brupdate_b2_uop_ctrl_is_sta),
    .io_lsu_brupdate_b2_uop_ctrl_is_std(dcache_io_lsu_brupdate_b2_uop_ctrl_is_std),
    .io_lsu_brupdate_b2_uop_ctrl_op3_sel(dcache_io_lsu_brupdate_b2_uop_ctrl_op3_sel),
    .io_lsu_brupdate_b2_uop_iw_state(dcache_io_lsu_brupdate_b2_uop_iw_state),
    .io_lsu_brupdate_b2_uop_iw_p1_poisoned(dcache_io_lsu_brupdate_b2_uop_iw_p1_poisoned),
    .io_lsu_brupdate_b2_uop_iw_p2_poisoned(dcache_io_lsu_brupdate_b2_uop_iw_p2_poisoned),
    .io_lsu_brupdate_b2_uop_is_br(dcache_io_lsu_brupdate_b2_uop_is_br),
    .io_lsu_brupdate_b2_uop_is_jalr(dcache_io_lsu_brupdate_b2_uop_is_jalr),
    .io_lsu_brupdate_b2_uop_is_jal(dcache_io_lsu_brupdate_b2_uop_is_jal),
    .io_lsu_brupdate_b2_uop_is_sfb(dcache_io_lsu_brupdate_b2_uop_is_sfb),
    .io_lsu_brupdate_b2_uop_br_mask(dcache_io_lsu_brupdate_b2_uop_br_mask),
    .io_lsu_brupdate_b2_uop_br_tag(dcache_io_lsu_brupdate_b2_uop_br_tag),
    .io_lsu_brupdate_b2_uop_ftq_idx(dcache_io_lsu_brupdate_b2_uop_ftq_idx),
    .io_lsu_brupdate_b2_uop_edge_inst(dcache_io_lsu_brupdate_b2_uop_edge_inst),
    .io_lsu_brupdate_b2_uop_pc_lob(dcache_io_lsu_brupdate_b2_uop_pc_lob),
    .io_lsu_brupdate_b2_uop_taken(dcache_io_lsu_brupdate_b2_uop_taken),
    .io_lsu_brupdate_b2_uop_imm_packed(dcache_io_lsu_brupdate_b2_uop_imm_packed),
    .io_lsu_brupdate_b2_uop_csr_addr(dcache_io_lsu_brupdate_b2_uop_csr_addr),
    .io_lsu_brupdate_b2_uop_rob_idx(dcache_io_lsu_brupdate_b2_uop_rob_idx),
    .io_lsu_brupdate_b2_uop_ldq_idx(dcache_io_lsu_brupdate_b2_uop_ldq_idx),
    .io_lsu_brupdate_b2_uop_stq_idx(dcache_io_lsu_brupdate_b2_uop_stq_idx),
    .io_lsu_brupdate_b2_uop_rxq_idx(dcache_io_lsu_brupdate_b2_uop_rxq_idx),
    .io_lsu_brupdate_b2_uop_pdst(dcache_io_lsu_brupdate_b2_uop_pdst),
    .io_lsu_brupdate_b2_uop_prs1(dcache_io_lsu_brupdate_b2_uop_prs1),
    .io_lsu_brupdate_b2_uop_prs2(dcache_io_lsu_brupdate_b2_uop_prs2),
    .io_lsu_brupdate_b2_uop_prs3(dcache_io_lsu_brupdate_b2_uop_prs3),
    .io_lsu_brupdate_b2_uop_ppred(dcache_io_lsu_brupdate_b2_uop_ppred),
    .io_lsu_brupdate_b2_uop_prs1_busy(dcache_io_lsu_brupdate_b2_uop_prs1_busy),
    .io_lsu_brupdate_b2_uop_prs2_busy(dcache_io_lsu_brupdate_b2_uop_prs2_busy),
    .io_lsu_brupdate_b2_uop_prs3_busy(dcache_io_lsu_brupdate_b2_uop_prs3_busy),
    .io_lsu_brupdate_b2_uop_ppred_busy(dcache_io_lsu_brupdate_b2_uop_ppred_busy),
    .io_lsu_brupdate_b2_uop_stale_pdst(dcache_io_lsu_brupdate_b2_uop_stale_pdst),
    .io_lsu_brupdate_b2_uop_exception(dcache_io_lsu_brupdate_b2_uop_exception),
    .io_lsu_brupdate_b2_uop_exc_cause(dcache_io_lsu_brupdate_b2_uop_exc_cause),
    .io_lsu_brupdate_b2_uop_bypassable(dcache_io_lsu_brupdate_b2_uop_bypassable),
    .io_lsu_brupdate_b2_uop_mem_cmd(dcache_io_lsu_brupdate_b2_uop_mem_cmd),
    .io_lsu_brupdate_b2_uop_mem_size(dcache_io_lsu_brupdate_b2_uop_mem_size),
    .io_lsu_brupdate_b2_uop_mem_signed(dcache_io_lsu_brupdate_b2_uop_mem_signed),
    .io_lsu_brupdate_b2_uop_is_fence(dcache_io_lsu_brupdate_b2_uop_is_fence),
    .io_lsu_brupdate_b2_uop_is_fencei(dcache_io_lsu_brupdate_b2_uop_is_fencei),
    .io_lsu_brupdate_b2_uop_is_amo(dcache_io_lsu_brupdate_b2_uop_is_amo),
    .io_lsu_brupdate_b2_uop_uses_ldq(dcache_io_lsu_brupdate_b2_uop_uses_ldq),
    .io_lsu_brupdate_b2_uop_uses_stq(dcache_io_lsu_brupdate_b2_uop_uses_stq),
    .io_lsu_brupdate_b2_uop_is_sys_pc2epc(dcache_io_lsu_brupdate_b2_uop_is_sys_pc2epc),
    .io_lsu_brupdate_b2_uop_is_unique(dcache_io_lsu_brupdate_b2_uop_is_unique),
    .io_lsu_brupdate_b2_uop_flush_on_commit(dcache_io_lsu_brupdate_b2_uop_flush_on_commit),
    .io_lsu_brupdate_b2_uop_ldst_is_rs1(dcache_io_lsu_brupdate_b2_uop_ldst_is_rs1),
    .io_lsu_brupdate_b2_uop_ldst(dcache_io_lsu_brupdate_b2_uop_ldst),
    .io_lsu_brupdate_b2_uop_lrs1(dcache_io_lsu_brupdate_b2_uop_lrs1),
    .io_lsu_brupdate_b2_uop_lrs2(dcache_io_lsu_brupdate_b2_uop_lrs2),
    .io_lsu_brupdate_b2_uop_lrs3(dcache_io_lsu_brupdate_b2_uop_lrs3),
    .io_lsu_brupdate_b2_uop_ldst_val(dcache_io_lsu_brupdate_b2_uop_ldst_val),
    .io_lsu_brupdate_b2_uop_dst_rtype(dcache_io_lsu_brupdate_b2_uop_dst_rtype),
    .io_lsu_brupdate_b2_uop_lrs1_rtype(dcache_io_lsu_brupdate_b2_uop_lrs1_rtype),
    .io_lsu_brupdate_b2_uop_lrs2_rtype(dcache_io_lsu_brupdate_b2_uop_lrs2_rtype),
    .io_lsu_brupdate_b2_uop_frs3_en(dcache_io_lsu_brupdate_b2_uop_frs3_en),
    .io_lsu_brupdate_b2_uop_fp_val(dcache_io_lsu_brupdate_b2_uop_fp_val),
    .io_lsu_brupdate_b2_uop_fp_single(dcache_io_lsu_brupdate_b2_uop_fp_single),
    .io_lsu_brupdate_b2_uop_xcpt_pf_if(dcache_io_lsu_brupdate_b2_uop_xcpt_pf_if),
    .io_lsu_brupdate_b2_uop_xcpt_ae_if(dcache_io_lsu_brupdate_b2_uop_xcpt_ae_if),
    .io_lsu_brupdate_b2_uop_xcpt_ma_if(dcache_io_lsu_brupdate_b2_uop_xcpt_ma_if),
    .io_lsu_brupdate_b2_uop_bp_debug_if(dcache_io_lsu_brupdate_b2_uop_bp_debug_if),
    .io_lsu_brupdate_b2_uop_bp_xcpt_if(dcache_io_lsu_brupdate_b2_uop_bp_xcpt_if),
    .io_lsu_brupdate_b2_uop_debug_fsrc(dcache_io_lsu_brupdate_b2_uop_debug_fsrc),
    .io_lsu_brupdate_b2_uop_debug_tsrc(dcache_io_lsu_brupdate_b2_uop_debug_tsrc),
    .io_lsu_brupdate_b2_valid(dcache_io_lsu_brupdate_b2_valid),
    .io_lsu_brupdate_b2_mispredict(dcache_io_lsu_brupdate_b2_mispredict),
    .io_lsu_brupdate_b2_taken(dcache_io_lsu_brupdate_b2_taken),
    .io_lsu_brupdate_b2_cfi_type(dcache_io_lsu_brupdate_b2_cfi_type),
    .io_lsu_brupdate_b2_pc_sel(dcache_io_lsu_brupdate_b2_pc_sel),
    .io_lsu_brupdate_b2_jalr_target(dcache_io_lsu_brupdate_b2_jalr_target),
    .io_lsu_brupdate_b2_target_offset(dcache_io_lsu_brupdate_b2_target_offset),
    .io_lsu_exception(dcache_io_lsu_exception),
    .io_lsu_rob_pnr_idx(dcache_io_lsu_rob_pnr_idx),
    .io_lsu_rob_head_idx(dcache_io_lsu_rob_head_idx),
    .io_lsu_release_ready(dcache_io_lsu_release_ready),
    .io_lsu_release_valid(dcache_io_lsu_release_valid),
    .io_lsu_release_bits_opcode(dcache_io_lsu_release_bits_opcode),
    .io_lsu_release_bits_param(dcache_io_lsu_release_bits_param),
    .io_lsu_release_bits_size(dcache_io_lsu_release_bits_size),
    .io_lsu_release_bits_source(dcache_io_lsu_release_bits_source),
    .io_lsu_release_bits_address(dcache_io_lsu_release_bits_address),
    .io_lsu_release_bits_data(dcache_io_lsu_release_bits_data),
    .io_lsu_release_bits_corrupt(dcache_io_lsu_release_bits_corrupt),
    .io_lsu_force_order(dcache_io_lsu_force_order),
    .io_lsu_ordered(dcache_io_lsu_ordered),
    .io_lsu_perf_acquire(dcache_io_lsu_perf_acquire),
    .io_lsu_perf_release(dcache_io_lsu_perf_release)
  );
  BoomFrontend frontend ( // @[tile.scala 140:28]
    .clock(frontend_clock),
    .reset(frontend_reset),
    .auto_icache_master_out_a_ready(frontend_auto_icache_master_out_a_ready),
    .auto_icache_master_out_a_valid(frontend_auto_icache_master_out_a_valid),
    .auto_icache_master_out_a_bits_opcode(frontend_auto_icache_master_out_a_bits_opcode),
    .auto_icache_master_out_a_bits_param(frontend_auto_icache_master_out_a_bits_param),
    .auto_icache_master_out_a_bits_size(frontend_auto_icache_master_out_a_bits_size),
    .auto_icache_master_out_a_bits_source(frontend_auto_icache_master_out_a_bits_source),
    .auto_icache_master_out_a_bits_address(frontend_auto_icache_master_out_a_bits_address),
    .auto_icache_master_out_a_bits_mask(frontend_auto_icache_master_out_a_bits_mask),
    .auto_icache_master_out_a_bits_data(frontend_auto_icache_master_out_a_bits_data),
    .auto_icache_master_out_a_bits_corrupt(frontend_auto_icache_master_out_a_bits_corrupt),
    .auto_icache_master_out_d_ready(frontend_auto_icache_master_out_d_ready),
    .auto_icache_master_out_d_valid(frontend_auto_icache_master_out_d_valid),
    .auto_icache_master_out_d_bits_opcode(frontend_auto_icache_master_out_d_bits_opcode),
    .auto_icache_master_out_d_bits_param(frontend_auto_icache_master_out_d_bits_param),
    .auto_icache_master_out_d_bits_size(frontend_auto_icache_master_out_d_bits_size),
    .auto_icache_master_out_d_bits_source(frontend_auto_icache_master_out_d_bits_source),
    .auto_icache_master_out_d_bits_sink(frontend_auto_icache_master_out_d_bits_sink),
    .auto_icache_master_out_d_bits_denied(frontend_auto_icache_master_out_d_bits_denied),
    .auto_icache_master_out_d_bits_data(frontend_auto_icache_master_out_d_bits_data),
    .auto_icache_master_out_d_bits_corrupt(frontend_auto_icache_master_out_d_bits_corrupt),
    .auto_reset_vector_sink_in(frontend_auto_reset_vector_sink_in),
    .io_cpu_fetchpacket_ready(frontend_io_cpu_fetchpacket_ready),
    .io_cpu_fetchpacket_valid(frontend_io_cpu_fetchpacket_valid),
    .io_cpu_fetchpacket_bits_uops_0_valid(frontend_io_cpu_fetchpacket_bits_uops_0_valid),
    .io_cpu_fetchpacket_bits_uops_0_bits_switch(frontend_io_cpu_fetchpacket_bits_uops_0_bits_switch),
    .io_cpu_fetchpacket_bits_uops_0_bits_switch_off(frontend_io_cpu_fetchpacket_bits_uops_0_bits_switch_off),
    .io_cpu_fetchpacket_bits_uops_0_bits_is_unicore(frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_unicore),
    .io_cpu_fetchpacket_bits_uops_0_bits_shift(frontend_io_cpu_fetchpacket_bits_uops_0_bits_shift),
    .io_cpu_fetchpacket_bits_uops_0_bits_lrs3_rtype(frontend_io_cpu_fetchpacket_bits_uops_0_bits_lrs3_rtype),
    .io_cpu_fetchpacket_bits_uops_0_bits_rflag(frontend_io_cpu_fetchpacket_bits_uops_0_bits_rflag),
    .io_cpu_fetchpacket_bits_uops_0_bits_wflag(frontend_io_cpu_fetchpacket_bits_uops_0_bits_wflag),
    .io_cpu_fetchpacket_bits_uops_0_bits_prflag(frontend_io_cpu_fetchpacket_bits_uops_0_bits_prflag),
    .io_cpu_fetchpacket_bits_uops_0_bits_pwflag(frontend_io_cpu_fetchpacket_bits_uops_0_bits_pwflag),
    .io_cpu_fetchpacket_bits_uops_0_bits_pflag_busy(frontend_io_cpu_fetchpacket_bits_uops_0_bits_pflag_busy),
    .io_cpu_fetchpacket_bits_uops_0_bits_stale_pflag(frontend_io_cpu_fetchpacket_bits_uops_0_bits_stale_pflag),
    .io_cpu_fetchpacket_bits_uops_0_bits_op1_sel(frontend_io_cpu_fetchpacket_bits_uops_0_bits_op1_sel),
    .io_cpu_fetchpacket_bits_uops_0_bits_op2_sel(frontend_io_cpu_fetchpacket_bits_uops_0_bits_op2_sel),
    .io_cpu_fetchpacket_bits_uops_0_bits_split_num(frontend_io_cpu_fetchpacket_bits_uops_0_bits_split_num),
    .io_cpu_fetchpacket_bits_uops_0_bits_self_index(frontend_io_cpu_fetchpacket_bits_uops_0_bits_self_index),
    .io_cpu_fetchpacket_bits_uops_0_bits_rob_inst_idx(frontend_io_cpu_fetchpacket_bits_uops_0_bits_rob_inst_idx),
    .io_cpu_fetchpacket_bits_uops_0_bits_address_num(frontend_io_cpu_fetchpacket_bits_uops_0_bits_address_num),
    .io_cpu_fetchpacket_bits_uops_0_bits_uopc(frontend_io_cpu_fetchpacket_bits_uops_0_bits_uopc),
    .io_cpu_fetchpacket_bits_uops_0_bits_inst(frontend_io_cpu_fetchpacket_bits_uops_0_bits_inst),
    .io_cpu_fetchpacket_bits_uops_0_bits_debug_inst(frontend_io_cpu_fetchpacket_bits_uops_0_bits_debug_inst),
    .io_cpu_fetchpacket_bits_uops_0_bits_is_rvc(frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_rvc),
    .io_cpu_fetchpacket_bits_uops_0_bits_debug_pc(frontend_io_cpu_fetchpacket_bits_uops_0_bits_debug_pc),
    .io_cpu_fetchpacket_bits_uops_0_bits_iq_type(frontend_io_cpu_fetchpacket_bits_uops_0_bits_iq_type),
    .io_cpu_fetchpacket_bits_uops_0_bits_fu_code(frontend_io_cpu_fetchpacket_bits_uops_0_bits_fu_code),
    .io_cpu_fetchpacket_bits_uops_0_bits_ctrl_br_type(frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_br_type),
    .io_cpu_fetchpacket_bits_uops_0_bits_ctrl_op1_sel(frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_op1_sel),
    .io_cpu_fetchpacket_bits_uops_0_bits_ctrl_op2_sel(frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_op2_sel),
    .io_cpu_fetchpacket_bits_uops_0_bits_ctrl_imm_sel(frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_imm_sel),
    .io_cpu_fetchpacket_bits_uops_0_bits_ctrl_op_fcn(frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_op_fcn),
    .io_cpu_fetchpacket_bits_uops_0_bits_ctrl_fcn_dw(frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_fcn_dw),
    .io_cpu_fetchpacket_bits_uops_0_bits_ctrl_csr_cmd(frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_csr_cmd),
    .io_cpu_fetchpacket_bits_uops_0_bits_ctrl_is_load(frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_is_load),
    .io_cpu_fetchpacket_bits_uops_0_bits_ctrl_is_sta(frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_is_sta),
    .io_cpu_fetchpacket_bits_uops_0_bits_ctrl_is_std(frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_is_std),
    .io_cpu_fetchpacket_bits_uops_0_bits_ctrl_op3_sel(frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_op3_sel),
    .io_cpu_fetchpacket_bits_uops_0_bits_iw_state(frontend_io_cpu_fetchpacket_bits_uops_0_bits_iw_state),
    .io_cpu_fetchpacket_bits_uops_0_bits_iw_p1_poisoned(frontend_io_cpu_fetchpacket_bits_uops_0_bits_iw_p1_poisoned),
    .io_cpu_fetchpacket_bits_uops_0_bits_iw_p2_poisoned(frontend_io_cpu_fetchpacket_bits_uops_0_bits_iw_p2_poisoned),
    .io_cpu_fetchpacket_bits_uops_0_bits_is_br(frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_br),
    .io_cpu_fetchpacket_bits_uops_0_bits_is_jalr(frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_jalr),
    .io_cpu_fetchpacket_bits_uops_0_bits_is_jal(frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_jal),
    .io_cpu_fetchpacket_bits_uops_0_bits_is_sfb(frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_sfb),
    .io_cpu_fetchpacket_bits_uops_0_bits_br_mask(frontend_io_cpu_fetchpacket_bits_uops_0_bits_br_mask),
    .io_cpu_fetchpacket_bits_uops_0_bits_br_tag(frontend_io_cpu_fetchpacket_bits_uops_0_bits_br_tag),
    .io_cpu_fetchpacket_bits_uops_0_bits_ftq_idx(frontend_io_cpu_fetchpacket_bits_uops_0_bits_ftq_idx),
    .io_cpu_fetchpacket_bits_uops_0_bits_edge_inst(frontend_io_cpu_fetchpacket_bits_uops_0_bits_edge_inst),
    .io_cpu_fetchpacket_bits_uops_0_bits_pc_lob(frontend_io_cpu_fetchpacket_bits_uops_0_bits_pc_lob),
    .io_cpu_fetchpacket_bits_uops_0_bits_taken(frontend_io_cpu_fetchpacket_bits_uops_0_bits_taken),
    .io_cpu_fetchpacket_bits_uops_0_bits_imm_packed(frontend_io_cpu_fetchpacket_bits_uops_0_bits_imm_packed),
    .io_cpu_fetchpacket_bits_uops_0_bits_csr_addr(frontend_io_cpu_fetchpacket_bits_uops_0_bits_csr_addr),
    .io_cpu_fetchpacket_bits_uops_0_bits_rob_idx(frontend_io_cpu_fetchpacket_bits_uops_0_bits_rob_idx),
    .io_cpu_fetchpacket_bits_uops_0_bits_ldq_idx(frontend_io_cpu_fetchpacket_bits_uops_0_bits_ldq_idx),
    .io_cpu_fetchpacket_bits_uops_0_bits_stq_idx(frontend_io_cpu_fetchpacket_bits_uops_0_bits_stq_idx),
    .io_cpu_fetchpacket_bits_uops_0_bits_rxq_idx(frontend_io_cpu_fetchpacket_bits_uops_0_bits_rxq_idx),
    .io_cpu_fetchpacket_bits_uops_0_bits_pdst(frontend_io_cpu_fetchpacket_bits_uops_0_bits_pdst),
    .io_cpu_fetchpacket_bits_uops_0_bits_prs1(frontend_io_cpu_fetchpacket_bits_uops_0_bits_prs1),
    .io_cpu_fetchpacket_bits_uops_0_bits_prs2(frontend_io_cpu_fetchpacket_bits_uops_0_bits_prs2),
    .io_cpu_fetchpacket_bits_uops_0_bits_prs3(frontend_io_cpu_fetchpacket_bits_uops_0_bits_prs3),
    .io_cpu_fetchpacket_bits_uops_0_bits_ppred(frontend_io_cpu_fetchpacket_bits_uops_0_bits_ppred),
    .io_cpu_fetchpacket_bits_uops_0_bits_prs1_busy(frontend_io_cpu_fetchpacket_bits_uops_0_bits_prs1_busy),
    .io_cpu_fetchpacket_bits_uops_0_bits_prs2_busy(frontend_io_cpu_fetchpacket_bits_uops_0_bits_prs2_busy),
    .io_cpu_fetchpacket_bits_uops_0_bits_prs3_busy(frontend_io_cpu_fetchpacket_bits_uops_0_bits_prs3_busy),
    .io_cpu_fetchpacket_bits_uops_0_bits_ppred_busy(frontend_io_cpu_fetchpacket_bits_uops_0_bits_ppred_busy),
    .io_cpu_fetchpacket_bits_uops_0_bits_stale_pdst(frontend_io_cpu_fetchpacket_bits_uops_0_bits_stale_pdst),
    .io_cpu_fetchpacket_bits_uops_0_bits_exception(frontend_io_cpu_fetchpacket_bits_uops_0_bits_exception),
    .io_cpu_fetchpacket_bits_uops_0_bits_exc_cause(frontend_io_cpu_fetchpacket_bits_uops_0_bits_exc_cause),
    .io_cpu_fetchpacket_bits_uops_0_bits_bypassable(frontend_io_cpu_fetchpacket_bits_uops_0_bits_bypassable),
    .io_cpu_fetchpacket_bits_uops_0_bits_mem_cmd(frontend_io_cpu_fetchpacket_bits_uops_0_bits_mem_cmd),
    .io_cpu_fetchpacket_bits_uops_0_bits_mem_size(frontend_io_cpu_fetchpacket_bits_uops_0_bits_mem_size),
    .io_cpu_fetchpacket_bits_uops_0_bits_mem_signed(frontend_io_cpu_fetchpacket_bits_uops_0_bits_mem_signed),
    .io_cpu_fetchpacket_bits_uops_0_bits_is_fence(frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_fence),
    .io_cpu_fetchpacket_bits_uops_0_bits_is_fencei(frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_fencei),
    .io_cpu_fetchpacket_bits_uops_0_bits_is_amo(frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_amo),
    .io_cpu_fetchpacket_bits_uops_0_bits_uses_ldq(frontend_io_cpu_fetchpacket_bits_uops_0_bits_uses_ldq),
    .io_cpu_fetchpacket_bits_uops_0_bits_uses_stq(frontend_io_cpu_fetchpacket_bits_uops_0_bits_uses_stq),
    .io_cpu_fetchpacket_bits_uops_0_bits_is_sys_pc2epc(frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_sys_pc2epc),
    .io_cpu_fetchpacket_bits_uops_0_bits_is_unique(frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_unique),
    .io_cpu_fetchpacket_bits_uops_0_bits_flush_on_commit(frontend_io_cpu_fetchpacket_bits_uops_0_bits_flush_on_commit),
    .io_cpu_fetchpacket_bits_uops_0_bits_ldst_is_rs1(frontend_io_cpu_fetchpacket_bits_uops_0_bits_ldst_is_rs1),
    .io_cpu_fetchpacket_bits_uops_0_bits_ldst(frontend_io_cpu_fetchpacket_bits_uops_0_bits_ldst),
    .io_cpu_fetchpacket_bits_uops_0_bits_lrs1(frontend_io_cpu_fetchpacket_bits_uops_0_bits_lrs1),
    .io_cpu_fetchpacket_bits_uops_0_bits_lrs2(frontend_io_cpu_fetchpacket_bits_uops_0_bits_lrs2),
    .io_cpu_fetchpacket_bits_uops_0_bits_lrs3(frontend_io_cpu_fetchpacket_bits_uops_0_bits_lrs3),
    .io_cpu_fetchpacket_bits_uops_0_bits_ldst_val(frontend_io_cpu_fetchpacket_bits_uops_0_bits_ldst_val),
    .io_cpu_fetchpacket_bits_uops_0_bits_dst_rtype(frontend_io_cpu_fetchpacket_bits_uops_0_bits_dst_rtype),
    .io_cpu_fetchpacket_bits_uops_0_bits_lrs1_rtype(frontend_io_cpu_fetchpacket_bits_uops_0_bits_lrs1_rtype),
    .io_cpu_fetchpacket_bits_uops_0_bits_lrs2_rtype(frontend_io_cpu_fetchpacket_bits_uops_0_bits_lrs2_rtype),
    .io_cpu_fetchpacket_bits_uops_0_bits_frs3_en(frontend_io_cpu_fetchpacket_bits_uops_0_bits_frs3_en),
    .io_cpu_fetchpacket_bits_uops_0_bits_fp_val(frontend_io_cpu_fetchpacket_bits_uops_0_bits_fp_val),
    .io_cpu_fetchpacket_bits_uops_0_bits_fp_single(frontend_io_cpu_fetchpacket_bits_uops_0_bits_fp_single),
    .io_cpu_fetchpacket_bits_uops_0_bits_xcpt_pf_if(frontend_io_cpu_fetchpacket_bits_uops_0_bits_xcpt_pf_if),
    .io_cpu_fetchpacket_bits_uops_0_bits_xcpt_ae_if(frontend_io_cpu_fetchpacket_bits_uops_0_bits_xcpt_ae_if),
    .io_cpu_fetchpacket_bits_uops_0_bits_xcpt_ma_if(frontend_io_cpu_fetchpacket_bits_uops_0_bits_xcpt_ma_if),
    .io_cpu_fetchpacket_bits_uops_0_bits_bp_debug_if(frontend_io_cpu_fetchpacket_bits_uops_0_bits_bp_debug_if),
    .io_cpu_fetchpacket_bits_uops_0_bits_bp_xcpt_if(frontend_io_cpu_fetchpacket_bits_uops_0_bits_bp_xcpt_if),
    .io_cpu_fetchpacket_bits_uops_0_bits_debug_fsrc(frontend_io_cpu_fetchpacket_bits_uops_0_bits_debug_fsrc),
    .io_cpu_fetchpacket_bits_uops_0_bits_debug_tsrc(frontend_io_cpu_fetchpacket_bits_uops_0_bits_debug_tsrc),
    .io_cpu_fetchpacket_bits_uops_1_valid(frontend_io_cpu_fetchpacket_bits_uops_1_valid),
    .io_cpu_fetchpacket_bits_uops_1_bits_switch(frontend_io_cpu_fetchpacket_bits_uops_1_bits_switch),
    .io_cpu_fetchpacket_bits_uops_1_bits_switch_off(frontend_io_cpu_fetchpacket_bits_uops_1_bits_switch_off),
    .io_cpu_fetchpacket_bits_uops_1_bits_is_unicore(frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_unicore),
    .io_cpu_fetchpacket_bits_uops_1_bits_shift(frontend_io_cpu_fetchpacket_bits_uops_1_bits_shift),
    .io_cpu_fetchpacket_bits_uops_1_bits_lrs3_rtype(frontend_io_cpu_fetchpacket_bits_uops_1_bits_lrs3_rtype),
    .io_cpu_fetchpacket_bits_uops_1_bits_rflag(frontend_io_cpu_fetchpacket_bits_uops_1_bits_rflag),
    .io_cpu_fetchpacket_bits_uops_1_bits_wflag(frontend_io_cpu_fetchpacket_bits_uops_1_bits_wflag),
    .io_cpu_fetchpacket_bits_uops_1_bits_prflag(frontend_io_cpu_fetchpacket_bits_uops_1_bits_prflag),
    .io_cpu_fetchpacket_bits_uops_1_bits_pwflag(frontend_io_cpu_fetchpacket_bits_uops_1_bits_pwflag),
    .io_cpu_fetchpacket_bits_uops_1_bits_pflag_busy(frontend_io_cpu_fetchpacket_bits_uops_1_bits_pflag_busy),
    .io_cpu_fetchpacket_bits_uops_1_bits_stale_pflag(frontend_io_cpu_fetchpacket_bits_uops_1_bits_stale_pflag),
    .io_cpu_fetchpacket_bits_uops_1_bits_op1_sel(frontend_io_cpu_fetchpacket_bits_uops_1_bits_op1_sel),
    .io_cpu_fetchpacket_bits_uops_1_bits_op2_sel(frontend_io_cpu_fetchpacket_bits_uops_1_bits_op2_sel),
    .io_cpu_fetchpacket_bits_uops_1_bits_split_num(frontend_io_cpu_fetchpacket_bits_uops_1_bits_split_num),
    .io_cpu_fetchpacket_bits_uops_1_bits_self_index(frontend_io_cpu_fetchpacket_bits_uops_1_bits_self_index),
    .io_cpu_fetchpacket_bits_uops_1_bits_rob_inst_idx(frontend_io_cpu_fetchpacket_bits_uops_1_bits_rob_inst_idx),
    .io_cpu_fetchpacket_bits_uops_1_bits_address_num(frontend_io_cpu_fetchpacket_bits_uops_1_bits_address_num),
    .io_cpu_fetchpacket_bits_uops_1_bits_uopc(frontend_io_cpu_fetchpacket_bits_uops_1_bits_uopc),
    .io_cpu_fetchpacket_bits_uops_1_bits_inst(frontend_io_cpu_fetchpacket_bits_uops_1_bits_inst),
    .io_cpu_fetchpacket_bits_uops_1_bits_debug_inst(frontend_io_cpu_fetchpacket_bits_uops_1_bits_debug_inst),
    .io_cpu_fetchpacket_bits_uops_1_bits_is_rvc(frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_rvc),
    .io_cpu_fetchpacket_bits_uops_1_bits_debug_pc(frontend_io_cpu_fetchpacket_bits_uops_1_bits_debug_pc),
    .io_cpu_fetchpacket_bits_uops_1_bits_iq_type(frontend_io_cpu_fetchpacket_bits_uops_1_bits_iq_type),
    .io_cpu_fetchpacket_bits_uops_1_bits_fu_code(frontend_io_cpu_fetchpacket_bits_uops_1_bits_fu_code),
    .io_cpu_fetchpacket_bits_uops_1_bits_ctrl_br_type(frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_br_type),
    .io_cpu_fetchpacket_bits_uops_1_bits_ctrl_op1_sel(frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_op1_sel),
    .io_cpu_fetchpacket_bits_uops_1_bits_ctrl_op2_sel(frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_op2_sel),
    .io_cpu_fetchpacket_bits_uops_1_bits_ctrl_imm_sel(frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_imm_sel),
    .io_cpu_fetchpacket_bits_uops_1_bits_ctrl_op_fcn(frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_op_fcn),
    .io_cpu_fetchpacket_bits_uops_1_bits_ctrl_fcn_dw(frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_fcn_dw),
    .io_cpu_fetchpacket_bits_uops_1_bits_ctrl_csr_cmd(frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_csr_cmd),
    .io_cpu_fetchpacket_bits_uops_1_bits_ctrl_is_load(frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_is_load),
    .io_cpu_fetchpacket_bits_uops_1_bits_ctrl_is_sta(frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_is_sta),
    .io_cpu_fetchpacket_bits_uops_1_bits_ctrl_is_std(frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_is_std),
    .io_cpu_fetchpacket_bits_uops_1_bits_ctrl_op3_sel(frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_op3_sel),
    .io_cpu_fetchpacket_bits_uops_1_bits_iw_state(frontend_io_cpu_fetchpacket_bits_uops_1_bits_iw_state),
    .io_cpu_fetchpacket_bits_uops_1_bits_iw_p1_poisoned(frontend_io_cpu_fetchpacket_bits_uops_1_bits_iw_p1_poisoned),
    .io_cpu_fetchpacket_bits_uops_1_bits_iw_p2_poisoned(frontend_io_cpu_fetchpacket_bits_uops_1_bits_iw_p2_poisoned),
    .io_cpu_fetchpacket_bits_uops_1_bits_is_br(frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_br),
    .io_cpu_fetchpacket_bits_uops_1_bits_is_jalr(frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_jalr),
    .io_cpu_fetchpacket_bits_uops_1_bits_is_jal(frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_jal),
    .io_cpu_fetchpacket_bits_uops_1_bits_is_sfb(frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_sfb),
    .io_cpu_fetchpacket_bits_uops_1_bits_br_mask(frontend_io_cpu_fetchpacket_bits_uops_1_bits_br_mask),
    .io_cpu_fetchpacket_bits_uops_1_bits_br_tag(frontend_io_cpu_fetchpacket_bits_uops_1_bits_br_tag),
    .io_cpu_fetchpacket_bits_uops_1_bits_ftq_idx(frontend_io_cpu_fetchpacket_bits_uops_1_bits_ftq_idx),
    .io_cpu_fetchpacket_bits_uops_1_bits_edge_inst(frontend_io_cpu_fetchpacket_bits_uops_1_bits_edge_inst),
    .io_cpu_fetchpacket_bits_uops_1_bits_pc_lob(frontend_io_cpu_fetchpacket_bits_uops_1_bits_pc_lob),
    .io_cpu_fetchpacket_bits_uops_1_bits_taken(frontend_io_cpu_fetchpacket_bits_uops_1_bits_taken),
    .io_cpu_fetchpacket_bits_uops_1_bits_imm_packed(frontend_io_cpu_fetchpacket_bits_uops_1_bits_imm_packed),
    .io_cpu_fetchpacket_bits_uops_1_bits_csr_addr(frontend_io_cpu_fetchpacket_bits_uops_1_bits_csr_addr),
    .io_cpu_fetchpacket_bits_uops_1_bits_rob_idx(frontend_io_cpu_fetchpacket_bits_uops_1_bits_rob_idx),
    .io_cpu_fetchpacket_bits_uops_1_bits_ldq_idx(frontend_io_cpu_fetchpacket_bits_uops_1_bits_ldq_idx),
    .io_cpu_fetchpacket_bits_uops_1_bits_stq_idx(frontend_io_cpu_fetchpacket_bits_uops_1_bits_stq_idx),
    .io_cpu_fetchpacket_bits_uops_1_bits_rxq_idx(frontend_io_cpu_fetchpacket_bits_uops_1_bits_rxq_idx),
    .io_cpu_fetchpacket_bits_uops_1_bits_pdst(frontend_io_cpu_fetchpacket_bits_uops_1_bits_pdst),
    .io_cpu_fetchpacket_bits_uops_1_bits_prs1(frontend_io_cpu_fetchpacket_bits_uops_1_bits_prs1),
    .io_cpu_fetchpacket_bits_uops_1_bits_prs2(frontend_io_cpu_fetchpacket_bits_uops_1_bits_prs2),
    .io_cpu_fetchpacket_bits_uops_1_bits_prs3(frontend_io_cpu_fetchpacket_bits_uops_1_bits_prs3),
    .io_cpu_fetchpacket_bits_uops_1_bits_ppred(frontend_io_cpu_fetchpacket_bits_uops_1_bits_ppred),
    .io_cpu_fetchpacket_bits_uops_1_bits_prs1_busy(frontend_io_cpu_fetchpacket_bits_uops_1_bits_prs1_busy),
    .io_cpu_fetchpacket_bits_uops_1_bits_prs2_busy(frontend_io_cpu_fetchpacket_bits_uops_1_bits_prs2_busy),
    .io_cpu_fetchpacket_bits_uops_1_bits_prs3_busy(frontend_io_cpu_fetchpacket_bits_uops_1_bits_prs3_busy),
    .io_cpu_fetchpacket_bits_uops_1_bits_ppred_busy(frontend_io_cpu_fetchpacket_bits_uops_1_bits_ppred_busy),
    .io_cpu_fetchpacket_bits_uops_1_bits_stale_pdst(frontend_io_cpu_fetchpacket_bits_uops_1_bits_stale_pdst),
    .io_cpu_fetchpacket_bits_uops_1_bits_exception(frontend_io_cpu_fetchpacket_bits_uops_1_bits_exception),
    .io_cpu_fetchpacket_bits_uops_1_bits_exc_cause(frontend_io_cpu_fetchpacket_bits_uops_1_bits_exc_cause),
    .io_cpu_fetchpacket_bits_uops_1_bits_bypassable(frontend_io_cpu_fetchpacket_bits_uops_1_bits_bypassable),
    .io_cpu_fetchpacket_bits_uops_1_bits_mem_cmd(frontend_io_cpu_fetchpacket_bits_uops_1_bits_mem_cmd),
    .io_cpu_fetchpacket_bits_uops_1_bits_mem_size(frontend_io_cpu_fetchpacket_bits_uops_1_bits_mem_size),
    .io_cpu_fetchpacket_bits_uops_1_bits_mem_signed(frontend_io_cpu_fetchpacket_bits_uops_1_bits_mem_signed),
    .io_cpu_fetchpacket_bits_uops_1_bits_is_fence(frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_fence),
    .io_cpu_fetchpacket_bits_uops_1_bits_is_fencei(frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_fencei),
    .io_cpu_fetchpacket_bits_uops_1_bits_is_amo(frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_amo),
    .io_cpu_fetchpacket_bits_uops_1_bits_uses_ldq(frontend_io_cpu_fetchpacket_bits_uops_1_bits_uses_ldq),
    .io_cpu_fetchpacket_bits_uops_1_bits_uses_stq(frontend_io_cpu_fetchpacket_bits_uops_1_bits_uses_stq),
    .io_cpu_fetchpacket_bits_uops_1_bits_is_sys_pc2epc(frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_sys_pc2epc),
    .io_cpu_fetchpacket_bits_uops_1_bits_is_unique(frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_unique),
    .io_cpu_fetchpacket_bits_uops_1_bits_flush_on_commit(frontend_io_cpu_fetchpacket_bits_uops_1_bits_flush_on_commit),
    .io_cpu_fetchpacket_bits_uops_1_bits_ldst_is_rs1(frontend_io_cpu_fetchpacket_bits_uops_1_bits_ldst_is_rs1),
    .io_cpu_fetchpacket_bits_uops_1_bits_ldst(frontend_io_cpu_fetchpacket_bits_uops_1_bits_ldst),
    .io_cpu_fetchpacket_bits_uops_1_bits_lrs1(frontend_io_cpu_fetchpacket_bits_uops_1_bits_lrs1),
    .io_cpu_fetchpacket_bits_uops_1_bits_lrs2(frontend_io_cpu_fetchpacket_bits_uops_1_bits_lrs2),
    .io_cpu_fetchpacket_bits_uops_1_bits_lrs3(frontend_io_cpu_fetchpacket_bits_uops_1_bits_lrs3),
    .io_cpu_fetchpacket_bits_uops_1_bits_ldst_val(frontend_io_cpu_fetchpacket_bits_uops_1_bits_ldst_val),
    .io_cpu_fetchpacket_bits_uops_1_bits_dst_rtype(frontend_io_cpu_fetchpacket_bits_uops_1_bits_dst_rtype),
    .io_cpu_fetchpacket_bits_uops_1_bits_lrs1_rtype(frontend_io_cpu_fetchpacket_bits_uops_1_bits_lrs1_rtype),
    .io_cpu_fetchpacket_bits_uops_1_bits_lrs2_rtype(frontend_io_cpu_fetchpacket_bits_uops_1_bits_lrs2_rtype),
    .io_cpu_fetchpacket_bits_uops_1_bits_frs3_en(frontend_io_cpu_fetchpacket_bits_uops_1_bits_frs3_en),
    .io_cpu_fetchpacket_bits_uops_1_bits_fp_val(frontend_io_cpu_fetchpacket_bits_uops_1_bits_fp_val),
    .io_cpu_fetchpacket_bits_uops_1_bits_fp_single(frontend_io_cpu_fetchpacket_bits_uops_1_bits_fp_single),
    .io_cpu_fetchpacket_bits_uops_1_bits_xcpt_pf_if(frontend_io_cpu_fetchpacket_bits_uops_1_bits_xcpt_pf_if),
    .io_cpu_fetchpacket_bits_uops_1_bits_xcpt_ae_if(frontend_io_cpu_fetchpacket_bits_uops_1_bits_xcpt_ae_if),
    .io_cpu_fetchpacket_bits_uops_1_bits_xcpt_ma_if(frontend_io_cpu_fetchpacket_bits_uops_1_bits_xcpt_ma_if),
    .io_cpu_fetchpacket_bits_uops_1_bits_bp_debug_if(frontend_io_cpu_fetchpacket_bits_uops_1_bits_bp_debug_if),
    .io_cpu_fetchpacket_bits_uops_1_bits_bp_xcpt_if(frontend_io_cpu_fetchpacket_bits_uops_1_bits_bp_xcpt_if),
    .io_cpu_fetchpacket_bits_uops_1_bits_debug_fsrc(frontend_io_cpu_fetchpacket_bits_uops_1_bits_debug_fsrc),
    .io_cpu_fetchpacket_bits_uops_1_bits_debug_tsrc(frontend_io_cpu_fetchpacket_bits_uops_1_bits_debug_tsrc),
    .io_cpu_get_pc_0_ftq_idx(frontend_io_cpu_get_pc_0_ftq_idx),
    .io_cpu_get_pc_0_entry_cfi_idx_valid(frontend_io_cpu_get_pc_0_entry_cfi_idx_valid),
    .io_cpu_get_pc_0_entry_cfi_idx_bits(frontend_io_cpu_get_pc_0_entry_cfi_idx_bits),
    .io_cpu_get_pc_0_entry_cfi_taken(frontend_io_cpu_get_pc_0_entry_cfi_taken),
    .io_cpu_get_pc_0_entry_cfi_mispredicted(frontend_io_cpu_get_pc_0_entry_cfi_mispredicted),
    .io_cpu_get_pc_0_entry_cfi_type(frontend_io_cpu_get_pc_0_entry_cfi_type),
    .io_cpu_get_pc_0_entry_br_mask(frontend_io_cpu_get_pc_0_entry_br_mask),
    .io_cpu_get_pc_0_entry_cfi_is_call(frontend_io_cpu_get_pc_0_entry_cfi_is_call),
    .io_cpu_get_pc_0_entry_cfi_is_ret(frontend_io_cpu_get_pc_0_entry_cfi_is_ret),
    .io_cpu_get_pc_0_entry_cfi_npc_plus4(frontend_io_cpu_get_pc_0_entry_cfi_npc_plus4),
    .io_cpu_get_pc_0_entry_ras_top(frontend_io_cpu_get_pc_0_entry_ras_top),
    .io_cpu_get_pc_0_entry_ras_idx(frontend_io_cpu_get_pc_0_entry_ras_idx),
    .io_cpu_get_pc_0_entry_start_bank(frontend_io_cpu_get_pc_0_entry_start_bank),
    .io_cpu_get_pc_0_ghist_old_history(frontend_io_cpu_get_pc_0_ghist_old_history),
    .io_cpu_get_pc_0_ghist_current_saw_branch_not_taken(frontend_io_cpu_get_pc_0_ghist_current_saw_branch_not_taken),
    .io_cpu_get_pc_0_ghist_new_saw_branch_not_taken(frontend_io_cpu_get_pc_0_ghist_new_saw_branch_not_taken),
    .io_cpu_get_pc_0_ghist_new_saw_branch_taken(frontend_io_cpu_get_pc_0_ghist_new_saw_branch_taken),
    .io_cpu_get_pc_0_ghist_ras_idx(frontend_io_cpu_get_pc_0_ghist_ras_idx),
    .io_cpu_get_pc_0_pc(frontend_io_cpu_get_pc_0_pc),
    .io_cpu_get_pc_0_com_pc(frontend_io_cpu_get_pc_0_com_pc),
    .io_cpu_get_pc_0_next_val(frontend_io_cpu_get_pc_0_next_val),
    .io_cpu_get_pc_0_next_pc(frontend_io_cpu_get_pc_0_next_pc),
    .io_cpu_get_pc_1_ftq_idx(frontend_io_cpu_get_pc_1_ftq_idx),
    .io_cpu_get_pc_1_entry_cfi_idx_valid(frontend_io_cpu_get_pc_1_entry_cfi_idx_valid),
    .io_cpu_get_pc_1_entry_cfi_idx_bits(frontend_io_cpu_get_pc_1_entry_cfi_idx_bits),
    .io_cpu_get_pc_1_entry_cfi_taken(frontend_io_cpu_get_pc_1_entry_cfi_taken),
    .io_cpu_get_pc_1_entry_cfi_mispredicted(frontend_io_cpu_get_pc_1_entry_cfi_mispredicted),
    .io_cpu_get_pc_1_entry_cfi_type(frontend_io_cpu_get_pc_1_entry_cfi_type),
    .io_cpu_get_pc_1_entry_br_mask(frontend_io_cpu_get_pc_1_entry_br_mask),
    .io_cpu_get_pc_1_entry_cfi_is_call(frontend_io_cpu_get_pc_1_entry_cfi_is_call),
    .io_cpu_get_pc_1_entry_cfi_is_ret(frontend_io_cpu_get_pc_1_entry_cfi_is_ret),
    .io_cpu_get_pc_1_entry_cfi_npc_plus4(frontend_io_cpu_get_pc_1_entry_cfi_npc_plus4),
    .io_cpu_get_pc_1_entry_ras_top(frontend_io_cpu_get_pc_1_entry_ras_top),
    .io_cpu_get_pc_1_entry_ras_idx(frontend_io_cpu_get_pc_1_entry_ras_idx),
    .io_cpu_get_pc_1_entry_start_bank(frontend_io_cpu_get_pc_1_entry_start_bank),
    .io_cpu_get_pc_1_ghist_old_history(frontend_io_cpu_get_pc_1_ghist_old_history),
    .io_cpu_get_pc_1_ghist_current_saw_branch_not_taken(frontend_io_cpu_get_pc_1_ghist_current_saw_branch_not_taken),
    .io_cpu_get_pc_1_ghist_new_saw_branch_not_taken(frontend_io_cpu_get_pc_1_ghist_new_saw_branch_not_taken),
    .io_cpu_get_pc_1_ghist_new_saw_branch_taken(frontend_io_cpu_get_pc_1_ghist_new_saw_branch_taken),
    .io_cpu_get_pc_1_ghist_ras_idx(frontend_io_cpu_get_pc_1_ghist_ras_idx),
    .io_cpu_get_pc_1_pc(frontend_io_cpu_get_pc_1_pc),
    .io_cpu_get_pc_1_com_pc(frontend_io_cpu_get_pc_1_com_pc),
    .io_cpu_get_pc_1_next_val(frontend_io_cpu_get_pc_1_next_val),
    .io_cpu_get_pc_1_next_pc(frontend_io_cpu_get_pc_1_next_pc),
    .io_cpu_get_pc_2_ftq_idx(frontend_io_cpu_get_pc_2_ftq_idx),
    .io_cpu_get_pc_2_entry_cfi_idx_valid(frontend_io_cpu_get_pc_2_entry_cfi_idx_valid),
    .io_cpu_get_pc_2_entry_cfi_idx_bits(frontend_io_cpu_get_pc_2_entry_cfi_idx_bits),
    .io_cpu_get_pc_2_entry_cfi_taken(frontend_io_cpu_get_pc_2_entry_cfi_taken),
    .io_cpu_get_pc_2_entry_cfi_mispredicted(frontend_io_cpu_get_pc_2_entry_cfi_mispredicted),
    .io_cpu_get_pc_2_entry_cfi_type(frontend_io_cpu_get_pc_2_entry_cfi_type),
    .io_cpu_get_pc_2_entry_br_mask(frontend_io_cpu_get_pc_2_entry_br_mask),
    .io_cpu_get_pc_2_entry_cfi_is_call(frontend_io_cpu_get_pc_2_entry_cfi_is_call),
    .io_cpu_get_pc_2_entry_cfi_is_ret(frontend_io_cpu_get_pc_2_entry_cfi_is_ret),
    .io_cpu_get_pc_2_entry_cfi_npc_plus4(frontend_io_cpu_get_pc_2_entry_cfi_npc_plus4),
    .io_cpu_get_pc_2_entry_ras_top(frontend_io_cpu_get_pc_2_entry_ras_top),
    .io_cpu_get_pc_2_entry_ras_idx(frontend_io_cpu_get_pc_2_entry_ras_idx),
    .io_cpu_get_pc_2_entry_start_bank(frontend_io_cpu_get_pc_2_entry_start_bank),
    .io_cpu_get_pc_2_ghist_old_history(frontend_io_cpu_get_pc_2_ghist_old_history),
    .io_cpu_get_pc_2_ghist_current_saw_branch_not_taken(frontend_io_cpu_get_pc_2_ghist_current_saw_branch_not_taken),
    .io_cpu_get_pc_2_ghist_new_saw_branch_not_taken(frontend_io_cpu_get_pc_2_ghist_new_saw_branch_not_taken),
    .io_cpu_get_pc_2_ghist_new_saw_branch_taken(frontend_io_cpu_get_pc_2_ghist_new_saw_branch_taken),
    .io_cpu_get_pc_2_ghist_ras_idx(frontend_io_cpu_get_pc_2_ghist_ras_idx),
    .io_cpu_get_pc_2_pc(frontend_io_cpu_get_pc_2_pc),
    .io_cpu_get_pc_2_com_pc(frontend_io_cpu_get_pc_2_com_pc),
    .io_cpu_get_pc_2_next_val(frontend_io_cpu_get_pc_2_next_val),
    .io_cpu_get_pc_2_next_pc(frontend_io_cpu_get_pc_2_next_pc),
    .io_cpu_get_pc_3_ftq_idx(frontend_io_cpu_get_pc_3_ftq_idx),
    .io_cpu_get_pc_3_entry_cfi_idx_valid(frontend_io_cpu_get_pc_3_entry_cfi_idx_valid),
    .io_cpu_get_pc_3_entry_cfi_idx_bits(frontend_io_cpu_get_pc_3_entry_cfi_idx_bits),
    .io_cpu_get_pc_3_entry_cfi_taken(frontend_io_cpu_get_pc_3_entry_cfi_taken),
    .io_cpu_get_pc_3_entry_cfi_mispredicted(frontend_io_cpu_get_pc_3_entry_cfi_mispredicted),
    .io_cpu_get_pc_3_entry_cfi_type(frontend_io_cpu_get_pc_3_entry_cfi_type),
    .io_cpu_get_pc_3_entry_br_mask(frontend_io_cpu_get_pc_3_entry_br_mask),
    .io_cpu_get_pc_3_entry_cfi_is_call(frontend_io_cpu_get_pc_3_entry_cfi_is_call),
    .io_cpu_get_pc_3_entry_cfi_is_ret(frontend_io_cpu_get_pc_3_entry_cfi_is_ret),
    .io_cpu_get_pc_3_entry_cfi_npc_plus4(frontend_io_cpu_get_pc_3_entry_cfi_npc_plus4),
    .io_cpu_get_pc_3_entry_ras_top(frontend_io_cpu_get_pc_3_entry_ras_top),
    .io_cpu_get_pc_3_entry_ras_idx(frontend_io_cpu_get_pc_3_entry_ras_idx),
    .io_cpu_get_pc_3_entry_start_bank(frontend_io_cpu_get_pc_3_entry_start_bank),
    .io_cpu_get_pc_3_ghist_old_history(frontend_io_cpu_get_pc_3_ghist_old_history),
    .io_cpu_get_pc_3_ghist_current_saw_branch_not_taken(frontend_io_cpu_get_pc_3_ghist_current_saw_branch_not_taken),
    .io_cpu_get_pc_3_ghist_new_saw_branch_not_taken(frontend_io_cpu_get_pc_3_ghist_new_saw_branch_not_taken),
    .io_cpu_get_pc_3_ghist_new_saw_branch_taken(frontend_io_cpu_get_pc_3_ghist_new_saw_branch_taken),
    .io_cpu_get_pc_3_ghist_ras_idx(frontend_io_cpu_get_pc_3_ghist_ras_idx),
    .io_cpu_get_pc_3_pc(frontend_io_cpu_get_pc_3_pc),
    .io_cpu_get_pc_3_com_pc(frontend_io_cpu_get_pc_3_com_pc),
    .io_cpu_get_pc_3_next_val(frontend_io_cpu_get_pc_3_next_val),
    .io_cpu_get_pc_3_next_pc(frontend_io_cpu_get_pc_3_next_pc),
    .io_cpu_debug_ftq_idx_0(frontend_io_cpu_debug_ftq_idx_0),
    .io_cpu_debug_ftq_idx_1(frontend_io_cpu_debug_ftq_idx_1),
    .io_cpu_debug_fetch_pc_0(frontend_io_cpu_debug_fetch_pc_0),
    .io_cpu_debug_fetch_pc_1(frontend_io_cpu_debug_fetch_pc_1),
    .io_cpu_status_debug(frontend_io_cpu_status_debug),
    .io_cpu_status_cease(frontend_io_cpu_status_cease),
    .io_cpu_status_wfi(frontend_io_cpu_status_wfi),
    .io_cpu_status_isa(frontend_io_cpu_status_isa),
    .io_cpu_status_dprv(frontend_io_cpu_status_dprv),
    .io_cpu_status_prv(frontend_io_cpu_status_prv),
    .io_cpu_status_sd(frontend_io_cpu_status_sd),
    .io_cpu_status_zero2(frontend_io_cpu_status_zero2),
    .io_cpu_status_sxl(frontend_io_cpu_status_sxl),
    .io_cpu_status_uxl(frontend_io_cpu_status_uxl),
    .io_cpu_status_sd_rv32(frontend_io_cpu_status_sd_rv32),
    .io_cpu_status_zero1(frontend_io_cpu_status_zero1),
    .io_cpu_status_tsr(frontend_io_cpu_status_tsr),
    .io_cpu_status_tw(frontend_io_cpu_status_tw),
    .io_cpu_status_tvm(frontend_io_cpu_status_tvm),
    .io_cpu_status_mxr(frontend_io_cpu_status_mxr),
    .io_cpu_status_sum(frontend_io_cpu_status_sum),
    .io_cpu_status_mprv(frontend_io_cpu_status_mprv),
    .io_cpu_status_xs(frontend_io_cpu_status_xs),
    .io_cpu_status_fs(frontend_io_cpu_status_fs),
    .io_cpu_status_mpp(frontend_io_cpu_status_mpp),
    .io_cpu_status_vs(frontend_io_cpu_status_vs),
    .io_cpu_status_spp(frontend_io_cpu_status_spp),
    .io_cpu_status_mpie(frontend_io_cpu_status_mpie),
    .io_cpu_status_hpie(frontend_io_cpu_status_hpie),
    .io_cpu_status_spie(frontend_io_cpu_status_spie),
    .io_cpu_status_upie(frontend_io_cpu_status_upie),
    .io_cpu_status_mie(frontend_io_cpu_status_mie),
    .io_cpu_status_hie(frontend_io_cpu_status_hie),
    .io_cpu_status_sie(frontend_io_cpu_status_sie),
    .io_cpu_status_uie(frontend_io_cpu_status_uie),
    .io_cpu_sfence_valid(frontend_io_cpu_sfence_valid),
    .io_cpu_sfence_bits_rs1(frontend_io_cpu_sfence_bits_rs1),
    .io_cpu_sfence_bits_rs2(frontend_io_cpu_sfence_bits_rs2),
    .io_cpu_sfence_bits_addr(frontend_io_cpu_sfence_bits_addr),
    .io_cpu_sfence_bits_asid(frontend_io_cpu_sfence_bits_asid),
    .io_cpu_brupdate_b1_resolve_mask(frontend_io_cpu_brupdate_b1_resolve_mask),
    .io_cpu_brupdate_b1_mispredict_mask(frontend_io_cpu_brupdate_b1_mispredict_mask),
    .io_cpu_brupdate_b2_uop_switch(frontend_io_cpu_brupdate_b2_uop_switch),
    .io_cpu_brupdate_b2_uop_switch_off(frontend_io_cpu_brupdate_b2_uop_switch_off),
    .io_cpu_brupdate_b2_uop_is_unicore(frontend_io_cpu_brupdate_b2_uop_is_unicore),
    .io_cpu_brupdate_b2_uop_shift(frontend_io_cpu_brupdate_b2_uop_shift),
    .io_cpu_brupdate_b2_uop_lrs3_rtype(frontend_io_cpu_brupdate_b2_uop_lrs3_rtype),
    .io_cpu_brupdate_b2_uop_rflag(frontend_io_cpu_brupdate_b2_uop_rflag),
    .io_cpu_brupdate_b2_uop_wflag(frontend_io_cpu_brupdate_b2_uop_wflag),
    .io_cpu_brupdate_b2_uop_prflag(frontend_io_cpu_brupdate_b2_uop_prflag),
    .io_cpu_brupdate_b2_uop_pwflag(frontend_io_cpu_brupdate_b2_uop_pwflag),
    .io_cpu_brupdate_b2_uop_pflag_busy(frontend_io_cpu_brupdate_b2_uop_pflag_busy),
    .io_cpu_brupdate_b2_uop_stale_pflag(frontend_io_cpu_brupdate_b2_uop_stale_pflag),
    .io_cpu_brupdate_b2_uop_op1_sel(frontend_io_cpu_brupdate_b2_uop_op1_sel),
    .io_cpu_brupdate_b2_uop_op2_sel(frontend_io_cpu_brupdate_b2_uop_op2_sel),
    .io_cpu_brupdate_b2_uop_split_num(frontend_io_cpu_brupdate_b2_uop_split_num),
    .io_cpu_brupdate_b2_uop_self_index(frontend_io_cpu_brupdate_b2_uop_self_index),
    .io_cpu_brupdate_b2_uop_rob_inst_idx(frontend_io_cpu_brupdate_b2_uop_rob_inst_idx),
    .io_cpu_brupdate_b2_uop_address_num(frontend_io_cpu_brupdate_b2_uop_address_num),
    .io_cpu_brupdate_b2_uop_uopc(frontend_io_cpu_brupdate_b2_uop_uopc),
    .io_cpu_brupdate_b2_uop_inst(frontend_io_cpu_brupdate_b2_uop_inst),
    .io_cpu_brupdate_b2_uop_debug_inst(frontend_io_cpu_brupdate_b2_uop_debug_inst),
    .io_cpu_brupdate_b2_uop_is_rvc(frontend_io_cpu_brupdate_b2_uop_is_rvc),
    .io_cpu_brupdate_b2_uop_debug_pc(frontend_io_cpu_brupdate_b2_uop_debug_pc),
    .io_cpu_brupdate_b2_uop_iq_type(frontend_io_cpu_brupdate_b2_uop_iq_type),
    .io_cpu_brupdate_b2_uop_fu_code(frontend_io_cpu_brupdate_b2_uop_fu_code),
    .io_cpu_brupdate_b2_uop_ctrl_br_type(frontend_io_cpu_brupdate_b2_uop_ctrl_br_type),
    .io_cpu_brupdate_b2_uop_ctrl_op1_sel(frontend_io_cpu_brupdate_b2_uop_ctrl_op1_sel),
    .io_cpu_brupdate_b2_uop_ctrl_op2_sel(frontend_io_cpu_brupdate_b2_uop_ctrl_op2_sel),
    .io_cpu_brupdate_b2_uop_ctrl_imm_sel(frontend_io_cpu_brupdate_b2_uop_ctrl_imm_sel),
    .io_cpu_brupdate_b2_uop_ctrl_op_fcn(frontend_io_cpu_brupdate_b2_uop_ctrl_op_fcn),
    .io_cpu_brupdate_b2_uop_ctrl_fcn_dw(frontend_io_cpu_brupdate_b2_uop_ctrl_fcn_dw),
    .io_cpu_brupdate_b2_uop_ctrl_csr_cmd(frontend_io_cpu_brupdate_b2_uop_ctrl_csr_cmd),
    .io_cpu_brupdate_b2_uop_ctrl_is_load(frontend_io_cpu_brupdate_b2_uop_ctrl_is_load),
    .io_cpu_brupdate_b2_uop_ctrl_is_sta(frontend_io_cpu_brupdate_b2_uop_ctrl_is_sta),
    .io_cpu_brupdate_b2_uop_ctrl_is_std(frontend_io_cpu_brupdate_b2_uop_ctrl_is_std),
    .io_cpu_brupdate_b2_uop_ctrl_op3_sel(frontend_io_cpu_brupdate_b2_uop_ctrl_op3_sel),
    .io_cpu_brupdate_b2_uop_iw_state(frontend_io_cpu_brupdate_b2_uop_iw_state),
    .io_cpu_brupdate_b2_uop_iw_p1_poisoned(frontend_io_cpu_brupdate_b2_uop_iw_p1_poisoned),
    .io_cpu_brupdate_b2_uop_iw_p2_poisoned(frontend_io_cpu_brupdate_b2_uop_iw_p2_poisoned),
    .io_cpu_brupdate_b2_uop_is_br(frontend_io_cpu_brupdate_b2_uop_is_br),
    .io_cpu_brupdate_b2_uop_is_jalr(frontend_io_cpu_brupdate_b2_uop_is_jalr),
    .io_cpu_brupdate_b2_uop_is_jal(frontend_io_cpu_brupdate_b2_uop_is_jal),
    .io_cpu_brupdate_b2_uop_is_sfb(frontend_io_cpu_brupdate_b2_uop_is_sfb),
    .io_cpu_brupdate_b2_uop_br_mask(frontend_io_cpu_brupdate_b2_uop_br_mask),
    .io_cpu_brupdate_b2_uop_br_tag(frontend_io_cpu_brupdate_b2_uop_br_tag),
    .io_cpu_brupdate_b2_uop_ftq_idx(frontend_io_cpu_brupdate_b2_uop_ftq_idx),
    .io_cpu_brupdate_b2_uop_edge_inst(frontend_io_cpu_brupdate_b2_uop_edge_inst),
    .io_cpu_brupdate_b2_uop_pc_lob(frontend_io_cpu_brupdate_b2_uop_pc_lob),
    .io_cpu_brupdate_b2_uop_taken(frontend_io_cpu_brupdate_b2_uop_taken),
    .io_cpu_brupdate_b2_uop_imm_packed(frontend_io_cpu_brupdate_b2_uop_imm_packed),
    .io_cpu_brupdate_b2_uop_csr_addr(frontend_io_cpu_brupdate_b2_uop_csr_addr),
    .io_cpu_brupdate_b2_uop_rob_idx(frontend_io_cpu_brupdate_b2_uop_rob_idx),
    .io_cpu_brupdate_b2_uop_ldq_idx(frontend_io_cpu_brupdate_b2_uop_ldq_idx),
    .io_cpu_brupdate_b2_uop_stq_idx(frontend_io_cpu_brupdate_b2_uop_stq_idx),
    .io_cpu_brupdate_b2_uop_rxq_idx(frontend_io_cpu_brupdate_b2_uop_rxq_idx),
    .io_cpu_brupdate_b2_uop_pdst(frontend_io_cpu_brupdate_b2_uop_pdst),
    .io_cpu_brupdate_b2_uop_prs1(frontend_io_cpu_brupdate_b2_uop_prs1),
    .io_cpu_brupdate_b2_uop_prs2(frontend_io_cpu_brupdate_b2_uop_prs2),
    .io_cpu_brupdate_b2_uop_prs3(frontend_io_cpu_brupdate_b2_uop_prs3),
    .io_cpu_brupdate_b2_uop_ppred(frontend_io_cpu_brupdate_b2_uop_ppred),
    .io_cpu_brupdate_b2_uop_prs1_busy(frontend_io_cpu_brupdate_b2_uop_prs1_busy),
    .io_cpu_brupdate_b2_uop_prs2_busy(frontend_io_cpu_brupdate_b2_uop_prs2_busy),
    .io_cpu_brupdate_b2_uop_prs3_busy(frontend_io_cpu_brupdate_b2_uop_prs3_busy),
    .io_cpu_brupdate_b2_uop_ppred_busy(frontend_io_cpu_brupdate_b2_uop_ppred_busy),
    .io_cpu_brupdate_b2_uop_stale_pdst(frontend_io_cpu_brupdate_b2_uop_stale_pdst),
    .io_cpu_brupdate_b2_uop_exception(frontend_io_cpu_brupdate_b2_uop_exception),
    .io_cpu_brupdate_b2_uop_exc_cause(frontend_io_cpu_brupdate_b2_uop_exc_cause),
    .io_cpu_brupdate_b2_uop_bypassable(frontend_io_cpu_brupdate_b2_uop_bypassable),
    .io_cpu_brupdate_b2_uop_mem_cmd(frontend_io_cpu_brupdate_b2_uop_mem_cmd),
    .io_cpu_brupdate_b2_uop_mem_size(frontend_io_cpu_brupdate_b2_uop_mem_size),
    .io_cpu_brupdate_b2_uop_mem_signed(frontend_io_cpu_brupdate_b2_uop_mem_signed),
    .io_cpu_brupdate_b2_uop_is_fence(frontend_io_cpu_brupdate_b2_uop_is_fence),
    .io_cpu_brupdate_b2_uop_is_fencei(frontend_io_cpu_brupdate_b2_uop_is_fencei),
    .io_cpu_brupdate_b2_uop_is_amo(frontend_io_cpu_brupdate_b2_uop_is_amo),
    .io_cpu_brupdate_b2_uop_uses_ldq(frontend_io_cpu_brupdate_b2_uop_uses_ldq),
    .io_cpu_brupdate_b2_uop_uses_stq(frontend_io_cpu_brupdate_b2_uop_uses_stq),
    .io_cpu_brupdate_b2_uop_is_sys_pc2epc(frontend_io_cpu_brupdate_b2_uop_is_sys_pc2epc),
    .io_cpu_brupdate_b2_uop_is_unique(frontend_io_cpu_brupdate_b2_uop_is_unique),
    .io_cpu_brupdate_b2_uop_flush_on_commit(frontend_io_cpu_brupdate_b2_uop_flush_on_commit),
    .io_cpu_brupdate_b2_uop_ldst_is_rs1(frontend_io_cpu_brupdate_b2_uop_ldst_is_rs1),
    .io_cpu_brupdate_b2_uop_ldst(frontend_io_cpu_brupdate_b2_uop_ldst),
    .io_cpu_brupdate_b2_uop_lrs1(frontend_io_cpu_brupdate_b2_uop_lrs1),
    .io_cpu_brupdate_b2_uop_lrs2(frontend_io_cpu_brupdate_b2_uop_lrs2),
    .io_cpu_brupdate_b2_uop_lrs3(frontend_io_cpu_brupdate_b2_uop_lrs3),
    .io_cpu_brupdate_b2_uop_ldst_val(frontend_io_cpu_brupdate_b2_uop_ldst_val),
    .io_cpu_brupdate_b2_uop_dst_rtype(frontend_io_cpu_brupdate_b2_uop_dst_rtype),
    .io_cpu_brupdate_b2_uop_lrs1_rtype(frontend_io_cpu_brupdate_b2_uop_lrs1_rtype),
    .io_cpu_brupdate_b2_uop_lrs2_rtype(frontend_io_cpu_brupdate_b2_uop_lrs2_rtype),
    .io_cpu_brupdate_b2_uop_frs3_en(frontend_io_cpu_brupdate_b2_uop_frs3_en),
    .io_cpu_brupdate_b2_uop_fp_val(frontend_io_cpu_brupdate_b2_uop_fp_val),
    .io_cpu_brupdate_b2_uop_fp_single(frontend_io_cpu_brupdate_b2_uop_fp_single),
    .io_cpu_brupdate_b2_uop_xcpt_pf_if(frontend_io_cpu_brupdate_b2_uop_xcpt_pf_if),
    .io_cpu_brupdate_b2_uop_xcpt_ae_if(frontend_io_cpu_brupdate_b2_uop_xcpt_ae_if),
    .io_cpu_brupdate_b2_uop_xcpt_ma_if(frontend_io_cpu_brupdate_b2_uop_xcpt_ma_if),
    .io_cpu_brupdate_b2_uop_bp_debug_if(frontend_io_cpu_brupdate_b2_uop_bp_debug_if),
    .io_cpu_brupdate_b2_uop_bp_xcpt_if(frontend_io_cpu_brupdate_b2_uop_bp_xcpt_if),
    .io_cpu_brupdate_b2_uop_debug_fsrc(frontend_io_cpu_brupdate_b2_uop_debug_fsrc),
    .io_cpu_brupdate_b2_uop_debug_tsrc(frontend_io_cpu_brupdate_b2_uop_debug_tsrc),
    .io_cpu_brupdate_b2_valid(frontend_io_cpu_brupdate_b2_valid),
    .io_cpu_brupdate_b2_mispredict(frontend_io_cpu_brupdate_b2_mispredict),
    .io_cpu_brupdate_b2_taken(frontend_io_cpu_brupdate_b2_taken),
    .io_cpu_brupdate_b2_cfi_type(frontend_io_cpu_brupdate_b2_cfi_type),
    .io_cpu_brupdate_b2_pc_sel(frontend_io_cpu_brupdate_b2_pc_sel),
    .io_cpu_brupdate_b2_jalr_target(frontend_io_cpu_brupdate_b2_jalr_target),
    .io_cpu_brupdate_b2_target_offset(frontend_io_cpu_brupdate_b2_target_offset),
    .io_cpu_redirect_flush(frontend_io_cpu_redirect_flush),
    .io_cpu_redirect_val(frontend_io_cpu_redirect_val),
    .io_cpu_redirect_pc(frontend_io_cpu_redirect_pc),
    .io_cpu_redirect_ftq_idx(frontend_io_cpu_redirect_ftq_idx),
    .io_cpu_redirect_ghist_old_history(frontend_io_cpu_redirect_ghist_old_history),
    .io_cpu_redirect_ghist_current_saw_branch_not_taken(frontend_io_cpu_redirect_ghist_current_saw_branch_not_taken),
    .io_cpu_redirect_ghist_new_saw_branch_not_taken(frontend_io_cpu_redirect_ghist_new_saw_branch_not_taken),
    .io_cpu_redirect_ghist_new_saw_branch_taken(frontend_io_cpu_redirect_ghist_new_saw_branch_taken),
    .io_cpu_redirect_ghist_ras_idx(frontend_io_cpu_redirect_ghist_ras_idx),
    .io_cpu_commit_valid(frontend_io_cpu_commit_valid),
    .io_cpu_commit_bits(frontend_io_cpu_commit_bits),
    .io_cpu_flush_icache(frontend_io_cpu_flush_icache),
    .io_cpu_perf_acquire(frontend_io_cpu_perf_acquire),
    .io_cpu_perf_tlbMiss(frontend_io_cpu_perf_tlbMiss),
    .io_cpu_is_unicore(frontend_io_cpu_is_unicore),
    .io_ptw_req_ready(frontend_io_ptw_req_ready),
    .io_ptw_req_valid(frontend_io_ptw_req_valid),
    .io_ptw_req_bits_valid(frontend_io_ptw_req_bits_valid),
    .io_ptw_req_bits_bits_addr(frontend_io_ptw_req_bits_bits_addr),
    .io_ptw_resp_valid(frontend_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae(frontend_io_ptw_resp_bits_ae),
    .io_ptw_resp_bits_pte_ppn(frontend_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(frontend_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(frontend_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(frontend_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(frontend_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(frontend_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(frontend_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(frontend_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(frontend_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(frontend_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(frontend_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_fragmented_superpage(frontend_io_ptw_resp_bits_fragmented_superpage),
    .io_ptw_resp_bits_homogeneous(frontend_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(frontend_io_ptw_ptbr_mode),
    .io_ptw_ptbr_asid(frontend_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(frontend_io_ptw_ptbr_ppn),
    .io_ptw_status_debug(frontend_io_ptw_status_debug),
    .io_ptw_status_cease(frontend_io_ptw_status_cease),
    .io_ptw_status_wfi(frontend_io_ptw_status_wfi),
    .io_ptw_status_isa(frontend_io_ptw_status_isa),
    .io_ptw_status_dprv(frontend_io_ptw_status_dprv),
    .io_ptw_status_prv(frontend_io_ptw_status_prv),
    .io_ptw_status_sd(frontend_io_ptw_status_sd),
    .io_ptw_status_zero2(frontend_io_ptw_status_zero2),
    .io_ptw_status_sxl(frontend_io_ptw_status_sxl),
    .io_ptw_status_uxl(frontend_io_ptw_status_uxl),
    .io_ptw_status_sd_rv32(frontend_io_ptw_status_sd_rv32),
    .io_ptw_status_zero1(frontend_io_ptw_status_zero1),
    .io_ptw_status_tsr(frontend_io_ptw_status_tsr),
    .io_ptw_status_tw(frontend_io_ptw_status_tw),
    .io_ptw_status_tvm(frontend_io_ptw_status_tvm),
    .io_ptw_status_mxr(frontend_io_ptw_status_mxr),
    .io_ptw_status_sum(frontend_io_ptw_status_sum),
    .io_ptw_status_mprv(frontend_io_ptw_status_mprv),
    .io_ptw_status_xs(frontend_io_ptw_status_xs),
    .io_ptw_status_fs(frontend_io_ptw_status_fs),
    .io_ptw_status_mpp(frontend_io_ptw_status_mpp),
    .io_ptw_status_vs(frontend_io_ptw_status_vs),
    .io_ptw_status_spp(frontend_io_ptw_status_spp),
    .io_ptw_status_mpie(frontend_io_ptw_status_mpie),
    .io_ptw_status_hpie(frontend_io_ptw_status_hpie),
    .io_ptw_status_spie(frontend_io_ptw_status_spie),
    .io_ptw_status_upie(frontend_io_ptw_status_upie),
    .io_ptw_status_mie(frontend_io_ptw_status_mie),
    .io_ptw_status_hie(frontend_io_ptw_status_hie),
    .io_ptw_status_sie(frontend_io_ptw_status_sie),
    .io_ptw_status_uie(frontend_io_ptw_status_uie),
    .io_ptw_pmp_0_cfg_l(frontend_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_res(frontend_io_ptw_pmp_0_cfg_res),
    .io_ptw_pmp_0_cfg_a(frontend_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(frontend_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(frontend_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(frontend_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(frontend_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(frontend_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(frontend_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_res(frontend_io_ptw_pmp_1_cfg_res),
    .io_ptw_pmp_1_cfg_a(frontend_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(frontend_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(frontend_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(frontend_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(frontend_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(frontend_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(frontend_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_res(frontend_io_ptw_pmp_2_cfg_res),
    .io_ptw_pmp_2_cfg_a(frontend_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(frontend_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(frontend_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(frontend_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(frontend_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(frontend_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(frontend_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_res(frontend_io_ptw_pmp_3_cfg_res),
    .io_ptw_pmp_3_cfg_a(frontend_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(frontend_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(frontend_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(frontend_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(frontend_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(frontend_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(frontend_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_res(frontend_io_ptw_pmp_4_cfg_res),
    .io_ptw_pmp_4_cfg_a(frontend_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(frontend_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(frontend_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(frontend_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(frontend_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(frontend_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(frontend_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_res(frontend_io_ptw_pmp_5_cfg_res),
    .io_ptw_pmp_5_cfg_a(frontend_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(frontend_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(frontend_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(frontend_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(frontend_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(frontend_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(frontend_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_res(frontend_io_ptw_pmp_6_cfg_res),
    .io_ptw_pmp_6_cfg_a(frontend_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(frontend_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(frontend_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(frontend_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(frontend_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(frontend_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(frontend_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_res(frontend_io_ptw_pmp_7_cfg_res),
    .io_ptw_pmp_7_cfg_a(frontend_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(frontend_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(frontend_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(frontend_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(frontend_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(frontend_io_ptw_pmp_7_mask),
    .io_ptw_customCSRs_csrs_0_wen(frontend_io_ptw_customCSRs_csrs_0_wen),
    .io_ptw_customCSRs_csrs_0_wdata(frontend_io_ptw_customCSRs_csrs_0_wdata),
    .io_ptw_customCSRs_csrs_0_value(frontend_io_ptw_customCSRs_csrs_0_value),
    .io_errors_bus_valid(frontend_io_errors_bus_valid),
    .io_errors_bus_bits(frontend_io_errors_bus_bits)
  );
  BoomCore core ( // @[tile.scala 159:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_hartid(core_io_hartid),
    .io_interrupts_debug(core_io_interrupts_debug),
    .io_interrupts_mtip(core_io_interrupts_mtip),
    .io_interrupts_msip(core_io_interrupts_msip),
    .io_interrupts_meip(core_io_interrupts_meip),
    .io_interrupts_seip(core_io_interrupts_seip),
    .io_ifu_fetchpacket_ready(core_io_ifu_fetchpacket_ready),
    .io_ifu_fetchpacket_valid(core_io_ifu_fetchpacket_valid),
    .io_ifu_fetchpacket_bits_uops_0_valid(core_io_ifu_fetchpacket_bits_uops_0_valid),
    .io_ifu_fetchpacket_bits_uops_0_bits_switch(core_io_ifu_fetchpacket_bits_uops_0_bits_switch),
    .io_ifu_fetchpacket_bits_uops_0_bits_switch_off(core_io_ifu_fetchpacket_bits_uops_0_bits_switch_off),
    .io_ifu_fetchpacket_bits_uops_0_bits_is_unicore(core_io_ifu_fetchpacket_bits_uops_0_bits_is_unicore),
    .io_ifu_fetchpacket_bits_uops_0_bits_shift(core_io_ifu_fetchpacket_bits_uops_0_bits_shift),
    .io_ifu_fetchpacket_bits_uops_0_bits_lrs3_rtype(core_io_ifu_fetchpacket_bits_uops_0_bits_lrs3_rtype),
    .io_ifu_fetchpacket_bits_uops_0_bits_rflag(core_io_ifu_fetchpacket_bits_uops_0_bits_rflag),
    .io_ifu_fetchpacket_bits_uops_0_bits_wflag(core_io_ifu_fetchpacket_bits_uops_0_bits_wflag),
    .io_ifu_fetchpacket_bits_uops_0_bits_prflag(core_io_ifu_fetchpacket_bits_uops_0_bits_prflag),
    .io_ifu_fetchpacket_bits_uops_0_bits_pwflag(core_io_ifu_fetchpacket_bits_uops_0_bits_pwflag),
    .io_ifu_fetchpacket_bits_uops_0_bits_pflag_busy(core_io_ifu_fetchpacket_bits_uops_0_bits_pflag_busy),
    .io_ifu_fetchpacket_bits_uops_0_bits_stale_pflag(core_io_ifu_fetchpacket_bits_uops_0_bits_stale_pflag),
    .io_ifu_fetchpacket_bits_uops_0_bits_op1_sel(core_io_ifu_fetchpacket_bits_uops_0_bits_op1_sel),
    .io_ifu_fetchpacket_bits_uops_0_bits_op2_sel(core_io_ifu_fetchpacket_bits_uops_0_bits_op2_sel),
    .io_ifu_fetchpacket_bits_uops_0_bits_split_num(core_io_ifu_fetchpacket_bits_uops_0_bits_split_num),
    .io_ifu_fetchpacket_bits_uops_0_bits_self_index(core_io_ifu_fetchpacket_bits_uops_0_bits_self_index),
    .io_ifu_fetchpacket_bits_uops_0_bits_rob_inst_idx(core_io_ifu_fetchpacket_bits_uops_0_bits_rob_inst_idx),
    .io_ifu_fetchpacket_bits_uops_0_bits_address_num(core_io_ifu_fetchpacket_bits_uops_0_bits_address_num),
    .io_ifu_fetchpacket_bits_uops_0_bits_uopc(core_io_ifu_fetchpacket_bits_uops_0_bits_uopc),
    .io_ifu_fetchpacket_bits_uops_0_bits_inst(core_io_ifu_fetchpacket_bits_uops_0_bits_inst),
    .io_ifu_fetchpacket_bits_uops_0_bits_debug_inst(core_io_ifu_fetchpacket_bits_uops_0_bits_debug_inst),
    .io_ifu_fetchpacket_bits_uops_0_bits_is_rvc(core_io_ifu_fetchpacket_bits_uops_0_bits_is_rvc),
    .io_ifu_fetchpacket_bits_uops_0_bits_debug_pc(core_io_ifu_fetchpacket_bits_uops_0_bits_debug_pc),
    .io_ifu_fetchpacket_bits_uops_0_bits_iq_type(core_io_ifu_fetchpacket_bits_uops_0_bits_iq_type),
    .io_ifu_fetchpacket_bits_uops_0_bits_fu_code(core_io_ifu_fetchpacket_bits_uops_0_bits_fu_code),
    .io_ifu_fetchpacket_bits_uops_0_bits_ctrl_br_type(core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_br_type),
    .io_ifu_fetchpacket_bits_uops_0_bits_ctrl_op1_sel(core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_op1_sel),
    .io_ifu_fetchpacket_bits_uops_0_bits_ctrl_op2_sel(core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_op2_sel),
    .io_ifu_fetchpacket_bits_uops_0_bits_ctrl_imm_sel(core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_imm_sel),
    .io_ifu_fetchpacket_bits_uops_0_bits_ctrl_op_fcn(core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_op_fcn),
    .io_ifu_fetchpacket_bits_uops_0_bits_ctrl_fcn_dw(core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_fcn_dw),
    .io_ifu_fetchpacket_bits_uops_0_bits_ctrl_csr_cmd(core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_csr_cmd),
    .io_ifu_fetchpacket_bits_uops_0_bits_ctrl_is_load(core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_is_load),
    .io_ifu_fetchpacket_bits_uops_0_bits_ctrl_is_sta(core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_is_sta),
    .io_ifu_fetchpacket_bits_uops_0_bits_ctrl_is_std(core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_is_std),
    .io_ifu_fetchpacket_bits_uops_0_bits_ctrl_op3_sel(core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_op3_sel),
    .io_ifu_fetchpacket_bits_uops_0_bits_iw_state(core_io_ifu_fetchpacket_bits_uops_0_bits_iw_state),
    .io_ifu_fetchpacket_bits_uops_0_bits_iw_p1_poisoned(core_io_ifu_fetchpacket_bits_uops_0_bits_iw_p1_poisoned),
    .io_ifu_fetchpacket_bits_uops_0_bits_iw_p2_poisoned(core_io_ifu_fetchpacket_bits_uops_0_bits_iw_p2_poisoned),
    .io_ifu_fetchpacket_bits_uops_0_bits_is_br(core_io_ifu_fetchpacket_bits_uops_0_bits_is_br),
    .io_ifu_fetchpacket_bits_uops_0_bits_is_jalr(core_io_ifu_fetchpacket_bits_uops_0_bits_is_jalr),
    .io_ifu_fetchpacket_bits_uops_0_bits_is_jal(core_io_ifu_fetchpacket_bits_uops_0_bits_is_jal),
    .io_ifu_fetchpacket_bits_uops_0_bits_is_sfb(core_io_ifu_fetchpacket_bits_uops_0_bits_is_sfb),
    .io_ifu_fetchpacket_bits_uops_0_bits_br_mask(core_io_ifu_fetchpacket_bits_uops_0_bits_br_mask),
    .io_ifu_fetchpacket_bits_uops_0_bits_br_tag(core_io_ifu_fetchpacket_bits_uops_0_bits_br_tag),
    .io_ifu_fetchpacket_bits_uops_0_bits_ftq_idx(core_io_ifu_fetchpacket_bits_uops_0_bits_ftq_idx),
    .io_ifu_fetchpacket_bits_uops_0_bits_edge_inst(core_io_ifu_fetchpacket_bits_uops_0_bits_edge_inst),
    .io_ifu_fetchpacket_bits_uops_0_bits_pc_lob(core_io_ifu_fetchpacket_bits_uops_0_bits_pc_lob),
    .io_ifu_fetchpacket_bits_uops_0_bits_taken(core_io_ifu_fetchpacket_bits_uops_0_bits_taken),
    .io_ifu_fetchpacket_bits_uops_0_bits_imm_packed(core_io_ifu_fetchpacket_bits_uops_0_bits_imm_packed),
    .io_ifu_fetchpacket_bits_uops_0_bits_csr_addr(core_io_ifu_fetchpacket_bits_uops_0_bits_csr_addr),
    .io_ifu_fetchpacket_bits_uops_0_bits_rob_idx(core_io_ifu_fetchpacket_bits_uops_0_bits_rob_idx),
    .io_ifu_fetchpacket_bits_uops_0_bits_ldq_idx(core_io_ifu_fetchpacket_bits_uops_0_bits_ldq_idx),
    .io_ifu_fetchpacket_bits_uops_0_bits_stq_idx(core_io_ifu_fetchpacket_bits_uops_0_bits_stq_idx),
    .io_ifu_fetchpacket_bits_uops_0_bits_rxq_idx(core_io_ifu_fetchpacket_bits_uops_0_bits_rxq_idx),
    .io_ifu_fetchpacket_bits_uops_0_bits_pdst(core_io_ifu_fetchpacket_bits_uops_0_bits_pdst),
    .io_ifu_fetchpacket_bits_uops_0_bits_prs1(core_io_ifu_fetchpacket_bits_uops_0_bits_prs1),
    .io_ifu_fetchpacket_bits_uops_0_bits_prs2(core_io_ifu_fetchpacket_bits_uops_0_bits_prs2),
    .io_ifu_fetchpacket_bits_uops_0_bits_prs3(core_io_ifu_fetchpacket_bits_uops_0_bits_prs3),
    .io_ifu_fetchpacket_bits_uops_0_bits_ppred(core_io_ifu_fetchpacket_bits_uops_0_bits_ppred),
    .io_ifu_fetchpacket_bits_uops_0_bits_prs1_busy(core_io_ifu_fetchpacket_bits_uops_0_bits_prs1_busy),
    .io_ifu_fetchpacket_bits_uops_0_bits_prs2_busy(core_io_ifu_fetchpacket_bits_uops_0_bits_prs2_busy),
    .io_ifu_fetchpacket_bits_uops_0_bits_prs3_busy(core_io_ifu_fetchpacket_bits_uops_0_bits_prs3_busy),
    .io_ifu_fetchpacket_bits_uops_0_bits_ppred_busy(core_io_ifu_fetchpacket_bits_uops_0_bits_ppred_busy),
    .io_ifu_fetchpacket_bits_uops_0_bits_stale_pdst(core_io_ifu_fetchpacket_bits_uops_0_bits_stale_pdst),
    .io_ifu_fetchpacket_bits_uops_0_bits_exception(core_io_ifu_fetchpacket_bits_uops_0_bits_exception),
    .io_ifu_fetchpacket_bits_uops_0_bits_exc_cause(core_io_ifu_fetchpacket_bits_uops_0_bits_exc_cause),
    .io_ifu_fetchpacket_bits_uops_0_bits_bypassable(core_io_ifu_fetchpacket_bits_uops_0_bits_bypassable),
    .io_ifu_fetchpacket_bits_uops_0_bits_mem_cmd(core_io_ifu_fetchpacket_bits_uops_0_bits_mem_cmd),
    .io_ifu_fetchpacket_bits_uops_0_bits_mem_size(core_io_ifu_fetchpacket_bits_uops_0_bits_mem_size),
    .io_ifu_fetchpacket_bits_uops_0_bits_mem_signed(core_io_ifu_fetchpacket_bits_uops_0_bits_mem_signed),
    .io_ifu_fetchpacket_bits_uops_0_bits_is_fence(core_io_ifu_fetchpacket_bits_uops_0_bits_is_fence),
    .io_ifu_fetchpacket_bits_uops_0_bits_is_fencei(core_io_ifu_fetchpacket_bits_uops_0_bits_is_fencei),
    .io_ifu_fetchpacket_bits_uops_0_bits_is_amo(core_io_ifu_fetchpacket_bits_uops_0_bits_is_amo),
    .io_ifu_fetchpacket_bits_uops_0_bits_uses_ldq(core_io_ifu_fetchpacket_bits_uops_0_bits_uses_ldq),
    .io_ifu_fetchpacket_bits_uops_0_bits_uses_stq(core_io_ifu_fetchpacket_bits_uops_0_bits_uses_stq),
    .io_ifu_fetchpacket_bits_uops_0_bits_is_sys_pc2epc(core_io_ifu_fetchpacket_bits_uops_0_bits_is_sys_pc2epc),
    .io_ifu_fetchpacket_bits_uops_0_bits_is_unique(core_io_ifu_fetchpacket_bits_uops_0_bits_is_unique),
    .io_ifu_fetchpacket_bits_uops_0_bits_flush_on_commit(core_io_ifu_fetchpacket_bits_uops_0_bits_flush_on_commit),
    .io_ifu_fetchpacket_bits_uops_0_bits_ldst_is_rs1(core_io_ifu_fetchpacket_bits_uops_0_bits_ldst_is_rs1),
    .io_ifu_fetchpacket_bits_uops_0_bits_ldst(core_io_ifu_fetchpacket_bits_uops_0_bits_ldst),
    .io_ifu_fetchpacket_bits_uops_0_bits_lrs1(core_io_ifu_fetchpacket_bits_uops_0_bits_lrs1),
    .io_ifu_fetchpacket_bits_uops_0_bits_lrs2(core_io_ifu_fetchpacket_bits_uops_0_bits_lrs2),
    .io_ifu_fetchpacket_bits_uops_0_bits_lrs3(core_io_ifu_fetchpacket_bits_uops_0_bits_lrs3),
    .io_ifu_fetchpacket_bits_uops_0_bits_ldst_val(core_io_ifu_fetchpacket_bits_uops_0_bits_ldst_val),
    .io_ifu_fetchpacket_bits_uops_0_bits_dst_rtype(core_io_ifu_fetchpacket_bits_uops_0_bits_dst_rtype),
    .io_ifu_fetchpacket_bits_uops_0_bits_lrs1_rtype(core_io_ifu_fetchpacket_bits_uops_0_bits_lrs1_rtype),
    .io_ifu_fetchpacket_bits_uops_0_bits_lrs2_rtype(core_io_ifu_fetchpacket_bits_uops_0_bits_lrs2_rtype),
    .io_ifu_fetchpacket_bits_uops_0_bits_frs3_en(core_io_ifu_fetchpacket_bits_uops_0_bits_frs3_en),
    .io_ifu_fetchpacket_bits_uops_0_bits_fp_val(core_io_ifu_fetchpacket_bits_uops_0_bits_fp_val),
    .io_ifu_fetchpacket_bits_uops_0_bits_fp_single(core_io_ifu_fetchpacket_bits_uops_0_bits_fp_single),
    .io_ifu_fetchpacket_bits_uops_0_bits_xcpt_pf_if(core_io_ifu_fetchpacket_bits_uops_0_bits_xcpt_pf_if),
    .io_ifu_fetchpacket_bits_uops_0_bits_xcpt_ae_if(core_io_ifu_fetchpacket_bits_uops_0_bits_xcpt_ae_if),
    .io_ifu_fetchpacket_bits_uops_0_bits_xcpt_ma_if(core_io_ifu_fetchpacket_bits_uops_0_bits_xcpt_ma_if),
    .io_ifu_fetchpacket_bits_uops_0_bits_bp_debug_if(core_io_ifu_fetchpacket_bits_uops_0_bits_bp_debug_if),
    .io_ifu_fetchpacket_bits_uops_0_bits_bp_xcpt_if(core_io_ifu_fetchpacket_bits_uops_0_bits_bp_xcpt_if),
    .io_ifu_fetchpacket_bits_uops_0_bits_debug_fsrc(core_io_ifu_fetchpacket_bits_uops_0_bits_debug_fsrc),
    .io_ifu_fetchpacket_bits_uops_0_bits_debug_tsrc(core_io_ifu_fetchpacket_bits_uops_0_bits_debug_tsrc),
    .io_ifu_fetchpacket_bits_uops_1_valid(core_io_ifu_fetchpacket_bits_uops_1_valid),
    .io_ifu_fetchpacket_bits_uops_1_bits_switch(core_io_ifu_fetchpacket_bits_uops_1_bits_switch),
    .io_ifu_fetchpacket_bits_uops_1_bits_switch_off(core_io_ifu_fetchpacket_bits_uops_1_bits_switch_off),
    .io_ifu_fetchpacket_bits_uops_1_bits_is_unicore(core_io_ifu_fetchpacket_bits_uops_1_bits_is_unicore),
    .io_ifu_fetchpacket_bits_uops_1_bits_shift(core_io_ifu_fetchpacket_bits_uops_1_bits_shift),
    .io_ifu_fetchpacket_bits_uops_1_bits_lrs3_rtype(core_io_ifu_fetchpacket_bits_uops_1_bits_lrs3_rtype),
    .io_ifu_fetchpacket_bits_uops_1_bits_rflag(core_io_ifu_fetchpacket_bits_uops_1_bits_rflag),
    .io_ifu_fetchpacket_bits_uops_1_bits_wflag(core_io_ifu_fetchpacket_bits_uops_1_bits_wflag),
    .io_ifu_fetchpacket_bits_uops_1_bits_prflag(core_io_ifu_fetchpacket_bits_uops_1_bits_prflag),
    .io_ifu_fetchpacket_bits_uops_1_bits_pwflag(core_io_ifu_fetchpacket_bits_uops_1_bits_pwflag),
    .io_ifu_fetchpacket_bits_uops_1_bits_pflag_busy(core_io_ifu_fetchpacket_bits_uops_1_bits_pflag_busy),
    .io_ifu_fetchpacket_bits_uops_1_bits_stale_pflag(core_io_ifu_fetchpacket_bits_uops_1_bits_stale_pflag),
    .io_ifu_fetchpacket_bits_uops_1_bits_op1_sel(core_io_ifu_fetchpacket_bits_uops_1_bits_op1_sel),
    .io_ifu_fetchpacket_bits_uops_1_bits_op2_sel(core_io_ifu_fetchpacket_bits_uops_1_bits_op2_sel),
    .io_ifu_fetchpacket_bits_uops_1_bits_split_num(core_io_ifu_fetchpacket_bits_uops_1_bits_split_num),
    .io_ifu_fetchpacket_bits_uops_1_bits_self_index(core_io_ifu_fetchpacket_bits_uops_1_bits_self_index),
    .io_ifu_fetchpacket_bits_uops_1_bits_rob_inst_idx(core_io_ifu_fetchpacket_bits_uops_1_bits_rob_inst_idx),
    .io_ifu_fetchpacket_bits_uops_1_bits_address_num(core_io_ifu_fetchpacket_bits_uops_1_bits_address_num),
    .io_ifu_fetchpacket_bits_uops_1_bits_uopc(core_io_ifu_fetchpacket_bits_uops_1_bits_uopc),
    .io_ifu_fetchpacket_bits_uops_1_bits_inst(core_io_ifu_fetchpacket_bits_uops_1_bits_inst),
    .io_ifu_fetchpacket_bits_uops_1_bits_debug_inst(core_io_ifu_fetchpacket_bits_uops_1_bits_debug_inst),
    .io_ifu_fetchpacket_bits_uops_1_bits_is_rvc(core_io_ifu_fetchpacket_bits_uops_1_bits_is_rvc),
    .io_ifu_fetchpacket_bits_uops_1_bits_debug_pc(core_io_ifu_fetchpacket_bits_uops_1_bits_debug_pc),
    .io_ifu_fetchpacket_bits_uops_1_bits_iq_type(core_io_ifu_fetchpacket_bits_uops_1_bits_iq_type),
    .io_ifu_fetchpacket_bits_uops_1_bits_fu_code(core_io_ifu_fetchpacket_bits_uops_1_bits_fu_code),
    .io_ifu_fetchpacket_bits_uops_1_bits_ctrl_br_type(core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_br_type),
    .io_ifu_fetchpacket_bits_uops_1_bits_ctrl_op1_sel(core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_op1_sel),
    .io_ifu_fetchpacket_bits_uops_1_bits_ctrl_op2_sel(core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_op2_sel),
    .io_ifu_fetchpacket_bits_uops_1_bits_ctrl_imm_sel(core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_imm_sel),
    .io_ifu_fetchpacket_bits_uops_1_bits_ctrl_op_fcn(core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_op_fcn),
    .io_ifu_fetchpacket_bits_uops_1_bits_ctrl_fcn_dw(core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_fcn_dw),
    .io_ifu_fetchpacket_bits_uops_1_bits_ctrl_csr_cmd(core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_csr_cmd),
    .io_ifu_fetchpacket_bits_uops_1_bits_ctrl_is_load(core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_is_load),
    .io_ifu_fetchpacket_bits_uops_1_bits_ctrl_is_sta(core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_is_sta),
    .io_ifu_fetchpacket_bits_uops_1_bits_ctrl_is_std(core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_is_std),
    .io_ifu_fetchpacket_bits_uops_1_bits_ctrl_op3_sel(core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_op3_sel),
    .io_ifu_fetchpacket_bits_uops_1_bits_iw_state(core_io_ifu_fetchpacket_bits_uops_1_bits_iw_state),
    .io_ifu_fetchpacket_bits_uops_1_bits_iw_p1_poisoned(core_io_ifu_fetchpacket_bits_uops_1_bits_iw_p1_poisoned),
    .io_ifu_fetchpacket_bits_uops_1_bits_iw_p2_poisoned(core_io_ifu_fetchpacket_bits_uops_1_bits_iw_p2_poisoned),
    .io_ifu_fetchpacket_bits_uops_1_bits_is_br(core_io_ifu_fetchpacket_bits_uops_1_bits_is_br),
    .io_ifu_fetchpacket_bits_uops_1_bits_is_jalr(core_io_ifu_fetchpacket_bits_uops_1_bits_is_jalr),
    .io_ifu_fetchpacket_bits_uops_1_bits_is_jal(core_io_ifu_fetchpacket_bits_uops_1_bits_is_jal),
    .io_ifu_fetchpacket_bits_uops_1_bits_is_sfb(core_io_ifu_fetchpacket_bits_uops_1_bits_is_sfb),
    .io_ifu_fetchpacket_bits_uops_1_bits_br_mask(core_io_ifu_fetchpacket_bits_uops_1_bits_br_mask),
    .io_ifu_fetchpacket_bits_uops_1_bits_br_tag(core_io_ifu_fetchpacket_bits_uops_1_bits_br_tag),
    .io_ifu_fetchpacket_bits_uops_1_bits_ftq_idx(core_io_ifu_fetchpacket_bits_uops_1_bits_ftq_idx),
    .io_ifu_fetchpacket_bits_uops_1_bits_edge_inst(core_io_ifu_fetchpacket_bits_uops_1_bits_edge_inst),
    .io_ifu_fetchpacket_bits_uops_1_bits_pc_lob(core_io_ifu_fetchpacket_bits_uops_1_bits_pc_lob),
    .io_ifu_fetchpacket_bits_uops_1_bits_taken(core_io_ifu_fetchpacket_bits_uops_1_bits_taken),
    .io_ifu_fetchpacket_bits_uops_1_bits_imm_packed(core_io_ifu_fetchpacket_bits_uops_1_bits_imm_packed),
    .io_ifu_fetchpacket_bits_uops_1_bits_csr_addr(core_io_ifu_fetchpacket_bits_uops_1_bits_csr_addr),
    .io_ifu_fetchpacket_bits_uops_1_bits_rob_idx(core_io_ifu_fetchpacket_bits_uops_1_bits_rob_idx),
    .io_ifu_fetchpacket_bits_uops_1_bits_ldq_idx(core_io_ifu_fetchpacket_bits_uops_1_bits_ldq_idx),
    .io_ifu_fetchpacket_bits_uops_1_bits_stq_idx(core_io_ifu_fetchpacket_bits_uops_1_bits_stq_idx),
    .io_ifu_fetchpacket_bits_uops_1_bits_rxq_idx(core_io_ifu_fetchpacket_bits_uops_1_bits_rxq_idx),
    .io_ifu_fetchpacket_bits_uops_1_bits_pdst(core_io_ifu_fetchpacket_bits_uops_1_bits_pdst),
    .io_ifu_fetchpacket_bits_uops_1_bits_prs1(core_io_ifu_fetchpacket_bits_uops_1_bits_prs1),
    .io_ifu_fetchpacket_bits_uops_1_bits_prs2(core_io_ifu_fetchpacket_bits_uops_1_bits_prs2),
    .io_ifu_fetchpacket_bits_uops_1_bits_prs3(core_io_ifu_fetchpacket_bits_uops_1_bits_prs3),
    .io_ifu_fetchpacket_bits_uops_1_bits_ppred(core_io_ifu_fetchpacket_bits_uops_1_bits_ppred),
    .io_ifu_fetchpacket_bits_uops_1_bits_prs1_busy(core_io_ifu_fetchpacket_bits_uops_1_bits_prs1_busy),
    .io_ifu_fetchpacket_bits_uops_1_bits_prs2_busy(core_io_ifu_fetchpacket_bits_uops_1_bits_prs2_busy),
    .io_ifu_fetchpacket_bits_uops_1_bits_prs3_busy(core_io_ifu_fetchpacket_bits_uops_1_bits_prs3_busy),
    .io_ifu_fetchpacket_bits_uops_1_bits_ppred_busy(core_io_ifu_fetchpacket_bits_uops_1_bits_ppred_busy),
    .io_ifu_fetchpacket_bits_uops_1_bits_stale_pdst(core_io_ifu_fetchpacket_bits_uops_1_bits_stale_pdst),
    .io_ifu_fetchpacket_bits_uops_1_bits_exception(core_io_ifu_fetchpacket_bits_uops_1_bits_exception),
    .io_ifu_fetchpacket_bits_uops_1_bits_exc_cause(core_io_ifu_fetchpacket_bits_uops_1_bits_exc_cause),
    .io_ifu_fetchpacket_bits_uops_1_bits_bypassable(core_io_ifu_fetchpacket_bits_uops_1_bits_bypassable),
    .io_ifu_fetchpacket_bits_uops_1_bits_mem_cmd(core_io_ifu_fetchpacket_bits_uops_1_bits_mem_cmd),
    .io_ifu_fetchpacket_bits_uops_1_bits_mem_size(core_io_ifu_fetchpacket_bits_uops_1_bits_mem_size),
    .io_ifu_fetchpacket_bits_uops_1_bits_mem_signed(core_io_ifu_fetchpacket_bits_uops_1_bits_mem_signed),
    .io_ifu_fetchpacket_bits_uops_1_bits_is_fence(core_io_ifu_fetchpacket_bits_uops_1_bits_is_fence),
    .io_ifu_fetchpacket_bits_uops_1_bits_is_fencei(core_io_ifu_fetchpacket_bits_uops_1_bits_is_fencei),
    .io_ifu_fetchpacket_bits_uops_1_bits_is_amo(core_io_ifu_fetchpacket_bits_uops_1_bits_is_amo),
    .io_ifu_fetchpacket_bits_uops_1_bits_uses_ldq(core_io_ifu_fetchpacket_bits_uops_1_bits_uses_ldq),
    .io_ifu_fetchpacket_bits_uops_1_bits_uses_stq(core_io_ifu_fetchpacket_bits_uops_1_bits_uses_stq),
    .io_ifu_fetchpacket_bits_uops_1_bits_is_sys_pc2epc(core_io_ifu_fetchpacket_bits_uops_1_bits_is_sys_pc2epc),
    .io_ifu_fetchpacket_bits_uops_1_bits_is_unique(core_io_ifu_fetchpacket_bits_uops_1_bits_is_unique),
    .io_ifu_fetchpacket_bits_uops_1_bits_flush_on_commit(core_io_ifu_fetchpacket_bits_uops_1_bits_flush_on_commit),
    .io_ifu_fetchpacket_bits_uops_1_bits_ldst_is_rs1(core_io_ifu_fetchpacket_bits_uops_1_bits_ldst_is_rs1),
    .io_ifu_fetchpacket_bits_uops_1_bits_ldst(core_io_ifu_fetchpacket_bits_uops_1_bits_ldst),
    .io_ifu_fetchpacket_bits_uops_1_bits_lrs1(core_io_ifu_fetchpacket_bits_uops_1_bits_lrs1),
    .io_ifu_fetchpacket_bits_uops_1_bits_lrs2(core_io_ifu_fetchpacket_bits_uops_1_bits_lrs2),
    .io_ifu_fetchpacket_bits_uops_1_bits_lrs3(core_io_ifu_fetchpacket_bits_uops_1_bits_lrs3),
    .io_ifu_fetchpacket_bits_uops_1_bits_ldst_val(core_io_ifu_fetchpacket_bits_uops_1_bits_ldst_val),
    .io_ifu_fetchpacket_bits_uops_1_bits_dst_rtype(core_io_ifu_fetchpacket_bits_uops_1_bits_dst_rtype),
    .io_ifu_fetchpacket_bits_uops_1_bits_lrs1_rtype(core_io_ifu_fetchpacket_bits_uops_1_bits_lrs1_rtype),
    .io_ifu_fetchpacket_bits_uops_1_bits_lrs2_rtype(core_io_ifu_fetchpacket_bits_uops_1_bits_lrs2_rtype),
    .io_ifu_fetchpacket_bits_uops_1_bits_frs3_en(core_io_ifu_fetchpacket_bits_uops_1_bits_frs3_en),
    .io_ifu_fetchpacket_bits_uops_1_bits_fp_val(core_io_ifu_fetchpacket_bits_uops_1_bits_fp_val),
    .io_ifu_fetchpacket_bits_uops_1_bits_fp_single(core_io_ifu_fetchpacket_bits_uops_1_bits_fp_single),
    .io_ifu_fetchpacket_bits_uops_1_bits_xcpt_pf_if(core_io_ifu_fetchpacket_bits_uops_1_bits_xcpt_pf_if),
    .io_ifu_fetchpacket_bits_uops_1_bits_xcpt_ae_if(core_io_ifu_fetchpacket_bits_uops_1_bits_xcpt_ae_if),
    .io_ifu_fetchpacket_bits_uops_1_bits_xcpt_ma_if(core_io_ifu_fetchpacket_bits_uops_1_bits_xcpt_ma_if),
    .io_ifu_fetchpacket_bits_uops_1_bits_bp_debug_if(core_io_ifu_fetchpacket_bits_uops_1_bits_bp_debug_if),
    .io_ifu_fetchpacket_bits_uops_1_bits_bp_xcpt_if(core_io_ifu_fetchpacket_bits_uops_1_bits_bp_xcpt_if),
    .io_ifu_fetchpacket_bits_uops_1_bits_debug_fsrc(core_io_ifu_fetchpacket_bits_uops_1_bits_debug_fsrc),
    .io_ifu_fetchpacket_bits_uops_1_bits_debug_tsrc(core_io_ifu_fetchpacket_bits_uops_1_bits_debug_tsrc),
    .io_ifu_get_pc_0_ftq_idx(core_io_ifu_get_pc_0_ftq_idx),
    .io_ifu_get_pc_0_entry_cfi_idx_valid(core_io_ifu_get_pc_0_entry_cfi_idx_valid),
    .io_ifu_get_pc_0_entry_cfi_idx_bits(core_io_ifu_get_pc_0_entry_cfi_idx_bits),
    .io_ifu_get_pc_0_entry_cfi_taken(core_io_ifu_get_pc_0_entry_cfi_taken),
    .io_ifu_get_pc_0_entry_cfi_mispredicted(core_io_ifu_get_pc_0_entry_cfi_mispredicted),
    .io_ifu_get_pc_0_entry_cfi_type(core_io_ifu_get_pc_0_entry_cfi_type),
    .io_ifu_get_pc_0_entry_br_mask(core_io_ifu_get_pc_0_entry_br_mask),
    .io_ifu_get_pc_0_entry_cfi_is_call(core_io_ifu_get_pc_0_entry_cfi_is_call),
    .io_ifu_get_pc_0_entry_cfi_is_ret(core_io_ifu_get_pc_0_entry_cfi_is_ret),
    .io_ifu_get_pc_0_entry_cfi_npc_plus4(core_io_ifu_get_pc_0_entry_cfi_npc_plus4),
    .io_ifu_get_pc_0_entry_ras_top(core_io_ifu_get_pc_0_entry_ras_top),
    .io_ifu_get_pc_0_entry_ras_idx(core_io_ifu_get_pc_0_entry_ras_idx),
    .io_ifu_get_pc_0_entry_start_bank(core_io_ifu_get_pc_0_entry_start_bank),
    .io_ifu_get_pc_0_ghist_old_history(core_io_ifu_get_pc_0_ghist_old_history),
    .io_ifu_get_pc_0_ghist_current_saw_branch_not_taken(core_io_ifu_get_pc_0_ghist_current_saw_branch_not_taken),
    .io_ifu_get_pc_0_ghist_new_saw_branch_not_taken(core_io_ifu_get_pc_0_ghist_new_saw_branch_not_taken),
    .io_ifu_get_pc_0_ghist_new_saw_branch_taken(core_io_ifu_get_pc_0_ghist_new_saw_branch_taken),
    .io_ifu_get_pc_0_ghist_ras_idx(core_io_ifu_get_pc_0_ghist_ras_idx),
    .io_ifu_get_pc_0_pc(core_io_ifu_get_pc_0_pc),
    .io_ifu_get_pc_0_com_pc(core_io_ifu_get_pc_0_com_pc),
    .io_ifu_get_pc_0_next_val(core_io_ifu_get_pc_0_next_val),
    .io_ifu_get_pc_0_next_pc(core_io_ifu_get_pc_0_next_pc),
    .io_ifu_get_pc_1_ftq_idx(core_io_ifu_get_pc_1_ftq_idx),
    .io_ifu_get_pc_1_entry_cfi_idx_valid(core_io_ifu_get_pc_1_entry_cfi_idx_valid),
    .io_ifu_get_pc_1_entry_cfi_idx_bits(core_io_ifu_get_pc_1_entry_cfi_idx_bits),
    .io_ifu_get_pc_1_entry_cfi_taken(core_io_ifu_get_pc_1_entry_cfi_taken),
    .io_ifu_get_pc_1_entry_cfi_mispredicted(core_io_ifu_get_pc_1_entry_cfi_mispredicted),
    .io_ifu_get_pc_1_entry_cfi_type(core_io_ifu_get_pc_1_entry_cfi_type),
    .io_ifu_get_pc_1_entry_br_mask(core_io_ifu_get_pc_1_entry_br_mask),
    .io_ifu_get_pc_1_entry_cfi_is_call(core_io_ifu_get_pc_1_entry_cfi_is_call),
    .io_ifu_get_pc_1_entry_cfi_is_ret(core_io_ifu_get_pc_1_entry_cfi_is_ret),
    .io_ifu_get_pc_1_entry_cfi_npc_plus4(core_io_ifu_get_pc_1_entry_cfi_npc_plus4),
    .io_ifu_get_pc_1_entry_ras_top(core_io_ifu_get_pc_1_entry_ras_top),
    .io_ifu_get_pc_1_entry_ras_idx(core_io_ifu_get_pc_1_entry_ras_idx),
    .io_ifu_get_pc_1_entry_start_bank(core_io_ifu_get_pc_1_entry_start_bank),
    .io_ifu_get_pc_1_ghist_old_history(core_io_ifu_get_pc_1_ghist_old_history),
    .io_ifu_get_pc_1_ghist_current_saw_branch_not_taken(core_io_ifu_get_pc_1_ghist_current_saw_branch_not_taken),
    .io_ifu_get_pc_1_ghist_new_saw_branch_not_taken(core_io_ifu_get_pc_1_ghist_new_saw_branch_not_taken),
    .io_ifu_get_pc_1_ghist_new_saw_branch_taken(core_io_ifu_get_pc_1_ghist_new_saw_branch_taken),
    .io_ifu_get_pc_1_ghist_ras_idx(core_io_ifu_get_pc_1_ghist_ras_idx),
    .io_ifu_get_pc_1_pc(core_io_ifu_get_pc_1_pc),
    .io_ifu_get_pc_1_com_pc(core_io_ifu_get_pc_1_com_pc),
    .io_ifu_get_pc_1_next_val(core_io_ifu_get_pc_1_next_val),
    .io_ifu_get_pc_1_next_pc(core_io_ifu_get_pc_1_next_pc),
    .io_ifu_get_pc_2_ftq_idx(core_io_ifu_get_pc_2_ftq_idx),
    .io_ifu_get_pc_2_entry_cfi_idx_valid(core_io_ifu_get_pc_2_entry_cfi_idx_valid),
    .io_ifu_get_pc_2_entry_cfi_idx_bits(core_io_ifu_get_pc_2_entry_cfi_idx_bits),
    .io_ifu_get_pc_2_entry_cfi_taken(core_io_ifu_get_pc_2_entry_cfi_taken),
    .io_ifu_get_pc_2_entry_cfi_mispredicted(core_io_ifu_get_pc_2_entry_cfi_mispredicted),
    .io_ifu_get_pc_2_entry_cfi_type(core_io_ifu_get_pc_2_entry_cfi_type),
    .io_ifu_get_pc_2_entry_br_mask(core_io_ifu_get_pc_2_entry_br_mask),
    .io_ifu_get_pc_2_entry_cfi_is_call(core_io_ifu_get_pc_2_entry_cfi_is_call),
    .io_ifu_get_pc_2_entry_cfi_is_ret(core_io_ifu_get_pc_2_entry_cfi_is_ret),
    .io_ifu_get_pc_2_entry_cfi_npc_plus4(core_io_ifu_get_pc_2_entry_cfi_npc_plus4),
    .io_ifu_get_pc_2_entry_ras_top(core_io_ifu_get_pc_2_entry_ras_top),
    .io_ifu_get_pc_2_entry_ras_idx(core_io_ifu_get_pc_2_entry_ras_idx),
    .io_ifu_get_pc_2_entry_start_bank(core_io_ifu_get_pc_2_entry_start_bank),
    .io_ifu_get_pc_2_ghist_old_history(core_io_ifu_get_pc_2_ghist_old_history),
    .io_ifu_get_pc_2_ghist_current_saw_branch_not_taken(core_io_ifu_get_pc_2_ghist_current_saw_branch_not_taken),
    .io_ifu_get_pc_2_ghist_new_saw_branch_not_taken(core_io_ifu_get_pc_2_ghist_new_saw_branch_not_taken),
    .io_ifu_get_pc_2_ghist_new_saw_branch_taken(core_io_ifu_get_pc_2_ghist_new_saw_branch_taken),
    .io_ifu_get_pc_2_ghist_ras_idx(core_io_ifu_get_pc_2_ghist_ras_idx),
    .io_ifu_get_pc_2_pc(core_io_ifu_get_pc_2_pc),
    .io_ifu_get_pc_2_com_pc(core_io_ifu_get_pc_2_com_pc),
    .io_ifu_get_pc_2_next_val(core_io_ifu_get_pc_2_next_val),
    .io_ifu_get_pc_2_next_pc(core_io_ifu_get_pc_2_next_pc),
    .io_ifu_get_pc_3_ftq_idx(core_io_ifu_get_pc_3_ftq_idx),
    .io_ifu_get_pc_3_entry_cfi_idx_valid(core_io_ifu_get_pc_3_entry_cfi_idx_valid),
    .io_ifu_get_pc_3_entry_cfi_idx_bits(core_io_ifu_get_pc_3_entry_cfi_idx_bits),
    .io_ifu_get_pc_3_entry_cfi_taken(core_io_ifu_get_pc_3_entry_cfi_taken),
    .io_ifu_get_pc_3_entry_cfi_mispredicted(core_io_ifu_get_pc_3_entry_cfi_mispredicted),
    .io_ifu_get_pc_3_entry_cfi_type(core_io_ifu_get_pc_3_entry_cfi_type),
    .io_ifu_get_pc_3_entry_br_mask(core_io_ifu_get_pc_3_entry_br_mask),
    .io_ifu_get_pc_3_entry_cfi_is_call(core_io_ifu_get_pc_3_entry_cfi_is_call),
    .io_ifu_get_pc_3_entry_cfi_is_ret(core_io_ifu_get_pc_3_entry_cfi_is_ret),
    .io_ifu_get_pc_3_entry_cfi_npc_plus4(core_io_ifu_get_pc_3_entry_cfi_npc_plus4),
    .io_ifu_get_pc_3_entry_ras_top(core_io_ifu_get_pc_3_entry_ras_top),
    .io_ifu_get_pc_3_entry_ras_idx(core_io_ifu_get_pc_3_entry_ras_idx),
    .io_ifu_get_pc_3_entry_start_bank(core_io_ifu_get_pc_3_entry_start_bank),
    .io_ifu_get_pc_3_ghist_old_history(core_io_ifu_get_pc_3_ghist_old_history),
    .io_ifu_get_pc_3_ghist_current_saw_branch_not_taken(core_io_ifu_get_pc_3_ghist_current_saw_branch_not_taken),
    .io_ifu_get_pc_3_ghist_new_saw_branch_not_taken(core_io_ifu_get_pc_3_ghist_new_saw_branch_not_taken),
    .io_ifu_get_pc_3_ghist_new_saw_branch_taken(core_io_ifu_get_pc_3_ghist_new_saw_branch_taken),
    .io_ifu_get_pc_3_ghist_ras_idx(core_io_ifu_get_pc_3_ghist_ras_idx),
    .io_ifu_get_pc_3_pc(core_io_ifu_get_pc_3_pc),
    .io_ifu_get_pc_3_com_pc(core_io_ifu_get_pc_3_com_pc),
    .io_ifu_get_pc_3_next_val(core_io_ifu_get_pc_3_next_val),
    .io_ifu_get_pc_3_next_pc(core_io_ifu_get_pc_3_next_pc),
    .io_ifu_debug_ftq_idx_0(core_io_ifu_debug_ftq_idx_0),
    .io_ifu_debug_ftq_idx_1(core_io_ifu_debug_ftq_idx_1),
    .io_ifu_debug_fetch_pc_0(core_io_ifu_debug_fetch_pc_0),
    .io_ifu_debug_fetch_pc_1(core_io_ifu_debug_fetch_pc_1),
    .io_ifu_status_debug(core_io_ifu_status_debug),
    .io_ifu_status_cease(core_io_ifu_status_cease),
    .io_ifu_status_wfi(core_io_ifu_status_wfi),
    .io_ifu_status_isa(core_io_ifu_status_isa),
    .io_ifu_status_dprv(core_io_ifu_status_dprv),
    .io_ifu_status_prv(core_io_ifu_status_prv),
    .io_ifu_status_sd(core_io_ifu_status_sd),
    .io_ifu_status_zero2(core_io_ifu_status_zero2),
    .io_ifu_status_sxl(core_io_ifu_status_sxl),
    .io_ifu_status_uxl(core_io_ifu_status_uxl),
    .io_ifu_status_sd_rv32(core_io_ifu_status_sd_rv32),
    .io_ifu_status_zero1(core_io_ifu_status_zero1),
    .io_ifu_status_tsr(core_io_ifu_status_tsr),
    .io_ifu_status_tw(core_io_ifu_status_tw),
    .io_ifu_status_tvm(core_io_ifu_status_tvm),
    .io_ifu_status_mxr(core_io_ifu_status_mxr),
    .io_ifu_status_sum(core_io_ifu_status_sum),
    .io_ifu_status_mprv(core_io_ifu_status_mprv),
    .io_ifu_status_xs(core_io_ifu_status_xs),
    .io_ifu_status_fs(core_io_ifu_status_fs),
    .io_ifu_status_mpp(core_io_ifu_status_mpp),
    .io_ifu_status_vs(core_io_ifu_status_vs),
    .io_ifu_status_spp(core_io_ifu_status_spp),
    .io_ifu_status_mpie(core_io_ifu_status_mpie),
    .io_ifu_status_hpie(core_io_ifu_status_hpie),
    .io_ifu_status_spie(core_io_ifu_status_spie),
    .io_ifu_status_upie(core_io_ifu_status_upie),
    .io_ifu_status_mie(core_io_ifu_status_mie),
    .io_ifu_status_hie(core_io_ifu_status_hie),
    .io_ifu_status_sie(core_io_ifu_status_sie),
    .io_ifu_status_uie(core_io_ifu_status_uie),
    .io_ifu_sfence_valid(core_io_ifu_sfence_valid),
    .io_ifu_sfence_bits_rs1(core_io_ifu_sfence_bits_rs1),
    .io_ifu_sfence_bits_rs2(core_io_ifu_sfence_bits_rs2),
    .io_ifu_sfence_bits_addr(core_io_ifu_sfence_bits_addr),
    .io_ifu_sfence_bits_asid(core_io_ifu_sfence_bits_asid),
    .io_ifu_brupdate_b1_resolve_mask(core_io_ifu_brupdate_b1_resolve_mask),
    .io_ifu_brupdate_b1_mispredict_mask(core_io_ifu_brupdate_b1_mispredict_mask),
    .io_ifu_brupdate_b2_uop_switch(core_io_ifu_brupdate_b2_uop_switch),
    .io_ifu_brupdate_b2_uop_switch_off(core_io_ifu_brupdate_b2_uop_switch_off),
    .io_ifu_brupdate_b2_uop_is_unicore(core_io_ifu_brupdate_b2_uop_is_unicore),
    .io_ifu_brupdate_b2_uop_shift(core_io_ifu_brupdate_b2_uop_shift),
    .io_ifu_brupdate_b2_uop_lrs3_rtype(core_io_ifu_brupdate_b2_uop_lrs3_rtype),
    .io_ifu_brupdate_b2_uop_rflag(core_io_ifu_brupdate_b2_uop_rflag),
    .io_ifu_brupdate_b2_uop_wflag(core_io_ifu_brupdate_b2_uop_wflag),
    .io_ifu_brupdate_b2_uop_prflag(core_io_ifu_brupdate_b2_uop_prflag),
    .io_ifu_brupdate_b2_uop_pwflag(core_io_ifu_brupdate_b2_uop_pwflag),
    .io_ifu_brupdate_b2_uop_pflag_busy(core_io_ifu_brupdate_b2_uop_pflag_busy),
    .io_ifu_brupdate_b2_uop_stale_pflag(core_io_ifu_brupdate_b2_uop_stale_pflag),
    .io_ifu_brupdate_b2_uop_op1_sel(core_io_ifu_brupdate_b2_uop_op1_sel),
    .io_ifu_brupdate_b2_uop_op2_sel(core_io_ifu_brupdate_b2_uop_op2_sel),
    .io_ifu_brupdate_b2_uop_split_num(core_io_ifu_brupdate_b2_uop_split_num),
    .io_ifu_brupdate_b2_uop_self_index(core_io_ifu_brupdate_b2_uop_self_index),
    .io_ifu_brupdate_b2_uop_rob_inst_idx(core_io_ifu_brupdate_b2_uop_rob_inst_idx),
    .io_ifu_brupdate_b2_uop_address_num(core_io_ifu_brupdate_b2_uop_address_num),
    .io_ifu_brupdate_b2_uop_uopc(core_io_ifu_brupdate_b2_uop_uopc),
    .io_ifu_brupdate_b2_uop_inst(core_io_ifu_brupdate_b2_uop_inst),
    .io_ifu_brupdate_b2_uop_debug_inst(core_io_ifu_brupdate_b2_uop_debug_inst),
    .io_ifu_brupdate_b2_uop_is_rvc(core_io_ifu_brupdate_b2_uop_is_rvc),
    .io_ifu_brupdate_b2_uop_debug_pc(core_io_ifu_brupdate_b2_uop_debug_pc),
    .io_ifu_brupdate_b2_uop_iq_type(core_io_ifu_brupdate_b2_uop_iq_type),
    .io_ifu_brupdate_b2_uop_fu_code(core_io_ifu_brupdate_b2_uop_fu_code),
    .io_ifu_brupdate_b2_uop_ctrl_br_type(core_io_ifu_brupdate_b2_uop_ctrl_br_type),
    .io_ifu_brupdate_b2_uop_ctrl_op1_sel(core_io_ifu_brupdate_b2_uop_ctrl_op1_sel),
    .io_ifu_brupdate_b2_uop_ctrl_op2_sel(core_io_ifu_brupdate_b2_uop_ctrl_op2_sel),
    .io_ifu_brupdate_b2_uop_ctrl_imm_sel(core_io_ifu_brupdate_b2_uop_ctrl_imm_sel),
    .io_ifu_brupdate_b2_uop_ctrl_op_fcn(core_io_ifu_brupdate_b2_uop_ctrl_op_fcn),
    .io_ifu_brupdate_b2_uop_ctrl_fcn_dw(core_io_ifu_brupdate_b2_uop_ctrl_fcn_dw),
    .io_ifu_brupdate_b2_uop_ctrl_csr_cmd(core_io_ifu_brupdate_b2_uop_ctrl_csr_cmd),
    .io_ifu_brupdate_b2_uop_ctrl_is_load(core_io_ifu_brupdate_b2_uop_ctrl_is_load),
    .io_ifu_brupdate_b2_uop_ctrl_is_sta(core_io_ifu_brupdate_b2_uop_ctrl_is_sta),
    .io_ifu_brupdate_b2_uop_ctrl_is_std(core_io_ifu_brupdate_b2_uop_ctrl_is_std),
    .io_ifu_brupdate_b2_uop_ctrl_op3_sel(core_io_ifu_brupdate_b2_uop_ctrl_op3_sel),
    .io_ifu_brupdate_b2_uop_iw_state(core_io_ifu_brupdate_b2_uop_iw_state),
    .io_ifu_brupdate_b2_uop_iw_p1_poisoned(core_io_ifu_brupdate_b2_uop_iw_p1_poisoned),
    .io_ifu_brupdate_b2_uop_iw_p2_poisoned(core_io_ifu_brupdate_b2_uop_iw_p2_poisoned),
    .io_ifu_brupdate_b2_uop_is_br(core_io_ifu_brupdate_b2_uop_is_br),
    .io_ifu_brupdate_b2_uop_is_jalr(core_io_ifu_brupdate_b2_uop_is_jalr),
    .io_ifu_brupdate_b2_uop_is_jal(core_io_ifu_brupdate_b2_uop_is_jal),
    .io_ifu_brupdate_b2_uop_is_sfb(core_io_ifu_brupdate_b2_uop_is_sfb),
    .io_ifu_brupdate_b2_uop_br_mask(core_io_ifu_brupdate_b2_uop_br_mask),
    .io_ifu_brupdate_b2_uop_br_tag(core_io_ifu_brupdate_b2_uop_br_tag),
    .io_ifu_brupdate_b2_uop_ftq_idx(core_io_ifu_brupdate_b2_uop_ftq_idx),
    .io_ifu_brupdate_b2_uop_edge_inst(core_io_ifu_brupdate_b2_uop_edge_inst),
    .io_ifu_brupdate_b2_uop_pc_lob(core_io_ifu_brupdate_b2_uop_pc_lob),
    .io_ifu_brupdate_b2_uop_taken(core_io_ifu_brupdate_b2_uop_taken),
    .io_ifu_brupdate_b2_uop_imm_packed(core_io_ifu_brupdate_b2_uop_imm_packed),
    .io_ifu_brupdate_b2_uop_csr_addr(core_io_ifu_brupdate_b2_uop_csr_addr),
    .io_ifu_brupdate_b2_uop_rob_idx(core_io_ifu_brupdate_b2_uop_rob_idx),
    .io_ifu_brupdate_b2_uop_ldq_idx(core_io_ifu_brupdate_b2_uop_ldq_idx),
    .io_ifu_brupdate_b2_uop_stq_idx(core_io_ifu_brupdate_b2_uop_stq_idx),
    .io_ifu_brupdate_b2_uop_rxq_idx(core_io_ifu_brupdate_b2_uop_rxq_idx),
    .io_ifu_brupdate_b2_uop_pdst(core_io_ifu_brupdate_b2_uop_pdst),
    .io_ifu_brupdate_b2_uop_prs1(core_io_ifu_brupdate_b2_uop_prs1),
    .io_ifu_brupdate_b2_uop_prs2(core_io_ifu_brupdate_b2_uop_prs2),
    .io_ifu_brupdate_b2_uop_prs3(core_io_ifu_brupdate_b2_uop_prs3),
    .io_ifu_brupdate_b2_uop_ppred(core_io_ifu_brupdate_b2_uop_ppred),
    .io_ifu_brupdate_b2_uop_prs1_busy(core_io_ifu_brupdate_b2_uop_prs1_busy),
    .io_ifu_brupdate_b2_uop_prs2_busy(core_io_ifu_brupdate_b2_uop_prs2_busy),
    .io_ifu_brupdate_b2_uop_prs3_busy(core_io_ifu_brupdate_b2_uop_prs3_busy),
    .io_ifu_brupdate_b2_uop_ppred_busy(core_io_ifu_brupdate_b2_uop_ppred_busy),
    .io_ifu_brupdate_b2_uop_stale_pdst(core_io_ifu_brupdate_b2_uop_stale_pdst),
    .io_ifu_brupdate_b2_uop_exception(core_io_ifu_brupdate_b2_uop_exception),
    .io_ifu_brupdate_b2_uop_exc_cause(core_io_ifu_brupdate_b2_uop_exc_cause),
    .io_ifu_brupdate_b2_uop_bypassable(core_io_ifu_brupdate_b2_uop_bypassable),
    .io_ifu_brupdate_b2_uop_mem_cmd(core_io_ifu_brupdate_b2_uop_mem_cmd),
    .io_ifu_brupdate_b2_uop_mem_size(core_io_ifu_brupdate_b2_uop_mem_size),
    .io_ifu_brupdate_b2_uop_mem_signed(core_io_ifu_brupdate_b2_uop_mem_signed),
    .io_ifu_brupdate_b2_uop_is_fence(core_io_ifu_brupdate_b2_uop_is_fence),
    .io_ifu_brupdate_b2_uop_is_fencei(core_io_ifu_brupdate_b2_uop_is_fencei),
    .io_ifu_brupdate_b2_uop_is_amo(core_io_ifu_brupdate_b2_uop_is_amo),
    .io_ifu_brupdate_b2_uop_uses_ldq(core_io_ifu_brupdate_b2_uop_uses_ldq),
    .io_ifu_brupdate_b2_uop_uses_stq(core_io_ifu_brupdate_b2_uop_uses_stq),
    .io_ifu_brupdate_b2_uop_is_sys_pc2epc(core_io_ifu_brupdate_b2_uop_is_sys_pc2epc),
    .io_ifu_brupdate_b2_uop_is_unique(core_io_ifu_brupdate_b2_uop_is_unique),
    .io_ifu_brupdate_b2_uop_flush_on_commit(core_io_ifu_brupdate_b2_uop_flush_on_commit),
    .io_ifu_brupdate_b2_uop_ldst_is_rs1(core_io_ifu_brupdate_b2_uop_ldst_is_rs1),
    .io_ifu_brupdate_b2_uop_ldst(core_io_ifu_brupdate_b2_uop_ldst),
    .io_ifu_brupdate_b2_uop_lrs1(core_io_ifu_brupdate_b2_uop_lrs1),
    .io_ifu_brupdate_b2_uop_lrs2(core_io_ifu_brupdate_b2_uop_lrs2),
    .io_ifu_brupdate_b2_uop_lrs3(core_io_ifu_brupdate_b2_uop_lrs3),
    .io_ifu_brupdate_b2_uop_ldst_val(core_io_ifu_brupdate_b2_uop_ldst_val),
    .io_ifu_brupdate_b2_uop_dst_rtype(core_io_ifu_brupdate_b2_uop_dst_rtype),
    .io_ifu_brupdate_b2_uop_lrs1_rtype(core_io_ifu_brupdate_b2_uop_lrs1_rtype),
    .io_ifu_brupdate_b2_uop_lrs2_rtype(core_io_ifu_brupdate_b2_uop_lrs2_rtype),
    .io_ifu_brupdate_b2_uop_frs3_en(core_io_ifu_brupdate_b2_uop_frs3_en),
    .io_ifu_brupdate_b2_uop_fp_val(core_io_ifu_brupdate_b2_uop_fp_val),
    .io_ifu_brupdate_b2_uop_fp_single(core_io_ifu_brupdate_b2_uop_fp_single),
    .io_ifu_brupdate_b2_uop_xcpt_pf_if(core_io_ifu_brupdate_b2_uop_xcpt_pf_if),
    .io_ifu_brupdate_b2_uop_xcpt_ae_if(core_io_ifu_brupdate_b2_uop_xcpt_ae_if),
    .io_ifu_brupdate_b2_uop_xcpt_ma_if(core_io_ifu_brupdate_b2_uop_xcpt_ma_if),
    .io_ifu_brupdate_b2_uop_bp_debug_if(core_io_ifu_brupdate_b2_uop_bp_debug_if),
    .io_ifu_brupdate_b2_uop_bp_xcpt_if(core_io_ifu_brupdate_b2_uop_bp_xcpt_if),
    .io_ifu_brupdate_b2_uop_debug_fsrc(core_io_ifu_brupdate_b2_uop_debug_fsrc),
    .io_ifu_brupdate_b2_uop_debug_tsrc(core_io_ifu_brupdate_b2_uop_debug_tsrc),
    .io_ifu_brupdate_b2_valid(core_io_ifu_brupdate_b2_valid),
    .io_ifu_brupdate_b2_mispredict(core_io_ifu_brupdate_b2_mispredict),
    .io_ifu_brupdate_b2_taken(core_io_ifu_brupdate_b2_taken),
    .io_ifu_brupdate_b2_cfi_type(core_io_ifu_brupdate_b2_cfi_type),
    .io_ifu_brupdate_b2_pc_sel(core_io_ifu_brupdate_b2_pc_sel),
    .io_ifu_brupdate_b2_jalr_target(core_io_ifu_brupdate_b2_jalr_target),
    .io_ifu_brupdate_b2_target_offset(core_io_ifu_brupdate_b2_target_offset),
    .io_ifu_redirect_flush(core_io_ifu_redirect_flush),
    .io_ifu_redirect_val(core_io_ifu_redirect_val),
    .io_ifu_redirect_pc(core_io_ifu_redirect_pc),
    .io_ifu_redirect_ftq_idx(core_io_ifu_redirect_ftq_idx),
    .io_ifu_redirect_ghist_old_history(core_io_ifu_redirect_ghist_old_history),
    .io_ifu_redirect_ghist_current_saw_branch_not_taken(core_io_ifu_redirect_ghist_current_saw_branch_not_taken),
    .io_ifu_redirect_ghist_new_saw_branch_not_taken(core_io_ifu_redirect_ghist_new_saw_branch_not_taken),
    .io_ifu_redirect_ghist_new_saw_branch_taken(core_io_ifu_redirect_ghist_new_saw_branch_taken),
    .io_ifu_redirect_ghist_ras_idx(core_io_ifu_redirect_ghist_ras_idx),
    .io_ifu_commit_valid(core_io_ifu_commit_valid),
    .io_ifu_commit_bits(core_io_ifu_commit_bits),
    .io_ifu_flush_icache(core_io_ifu_flush_icache),
    .io_ifu_perf_acquire(core_io_ifu_perf_acquire),
    .io_ifu_perf_tlbMiss(core_io_ifu_perf_tlbMiss),
    .io_ifu_is_unicore(core_io_ifu_is_unicore),
    .io_ptw_ptbr_mode(core_io_ptw_ptbr_mode),
    .io_ptw_ptbr_asid(core_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(core_io_ptw_ptbr_ppn),
    .io_ptw_sfence_valid(core_io_ptw_sfence_valid),
    .io_ptw_sfence_bits_rs1(core_io_ptw_sfence_bits_rs1),
    .io_ptw_sfence_bits_rs2(core_io_ptw_sfence_bits_rs2),
    .io_ptw_sfence_bits_addr(core_io_ptw_sfence_bits_addr),
    .io_ptw_sfence_bits_asid(core_io_ptw_sfence_bits_asid),
    .io_ptw_status_debug(core_io_ptw_status_debug),
    .io_ptw_status_cease(core_io_ptw_status_cease),
    .io_ptw_status_wfi(core_io_ptw_status_wfi),
    .io_ptw_status_isa(core_io_ptw_status_isa),
    .io_ptw_status_dprv(core_io_ptw_status_dprv),
    .io_ptw_status_prv(core_io_ptw_status_prv),
    .io_ptw_status_sd(core_io_ptw_status_sd),
    .io_ptw_status_zero2(core_io_ptw_status_zero2),
    .io_ptw_status_sxl(core_io_ptw_status_sxl),
    .io_ptw_status_uxl(core_io_ptw_status_uxl),
    .io_ptw_status_sd_rv32(core_io_ptw_status_sd_rv32),
    .io_ptw_status_zero1(core_io_ptw_status_zero1),
    .io_ptw_status_tsr(core_io_ptw_status_tsr),
    .io_ptw_status_tw(core_io_ptw_status_tw),
    .io_ptw_status_tvm(core_io_ptw_status_tvm),
    .io_ptw_status_mxr(core_io_ptw_status_mxr),
    .io_ptw_status_sum(core_io_ptw_status_sum),
    .io_ptw_status_mprv(core_io_ptw_status_mprv),
    .io_ptw_status_xs(core_io_ptw_status_xs),
    .io_ptw_status_fs(core_io_ptw_status_fs),
    .io_ptw_status_mpp(core_io_ptw_status_mpp),
    .io_ptw_status_vs(core_io_ptw_status_vs),
    .io_ptw_status_spp(core_io_ptw_status_spp),
    .io_ptw_status_mpie(core_io_ptw_status_mpie),
    .io_ptw_status_hpie(core_io_ptw_status_hpie),
    .io_ptw_status_spie(core_io_ptw_status_spie),
    .io_ptw_status_upie(core_io_ptw_status_upie),
    .io_ptw_status_mie(core_io_ptw_status_mie),
    .io_ptw_status_hie(core_io_ptw_status_hie),
    .io_ptw_status_sie(core_io_ptw_status_sie),
    .io_ptw_status_uie(core_io_ptw_status_uie),
    .io_ptw_pmp_0_cfg_l(core_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_res(core_io_ptw_pmp_0_cfg_res),
    .io_ptw_pmp_0_cfg_a(core_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(core_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(core_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(core_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(core_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(core_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(core_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_res(core_io_ptw_pmp_1_cfg_res),
    .io_ptw_pmp_1_cfg_a(core_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(core_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(core_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(core_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(core_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(core_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(core_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_res(core_io_ptw_pmp_2_cfg_res),
    .io_ptw_pmp_2_cfg_a(core_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(core_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(core_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(core_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(core_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(core_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(core_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_res(core_io_ptw_pmp_3_cfg_res),
    .io_ptw_pmp_3_cfg_a(core_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(core_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(core_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(core_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(core_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(core_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(core_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_res(core_io_ptw_pmp_4_cfg_res),
    .io_ptw_pmp_4_cfg_a(core_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(core_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(core_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(core_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(core_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(core_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(core_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_res(core_io_ptw_pmp_5_cfg_res),
    .io_ptw_pmp_5_cfg_a(core_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(core_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(core_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(core_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(core_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(core_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(core_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_res(core_io_ptw_pmp_6_cfg_res),
    .io_ptw_pmp_6_cfg_a(core_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(core_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(core_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(core_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(core_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(core_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(core_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_res(core_io_ptw_pmp_7_cfg_res),
    .io_ptw_pmp_7_cfg_a(core_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(core_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(core_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(core_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(core_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(core_io_ptw_pmp_7_mask),
    .io_ptw_perf_l2miss(core_io_ptw_perf_l2miss),
    .io_ptw_perf_l2hit(core_io_ptw_perf_l2hit),
    .io_ptw_perf_pte_miss(core_io_ptw_perf_pte_miss),
    .io_ptw_perf_pte_hit(core_io_ptw_perf_pte_hit),
    .io_ptw_customCSRs_csrs_0_wen(core_io_ptw_customCSRs_csrs_0_wen),
    .io_ptw_customCSRs_csrs_0_wdata(core_io_ptw_customCSRs_csrs_0_wdata),
    .io_ptw_customCSRs_csrs_0_value(core_io_ptw_customCSRs_csrs_0_value),
    .io_ptw_clock_enabled(core_io_ptw_clock_enabled),
    .io_rocc_cmd_ready(core_io_rocc_cmd_ready),
    .io_rocc_cmd_valid(core_io_rocc_cmd_valid),
    .io_rocc_cmd_bits_inst_funct(core_io_rocc_cmd_bits_inst_funct),
    .io_rocc_cmd_bits_inst_rs2(core_io_rocc_cmd_bits_inst_rs2),
    .io_rocc_cmd_bits_inst_rs1(core_io_rocc_cmd_bits_inst_rs1),
    .io_rocc_cmd_bits_inst_xd(core_io_rocc_cmd_bits_inst_xd),
    .io_rocc_cmd_bits_inst_xs1(core_io_rocc_cmd_bits_inst_xs1),
    .io_rocc_cmd_bits_inst_xs2(core_io_rocc_cmd_bits_inst_xs2),
    .io_rocc_cmd_bits_inst_rd(core_io_rocc_cmd_bits_inst_rd),
    .io_rocc_cmd_bits_inst_opcode(core_io_rocc_cmd_bits_inst_opcode),
    .io_rocc_cmd_bits_rs1(core_io_rocc_cmd_bits_rs1),
    .io_rocc_cmd_bits_rs2(core_io_rocc_cmd_bits_rs2),
    .io_rocc_cmd_bits_status_debug(core_io_rocc_cmd_bits_status_debug),
    .io_rocc_cmd_bits_status_cease(core_io_rocc_cmd_bits_status_cease),
    .io_rocc_cmd_bits_status_wfi(core_io_rocc_cmd_bits_status_wfi),
    .io_rocc_cmd_bits_status_isa(core_io_rocc_cmd_bits_status_isa),
    .io_rocc_cmd_bits_status_dprv(core_io_rocc_cmd_bits_status_dprv),
    .io_rocc_cmd_bits_status_prv(core_io_rocc_cmd_bits_status_prv),
    .io_rocc_cmd_bits_status_sd(core_io_rocc_cmd_bits_status_sd),
    .io_rocc_cmd_bits_status_zero2(core_io_rocc_cmd_bits_status_zero2),
    .io_rocc_cmd_bits_status_sxl(core_io_rocc_cmd_bits_status_sxl),
    .io_rocc_cmd_bits_status_uxl(core_io_rocc_cmd_bits_status_uxl),
    .io_rocc_cmd_bits_status_sd_rv32(core_io_rocc_cmd_bits_status_sd_rv32),
    .io_rocc_cmd_bits_status_zero1(core_io_rocc_cmd_bits_status_zero1),
    .io_rocc_cmd_bits_status_tsr(core_io_rocc_cmd_bits_status_tsr),
    .io_rocc_cmd_bits_status_tw(core_io_rocc_cmd_bits_status_tw),
    .io_rocc_cmd_bits_status_tvm(core_io_rocc_cmd_bits_status_tvm),
    .io_rocc_cmd_bits_status_mxr(core_io_rocc_cmd_bits_status_mxr),
    .io_rocc_cmd_bits_status_sum(core_io_rocc_cmd_bits_status_sum),
    .io_rocc_cmd_bits_status_mprv(core_io_rocc_cmd_bits_status_mprv),
    .io_rocc_cmd_bits_status_xs(core_io_rocc_cmd_bits_status_xs),
    .io_rocc_cmd_bits_status_fs(core_io_rocc_cmd_bits_status_fs),
    .io_rocc_cmd_bits_status_mpp(core_io_rocc_cmd_bits_status_mpp),
    .io_rocc_cmd_bits_status_vs(core_io_rocc_cmd_bits_status_vs),
    .io_rocc_cmd_bits_status_spp(core_io_rocc_cmd_bits_status_spp),
    .io_rocc_cmd_bits_status_mpie(core_io_rocc_cmd_bits_status_mpie),
    .io_rocc_cmd_bits_status_hpie(core_io_rocc_cmd_bits_status_hpie),
    .io_rocc_cmd_bits_status_spie(core_io_rocc_cmd_bits_status_spie),
    .io_rocc_cmd_bits_status_upie(core_io_rocc_cmd_bits_status_upie),
    .io_rocc_cmd_bits_status_mie(core_io_rocc_cmd_bits_status_mie),
    .io_rocc_cmd_bits_status_hie(core_io_rocc_cmd_bits_status_hie),
    .io_rocc_cmd_bits_status_sie(core_io_rocc_cmd_bits_status_sie),
    .io_rocc_cmd_bits_status_uie(core_io_rocc_cmd_bits_status_uie),
    .io_rocc_resp_ready(core_io_rocc_resp_ready),
    .io_rocc_resp_valid(core_io_rocc_resp_valid),
    .io_rocc_resp_bits_rd(core_io_rocc_resp_bits_rd),
    .io_rocc_resp_bits_data(core_io_rocc_resp_bits_data),
    .io_rocc_mem_req_ready(core_io_rocc_mem_req_ready),
    .io_rocc_mem_req_valid(core_io_rocc_mem_req_valid),
    .io_rocc_mem_req_bits_addr(core_io_rocc_mem_req_bits_addr),
    .io_rocc_mem_req_bits_tag(core_io_rocc_mem_req_bits_tag),
    .io_rocc_mem_req_bits_cmd(core_io_rocc_mem_req_bits_cmd),
    .io_rocc_mem_req_bits_size(core_io_rocc_mem_req_bits_size),
    .io_rocc_mem_req_bits_signed(core_io_rocc_mem_req_bits_signed),
    .io_rocc_mem_req_bits_dprv(core_io_rocc_mem_req_bits_dprv),
    .io_rocc_mem_req_bits_phys(core_io_rocc_mem_req_bits_phys),
    .io_rocc_mem_req_bits_no_alloc(core_io_rocc_mem_req_bits_no_alloc),
    .io_rocc_mem_req_bits_no_xcpt(core_io_rocc_mem_req_bits_no_xcpt),
    .io_rocc_mem_req_bits_data(core_io_rocc_mem_req_bits_data),
    .io_rocc_mem_req_bits_mask(core_io_rocc_mem_req_bits_mask),
    .io_rocc_mem_s1_kill(core_io_rocc_mem_s1_kill),
    .io_rocc_mem_s1_data_data(core_io_rocc_mem_s1_data_data),
    .io_rocc_mem_s1_data_mask(core_io_rocc_mem_s1_data_mask),
    .io_rocc_mem_s2_nack(core_io_rocc_mem_s2_nack),
    .io_rocc_mem_s2_nack_cause_raw(core_io_rocc_mem_s2_nack_cause_raw),
    .io_rocc_mem_s2_kill(core_io_rocc_mem_s2_kill),
    .io_rocc_mem_s2_uncached(core_io_rocc_mem_s2_uncached),
    .io_rocc_mem_s2_paddr(core_io_rocc_mem_s2_paddr),
    .io_rocc_mem_resp_valid(core_io_rocc_mem_resp_valid),
    .io_rocc_mem_resp_bits_addr(core_io_rocc_mem_resp_bits_addr),
    .io_rocc_mem_resp_bits_tag(core_io_rocc_mem_resp_bits_tag),
    .io_rocc_mem_resp_bits_cmd(core_io_rocc_mem_resp_bits_cmd),
    .io_rocc_mem_resp_bits_size(core_io_rocc_mem_resp_bits_size),
    .io_rocc_mem_resp_bits_signed(core_io_rocc_mem_resp_bits_signed),
    .io_rocc_mem_resp_bits_dprv(core_io_rocc_mem_resp_bits_dprv),
    .io_rocc_mem_resp_bits_data(core_io_rocc_mem_resp_bits_data),
    .io_rocc_mem_resp_bits_mask(core_io_rocc_mem_resp_bits_mask),
    .io_rocc_mem_resp_bits_replay(core_io_rocc_mem_resp_bits_replay),
    .io_rocc_mem_resp_bits_has_data(core_io_rocc_mem_resp_bits_has_data),
    .io_rocc_mem_resp_bits_data_word_bypass(core_io_rocc_mem_resp_bits_data_word_bypass),
    .io_rocc_mem_resp_bits_data_raw(core_io_rocc_mem_resp_bits_data_raw),
    .io_rocc_mem_resp_bits_store_data(core_io_rocc_mem_resp_bits_store_data),
    .io_rocc_mem_replay_next(core_io_rocc_mem_replay_next),
    .io_rocc_mem_s2_xcpt_ma_ld(core_io_rocc_mem_s2_xcpt_ma_ld),
    .io_rocc_mem_s2_xcpt_ma_st(core_io_rocc_mem_s2_xcpt_ma_st),
    .io_rocc_mem_s2_xcpt_pf_ld(core_io_rocc_mem_s2_xcpt_pf_ld),
    .io_rocc_mem_s2_xcpt_pf_st(core_io_rocc_mem_s2_xcpt_pf_st),
    .io_rocc_mem_s2_xcpt_ae_ld(core_io_rocc_mem_s2_xcpt_ae_ld),
    .io_rocc_mem_s2_xcpt_ae_st(core_io_rocc_mem_s2_xcpt_ae_st),
    .io_rocc_mem_ordered(core_io_rocc_mem_ordered),
    .io_rocc_mem_perf_acquire(core_io_rocc_mem_perf_acquire),
    .io_rocc_mem_perf_release(core_io_rocc_mem_perf_release),
    .io_rocc_mem_perf_grant(core_io_rocc_mem_perf_grant),
    .io_rocc_mem_perf_tlbMiss(core_io_rocc_mem_perf_tlbMiss),
    .io_rocc_mem_perf_blocked(core_io_rocc_mem_perf_blocked),
    .io_rocc_mem_perf_canAcceptStoreThenLoad(core_io_rocc_mem_perf_canAcceptStoreThenLoad),
    .io_rocc_mem_perf_canAcceptStoreThenRMW(core_io_rocc_mem_perf_canAcceptStoreThenRMW),
    .io_rocc_mem_perf_canAcceptLoadThenLoad(core_io_rocc_mem_perf_canAcceptLoadThenLoad),
    .io_rocc_mem_perf_storeBufferEmptyAfterLoad(core_io_rocc_mem_perf_storeBufferEmptyAfterLoad),
    .io_rocc_mem_perf_storeBufferEmptyAfterStore(core_io_rocc_mem_perf_storeBufferEmptyAfterStore),
    .io_rocc_mem_keep_clock_enabled(core_io_rocc_mem_keep_clock_enabled),
    .io_rocc_mem_clock_enabled(core_io_rocc_mem_clock_enabled),
    .io_rocc_busy(core_io_rocc_busy),
    .io_rocc_interrupt(core_io_rocc_interrupt),
    .io_rocc_exception(core_io_rocc_exception),
    .io_lsu_exe_0_req_valid(core_io_lsu_exe_0_req_valid),
    .io_lsu_exe_0_req_bits_uop_switch(core_io_lsu_exe_0_req_bits_uop_switch),
    .io_lsu_exe_0_req_bits_uop_switch_off(core_io_lsu_exe_0_req_bits_uop_switch_off),
    .io_lsu_exe_0_req_bits_uop_is_unicore(core_io_lsu_exe_0_req_bits_uop_is_unicore),
    .io_lsu_exe_0_req_bits_uop_shift(core_io_lsu_exe_0_req_bits_uop_shift),
    .io_lsu_exe_0_req_bits_uop_lrs3_rtype(core_io_lsu_exe_0_req_bits_uop_lrs3_rtype),
    .io_lsu_exe_0_req_bits_uop_rflag(core_io_lsu_exe_0_req_bits_uop_rflag),
    .io_lsu_exe_0_req_bits_uop_wflag(core_io_lsu_exe_0_req_bits_uop_wflag),
    .io_lsu_exe_0_req_bits_uop_prflag(core_io_lsu_exe_0_req_bits_uop_prflag),
    .io_lsu_exe_0_req_bits_uop_pwflag(core_io_lsu_exe_0_req_bits_uop_pwflag),
    .io_lsu_exe_0_req_bits_uop_pflag_busy(core_io_lsu_exe_0_req_bits_uop_pflag_busy),
    .io_lsu_exe_0_req_bits_uop_stale_pflag(core_io_lsu_exe_0_req_bits_uop_stale_pflag),
    .io_lsu_exe_0_req_bits_uop_op1_sel(core_io_lsu_exe_0_req_bits_uop_op1_sel),
    .io_lsu_exe_0_req_bits_uop_op2_sel(core_io_lsu_exe_0_req_bits_uop_op2_sel),
    .io_lsu_exe_0_req_bits_uop_split_num(core_io_lsu_exe_0_req_bits_uop_split_num),
    .io_lsu_exe_0_req_bits_uop_self_index(core_io_lsu_exe_0_req_bits_uop_self_index),
    .io_lsu_exe_0_req_bits_uop_rob_inst_idx(core_io_lsu_exe_0_req_bits_uop_rob_inst_idx),
    .io_lsu_exe_0_req_bits_uop_address_num(core_io_lsu_exe_0_req_bits_uop_address_num),
    .io_lsu_exe_0_req_bits_uop_uopc(core_io_lsu_exe_0_req_bits_uop_uopc),
    .io_lsu_exe_0_req_bits_uop_inst(core_io_lsu_exe_0_req_bits_uop_inst),
    .io_lsu_exe_0_req_bits_uop_debug_inst(core_io_lsu_exe_0_req_bits_uop_debug_inst),
    .io_lsu_exe_0_req_bits_uop_is_rvc(core_io_lsu_exe_0_req_bits_uop_is_rvc),
    .io_lsu_exe_0_req_bits_uop_debug_pc(core_io_lsu_exe_0_req_bits_uop_debug_pc),
    .io_lsu_exe_0_req_bits_uop_iq_type(core_io_lsu_exe_0_req_bits_uop_iq_type),
    .io_lsu_exe_0_req_bits_uop_fu_code(core_io_lsu_exe_0_req_bits_uop_fu_code),
    .io_lsu_exe_0_req_bits_uop_ctrl_br_type(core_io_lsu_exe_0_req_bits_uop_ctrl_br_type),
    .io_lsu_exe_0_req_bits_uop_ctrl_op1_sel(core_io_lsu_exe_0_req_bits_uop_ctrl_op1_sel),
    .io_lsu_exe_0_req_bits_uop_ctrl_op2_sel(core_io_lsu_exe_0_req_bits_uop_ctrl_op2_sel),
    .io_lsu_exe_0_req_bits_uop_ctrl_imm_sel(core_io_lsu_exe_0_req_bits_uop_ctrl_imm_sel),
    .io_lsu_exe_0_req_bits_uop_ctrl_op_fcn(core_io_lsu_exe_0_req_bits_uop_ctrl_op_fcn),
    .io_lsu_exe_0_req_bits_uop_ctrl_fcn_dw(core_io_lsu_exe_0_req_bits_uop_ctrl_fcn_dw),
    .io_lsu_exe_0_req_bits_uop_ctrl_csr_cmd(core_io_lsu_exe_0_req_bits_uop_ctrl_csr_cmd),
    .io_lsu_exe_0_req_bits_uop_ctrl_is_load(core_io_lsu_exe_0_req_bits_uop_ctrl_is_load),
    .io_lsu_exe_0_req_bits_uop_ctrl_is_sta(core_io_lsu_exe_0_req_bits_uop_ctrl_is_sta),
    .io_lsu_exe_0_req_bits_uop_ctrl_is_std(core_io_lsu_exe_0_req_bits_uop_ctrl_is_std),
    .io_lsu_exe_0_req_bits_uop_ctrl_op3_sel(core_io_lsu_exe_0_req_bits_uop_ctrl_op3_sel),
    .io_lsu_exe_0_req_bits_uop_iw_state(core_io_lsu_exe_0_req_bits_uop_iw_state),
    .io_lsu_exe_0_req_bits_uop_iw_p1_poisoned(core_io_lsu_exe_0_req_bits_uop_iw_p1_poisoned),
    .io_lsu_exe_0_req_bits_uop_iw_p2_poisoned(core_io_lsu_exe_0_req_bits_uop_iw_p2_poisoned),
    .io_lsu_exe_0_req_bits_uop_is_br(core_io_lsu_exe_0_req_bits_uop_is_br),
    .io_lsu_exe_0_req_bits_uop_is_jalr(core_io_lsu_exe_0_req_bits_uop_is_jalr),
    .io_lsu_exe_0_req_bits_uop_is_jal(core_io_lsu_exe_0_req_bits_uop_is_jal),
    .io_lsu_exe_0_req_bits_uop_is_sfb(core_io_lsu_exe_0_req_bits_uop_is_sfb),
    .io_lsu_exe_0_req_bits_uop_br_mask(core_io_lsu_exe_0_req_bits_uop_br_mask),
    .io_lsu_exe_0_req_bits_uop_br_tag(core_io_lsu_exe_0_req_bits_uop_br_tag),
    .io_lsu_exe_0_req_bits_uop_ftq_idx(core_io_lsu_exe_0_req_bits_uop_ftq_idx),
    .io_lsu_exe_0_req_bits_uop_edge_inst(core_io_lsu_exe_0_req_bits_uop_edge_inst),
    .io_lsu_exe_0_req_bits_uop_pc_lob(core_io_lsu_exe_0_req_bits_uop_pc_lob),
    .io_lsu_exe_0_req_bits_uop_taken(core_io_lsu_exe_0_req_bits_uop_taken),
    .io_lsu_exe_0_req_bits_uop_imm_packed(core_io_lsu_exe_0_req_bits_uop_imm_packed),
    .io_lsu_exe_0_req_bits_uop_csr_addr(core_io_lsu_exe_0_req_bits_uop_csr_addr),
    .io_lsu_exe_0_req_bits_uop_rob_idx(core_io_lsu_exe_0_req_bits_uop_rob_idx),
    .io_lsu_exe_0_req_bits_uop_ldq_idx(core_io_lsu_exe_0_req_bits_uop_ldq_idx),
    .io_lsu_exe_0_req_bits_uop_stq_idx(core_io_lsu_exe_0_req_bits_uop_stq_idx),
    .io_lsu_exe_0_req_bits_uop_rxq_idx(core_io_lsu_exe_0_req_bits_uop_rxq_idx),
    .io_lsu_exe_0_req_bits_uop_pdst(core_io_lsu_exe_0_req_bits_uop_pdst),
    .io_lsu_exe_0_req_bits_uop_prs1(core_io_lsu_exe_0_req_bits_uop_prs1),
    .io_lsu_exe_0_req_bits_uop_prs2(core_io_lsu_exe_0_req_bits_uop_prs2),
    .io_lsu_exe_0_req_bits_uop_prs3(core_io_lsu_exe_0_req_bits_uop_prs3),
    .io_lsu_exe_0_req_bits_uop_ppred(core_io_lsu_exe_0_req_bits_uop_ppred),
    .io_lsu_exe_0_req_bits_uop_prs1_busy(core_io_lsu_exe_0_req_bits_uop_prs1_busy),
    .io_lsu_exe_0_req_bits_uop_prs2_busy(core_io_lsu_exe_0_req_bits_uop_prs2_busy),
    .io_lsu_exe_0_req_bits_uop_prs3_busy(core_io_lsu_exe_0_req_bits_uop_prs3_busy),
    .io_lsu_exe_0_req_bits_uop_ppred_busy(core_io_lsu_exe_0_req_bits_uop_ppred_busy),
    .io_lsu_exe_0_req_bits_uop_stale_pdst(core_io_lsu_exe_0_req_bits_uop_stale_pdst),
    .io_lsu_exe_0_req_bits_uop_exception(core_io_lsu_exe_0_req_bits_uop_exception),
    .io_lsu_exe_0_req_bits_uop_exc_cause(core_io_lsu_exe_0_req_bits_uop_exc_cause),
    .io_lsu_exe_0_req_bits_uop_bypassable(core_io_lsu_exe_0_req_bits_uop_bypassable),
    .io_lsu_exe_0_req_bits_uop_mem_cmd(core_io_lsu_exe_0_req_bits_uop_mem_cmd),
    .io_lsu_exe_0_req_bits_uop_mem_size(core_io_lsu_exe_0_req_bits_uop_mem_size),
    .io_lsu_exe_0_req_bits_uop_mem_signed(core_io_lsu_exe_0_req_bits_uop_mem_signed),
    .io_lsu_exe_0_req_bits_uop_is_fence(core_io_lsu_exe_0_req_bits_uop_is_fence),
    .io_lsu_exe_0_req_bits_uop_is_fencei(core_io_lsu_exe_0_req_bits_uop_is_fencei),
    .io_lsu_exe_0_req_bits_uop_is_amo(core_io_lsu_exe_0_req_bits_uop_is_amo),
    .io_lsu_exe_0_req_bits_uop_uses_ldq(core_io_lsu_exe_0_req_bits_uop_uses_ldq),
    .io_lsu_exe_0_req_bits_uop_uses_stq(core_io_lsu_exe_0_req_bits_uop_uses_stq),
    .io_lsu_exe_0_req_bits_uop_is_sys_pc2epc(core_io_lsu_exe_0_req_bits_uop_is_sys_pc2epc),
    .io_lsu_exe_0_req_bits_uop_is_unique(core_io_lsu_exe_0_req_bits_uop_is_unique),
    .io_lsu_exe_0_req_bits_uop_flush_on_commit(core_io_lsu_exe_0_req_bits_uop_flush_on_commit),
    .io_lsu_exe_0_req_bits_uop_ldst_is_rs1(core_io_lsu_exe_0_req_bits_uop_ldst_is_rs1),
    .io_lsu_exe_0_req_bits_uop_ldst(core_io_lsu_exe_0_req_bits_uop_ldst),
    .io_lsu_exe_0_req_bits_uop_lrs1(core_io_lsu_exe_0_req_bits_uop_lrs1),
    .io_lsu_exe_0_req_bits_uop_lrs2(core_io_lsu_exe_0_req_bits_uop_lrs2),
    .io_lsu_exe_0_req_bits_uop_lrs3(core_io_lsu_exe_0_req_bits_uop_lrs3),
    .io_lsu_exe_0_req_bits_uop_ldst_val(core_io_lsu_exe_0_req_bits_uop_ldst_val),
    .io_lsu_exe_0_req_bits_uop_dst_rtype(core_io_lsu_exe_0_req_bits_uop_dst_rtype),
    .io_lsu_exe_0_req_bits_uop_lrs1_rtype(core_io_lsu_exe_0_req_bits_uop_lrs1_rtype),
    .io_lsu_exe_0_req_bits_uop_lrs2_rtype(core_io_lsu_exe_0_req_bits_uop_lrs2_rtype),
    .io_lsu_exe_0_req_bits_uop_frs3_en(core_io_lsu_exe_0_req_bits_uop_frs3_en),
    .io_lsu_exe_0_req_bits_uop_fp_val(core_io_lsu_exe_0_req_bits_uop_fp_val),
    .io_lsu_exe_0_req_bits_uop_fp_single(core_io_lsu_exe_0_req_bits_uop_fp_single),
    .io_lsu_exe_0_req_bits_uop_xcpt_pf_if(core_io_lsu_exe_0_req_bits_uop_xcpt_pf_if),
    .io_lsu_exe_0_req_bits_uop_xcpt_ae_if(core_io_lsu_exe_0_req_bits_uop_xcpt_ae_if),
    .io_lsu_exe_0_req_bits_uop_xcpt_ma_if(core_io_lsu_exe_0_req_bits_uop_xcpt_ma_if),
    .io_lsu_exe_0_req_bits_uop_bp_debug_if(core_io_lsu_exe_0_req_bits_uop_bp_debug_if),
    .io_lsu_exe_0_req_bits_uop_bp_xcpt_if(core_io_lsu_exe_0_req_bits_uop_bp_xcpt_if),
    .io_lsu_exe_0_req_bits_uop_debug_fsrc(core_io_lsu_exe_0_req_bits_uop_debug_fsrc),
    .io_lsu_exe_0_req_bits_uop_debug_tsrc(core_io_lsu_exe_0_req_bits_uop_debug_tsrc),
    .io_lsu_exe_0_req_bits_predicated(core_io_lsu_exe_0_req_bits_predicated),
    .io_lsu_exe_0_req_bits_data(core_io_lsu_exe_0_req_bits_data),
    .io_lsu_exe_0_req_bits_fflags_valid(core_io_lsu_exe_0_req_bits_fflags_valid),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_switch(core_io_lsu_exe_0_req_bits_fflags_bits_uop_switch),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_switch_off(core_io_lsu_exe_0_req_bits_fflags_bits_uop_switch_off),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_is_unicore(core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_unicore),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_shift(core_io_lsu_exe_0_req_bits_fflags_bits_uop_shift),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_lrs3_rtype(core_io_lsu_exe_0_req_bits_fflags_bits_uop_lrs3_rtype),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_rflag(core_io_lsu_exe_0_req_bits_fflags_bits_uop_rflag),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_wflag(core_io_lsu_exe_0_req_bits_fflags_bits_uop_wflag),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_prflag(core_io_lsu_exe_0_req_bits_fflags_bits_uop_prflag),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_pwflag(core_io_lsu_exe_0_req_bits_fflags_bits_uop_pwflag),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_pflag_busy(core_io_lsu_exe_0_req_bits_fflags_bits_uop_pflag_busy),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_stale_pflag(core_io_lsu_exe_0_req_bits_fflags_bits_uop_stale_pflag),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_op1_sel(core_io_lsu_exe_0_req_bits_fflags_bits_uop_op1_sel),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_op2_sel(core_io_lsu_exe_0_req_bits_fflags_bits_uop_op2_sel),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_split_num(core_io_lsu_exe_0_req_bits_fflags_bits_uop_split_num),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_self_index(core_io_lsu_exe_0_req_bits_fflags_bits_uop_self_index),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_rob_inst_idx(core_io_lsu_exe_0_req_bits_fflags_bits_uop_rob_inst_idx),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_address_num(core_io_lsu_exe_0_req_bits_fflags_bits_uop_address_num),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_uopc(core_io_lsu_exe_0_req_bits_fflags_bits_uop_uopc),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_inst(core_io_lsu_exe_0_req_bits_fflags_bits_uop_inst),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_debug_inst(core_io_lsu_exe_0_req_bits_fflags_bits_uop_debug_inst),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_is_rvc(core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_rvc),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_debug_pc(core_io_lsu_exe_0_req_bits_fflags_bits_uop_debug_pc),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_iq_type(core_io_lsu_exe_0_req_bits_fflags_bits_uop_iq_type),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_fu_code(core_io_lsu_exe_0_req_bits_fflags_bits_uop_fu_code),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_br_type(core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_br_type),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_op1_sel(core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_op1_sel),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_op2_sel(core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_op2_sel),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_imm_sel(core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_imm_sel),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_op_fcn(core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_op_fcn),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_fcn_dw(core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_fcn_dw),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_csr_cmd(core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_csr_cmd),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_is_load(core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_is_load),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_is_sta(core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_is_sta),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_is_std(core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_is_std),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_op3_sel(core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_op3_sel),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_iw_state(core_io_lsu_exe_0_req_bits_fflags_bits_uop_iw_state),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_iw_p1_poisoned(core_io_lsu_exe_0_req_bits_fflags_bits_uop_iw_p1_poisoned),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_iw_p2_poisoned(core_io_lsu_exe_0_req_bits_fflags_bits_uop_iw_p2_poisoned),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_is_br(core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_br),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_is_jalr(core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_jalr),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_is_jal(core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_jal),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_is_sfb(core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_sfb),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_br_mask(core_io_lsu_exe_0_req_bits_fflags_bits_uop_br_mask),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_br_tag(core_io_lsu_exe_0_req_bits_fflags_bits_uop_br_tag),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_ftq_idx(core_io_lsu_exe_0_req_bits_fflags_bits_uop_ftq_idx),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_edge_inst(core_io_lsu_exe_0_req_bits_fflags_bits_uop_edge_inst),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_pc_lob(core_io_lsu_exe_0_req_bits_fflags_bits_uop_pc_lob),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_taken(core_io_lsu_exe_0_req_bits_fflags_bits_uop_taken),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_imm_packed(core_io_lsu_exe_0_req_bits_fflags_bits_uop_imm_packed),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_csr_addr(core_io_lsu_exe_0_req_bits_fflags_bits_uop_csr_addr),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_rob_idx(core_io_lsu_exe_0_req_bits_fflags_bits_uop_rob_idx),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_ldq_idx(core_io_lsu_exe_0_req_bits_fflags_bits_uop_ldq_idx),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_stq_idx(core_io_lsu_exe_0_req_bits_fflags_bits_uop_stq_idx),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_rxq_idx(core_io_lsu_exe_0_req_bits_fflags_bits_uop_rxq_idx),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_pdst(core_io_lsu_exe_0_req_bits_fflags_bits_uop_pdst),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_prs1(core_io_lsu_exe_0_req_bits_fflags_bits_uop_prs1),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_prs2(core_io_lsu_exe_0_req_bits_fflags_bits_uop_prs2),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_prs3(core_io_lsu_exe_0_req_bits_fflags_bits_uop_prs3),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_ppred(core_io_lsu_exe_0_req_bits_fflags_bits_uop_ppred),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_prs1_busy(core_io_lsu_exe_0_req_bits_fflags_bits_uop_prs1_busy),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_prs2_busy(core_io_lsu_exe_0_req_bits_fflags_bits_uop_prs2_busy),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_prs3_busy(core_io_lsu_exe_0_req_bits_fflags_bits_uop_prs3_busy),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_ppred_busy(core_io_lsu_exe_0_req_bits_fflags_bits_uop_ppred_busy),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_stale_pdst(core_io_lsu_exe_0_req_bits_fflags_bits_uop_stale_pdst),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_exception(core_io_lsu_exe_0_req_bits_fflags_bits_uop_exception),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_exc_cause(core_io_lsu_exe_0_req_bits_fflags_bits_uop_exc_cause),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_bypassable(core_io_lsu_exe_0_req_bits_fflags_bits_uop_bypassable),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_mem_cmd(core_io_lsu_exe_0_req_bits_fflags_bits_uop_mem_cmd),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_mem_size(core_io_lsu_exe_0_req_bits_fflags_bits_uop_mem_size),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_mem_signed(core_io_lsu_exe_0_req_bits_fflags_bits_uop_mem_signed),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_is_fence(core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_fence),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_is_fencei(core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_fencei),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_is_amo(core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_amo),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_uses_ldq(core_io_lsu_exe_0_req_bits_fflags_bits_uop_uses_ldq),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_uses_stq(core_io_lsu_exe_0_req_bits_fflags_bits_uop_uses_stq),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_is_sys_pc2epc(core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_sys_pc2epc),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_is_unique(core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_unique),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_flush_on_commit(core_io_lsu_exe_0_req_bits_fflags_bits_uop_flush_on_commit),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_ldst_is_rs1(core_io_lsu_exe_0_req_bits_fflags_bits_uop_ldst_is_rs1),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_ldst(core_io_lsu_exe_0_req_bits_fflags_bits_uop_ldst),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_lrs1(core_io_lsu_exe_0_req_bits_fflags_bits_uop_lrs1),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_lrs2(core_io_lsu_exe_0_req_bits_fflags_bits_uop_lrs2),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_lrs3(core_io_lsu_exe_0_req_bits_fflags_bits_uop_lrs3),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_ldst_val(core_io_lsu_exe_0_req_bits_fflags_bits_uop_ldst_val),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_dst_rtype(core_io_lsu_exe_0_req_bits_fflags_bits_uop_dst_rtype),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_lrs1_rtype(core_io_lsu_exe_0_req_bits_fflags_bits_uop_lrs1_rtype),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_lrs2_rtype(core_io_lsu_exe_0_req_bits_fflags_bits_uop_lrs2_rtype),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_frs3_en(core_io_lsu_exe_0_req_bits_fflags_bits_uop_frs3_en),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_fp_val(core_io_lsu_exe_0_req_bits_fflags_bits_uop_fp_val),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_fp_single(core_io_lsu_exe_0_req_bits_fflags_bits_uop_fp_single),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_xcpt_pf_if(core_io_lsu_exe_0_req_bits_fflags_bits_uop_xcpt_pf_if),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_xcpt_ae_if(core_io_lsu_exe_0_req_bits_fflags_bits_uop_xcpt_ae_if),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_xcpt_ma_if(core_io_lsu_exe_0_req_bits_fflags_bits_uop_xcpt_ma_if),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_bp_debug_if(core_io_lsu_exe_0_req_bits_fflags_bits_uop_bp_debug_if),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_bp_xcpt_if(core_io_lsu_exe_0_req_bits_fflags_bits_uop_bp_xcpt_if),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_debug_fsrc(core_io_lsu_exe_0_req_bits_fflags_bits_uop_debug_fsrc),
    .io_lsu_exe_0_req_bits_fflags_bits_uop_debug_tsrc(core_io_lsu_exe_0_req_bits_fflags_bits_uop_debug_tsrc),
    .io_lsu_exe_0_req_bits_fflags_bits_flags(core_io_lsu_exe_0_req_bits_fflags_bits_flags),
    .io_lsu_exe_0_req_bits_addr(core_io_lsu_exe_0_req_bits_addr),
    .io_lsu_exe_0_req_bits_mxcpt_valid(core_io_lsu_exe_0_req_bits_mxcpt_valid),
    .io_lsu_exe_0_req_bits_mxcpt_bits(core_io_lsu_exe_0_req_bits_mxcpt_bits),
    .io_lsu_exe_0_req_bits_sfence_valid(core_io_lsu_exe_0_req_bits_sfence_valid),
    .io_lsu_exe_0_req_bits_sfence_bits_rs1(core_io_lsu_exe_0_req_bits_sfence_bits_rs1),
    .io_lsu_exe_0_req_bits_sfence_bits_rs2(core_io_lsu_exe_0_req_bits_sfence_bits_rs2),
    .io_lsu_exe_0_req_bits_sfence_bits_addr(core_io_lsu_exe_0_req_bits_sfence_bits_addr),
    .io_lsu_exe_0_req_bits_sfence_bits_asid(core_io_lsu_exe_0_req_bits_sfence_bits_asid),
    .io_lsu_exe_0_req_bits_flagdata(core_io_lsu_exe_0_req_bits_flagdata),
    .io_lsu_exe_0_req_bits_fflagdata_valid(core_io_lsu_exe_0_req_bits_fflagdata_valid),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_switch(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_switch),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_switch_off(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_switch_off),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_unicore(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_unicore),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_shift(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_shift),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs3_rtype(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs3_rtype),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_rflag(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_rflag),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_wflag(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_wflag),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_prflag(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_prflag),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_pwflag(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_pwflag),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_pflag_busy(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_pflag_busy),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_stale_pflag(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_stale_pflag),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_op1_sel(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_op1_sel),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_op2_sel(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_op2_sel),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_split_num(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_split_num),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_self_index(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_self_index),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_rob_inst_idx(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_rob_inst_idx),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_address_num(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_address_num),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_uopc(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_uopc),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_inst(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_inst),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_debug_inst(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_debug_inst),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_rvc(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_rvc),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_debug_pc(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_debug_pc),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_iq_type(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_iq_type),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_fu_code(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_fu_code),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_br_type(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_br_type),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_op1_sel(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_op1_sel),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_op2_sel(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_op2_sel),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_imm_sel(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_imm_sel),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_op_fcn(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_op_fcn),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_fcn_dw(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_fcn_dw),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_csr_cmd(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_csr_cmd),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_load(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_load),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_sta(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_sta),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_std(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_std),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_op3_sel(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_op3_sel),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_iw_state(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_iw_state),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_iw_p1_poisoned(
      core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_iw_p1_poisoned),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_iw_p2_poisoned(
      core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_iw_p2_poisoned),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_br(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_br),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_jalr(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_jalr),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_jal(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_jal),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_sfb(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_sfb),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_br_mask(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_br_mask),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_br_tag(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_br_tag),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_ftq_idx(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ftq_idx),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_edge_inst(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_edge_inst),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_pc_lob(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_pc_lob),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_taken(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_taken),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_imm_packed(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_imm_packed),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_csr_addr(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_csr_addr),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_rob_idx(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_rob_idx),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_ldq_idx(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ldq_idx),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_stq_idx(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_stq_idx),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_rxq_idx(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_rxq_idx),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_pdst(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_pdst),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs1(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs1),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs2(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs2),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs3(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs3),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_ppred(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ppred),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs1_busy(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs1_busy),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs2_busy(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs2_busy),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs3_busy(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs3_busy),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_ppred_busy(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ppred_busy),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_stale_pdst(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_stale_pdst),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_exception(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_exception),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_exc_cause(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_exc_cause),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_bypassable(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_bypassable),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_mem_cmd(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_mem_cmd),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_mem_size(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_mem_size),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_mem_signed(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_mem_signed),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_fence(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_fence),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_fencei(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_fencei),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_amo(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_amo),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_uses_ldq(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_uses_ldq),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_uses_stq(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_uses_stq),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_sys_pc2epc(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_sys_pc2epc)
      ,
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_unique(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_unique),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_flush_on_commit(
      core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_flush_on_commit),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_ldst_is_rs1(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ldst_is_rs1),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_ldst(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ldst),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs1(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs1),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs2(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs2),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs3(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs3),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_ldst_val(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ldst_val),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_dst_rtype(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_dst_rtype),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs1_rtype(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs1_rtype),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs2_rtype(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs2_rtype),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_frs3_en(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_frs3_en),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_fp_val(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_fp_val),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_fp_single(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_fp_single),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_xcpt_pf_if(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_xcpt_pf_if),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_xcpt_ae_if(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_xcpt_ae_if),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_xcpt_ma_if(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_xcpt_ma_if),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_bp_debug_if(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_bp_debug_if),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_bp_xcpt_if(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_bp_xcpt_if),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_debug_fsrc(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_debug_fsrc),
    .io_lsu_exe_0_req_bits_fflagdata_bits_uop_debug_tsrc(core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_debug_tsrc),
    .io_lsu_exe_0_req_bits_fflagdata_bits_fflag(core_io_lsu_exe_0_req_bits_fflagdata_bits_fflag),
    .io_lsu_exe_0_iresp_ready(core_io_lsu_exe_0_iresp_ready),
    .io_lsu_exe_0_iresp_valid(core_io_lsu_exe_0_iresp_valid),
    .io_lsu_exe_0_iresp_bits_uop_switch(core_io_lsu_exe_0_iresp_bits_uop_switch),
    .io_lsu_exe_0_iresp_bits_uop_switch_off(core_io_lsu_exe_0_iresp_bits_uop_switch_off),
    .io_lsu_exe_0_iresp_bits_uop_is_unicore(core_io_lsu_exe_0_iresp_bits_uop_is_unicore),
    .io_lsu_exe_0_iresp_bits_uop_shift(core_io_lsu_exe_0_iresp_bits_uop_shift),
    .io_lsu_exe_0_iresp_bits_uop_lrs3_rtype(core_io_lsu_exe_0_iresp_bits_uop_lrs3_rtype),
    .io_lsu_exe_0_iresp_bits_uop_rflag(core_io_lsu_exe_0_iresp_bits_uop_rflag),
    .io_lsu_exe_0_iresp_bits_uop_wflag(core_io_lsu_exe_0_iresp_bits_uop_wflag),
    .io_lsu_exe_0_iresp_bits_uop_prflag(core_io_lsu_exe_0_iresp_bits_uop_prflag),
    .io_lsu_exe_0_iresp_bits_uop_pwflag(core_io_lsu_exe_0_iresp_bits_uop_pwflag),
    .io_lsu_exe_0_iresp_bits_uop_pflag_busy(core_io_lsu_exe_0_iresp_bits_uop_pflag_busy),
    .io_lsu_exe_0_iresp_bits_uop_stale_pflag(core_io_lsu_exe_0_iresp_bits_uop_stale_pflag),
    .io_lsu_exe_0_iresp_bits_uop_op1_sel(core_io_lsu_exe_0_iresp_bits_uop_op1_sel),
    .io_lsu_exe_0_iresp_bits_uop_op2_sel(core_io_lsu_exe_0_iresp_bits_uop_op2_sel),
    .io_lsu_exe_0_iresp_bits_uop_split_num(core_io_lsu_exe_0_iresp_bits_uop_split_num),
    .io_lsu_exe_0_iresp_bits_uop_self_index(core_io_lsu_exe_0_iresp_bits_uop_self_index),
    .io_lsu_exe_0_iresp_bits_uop_rob_inst_idx(core_io_lsu_exe_0_iresp_bits_uop_rob_inst_idx),
    .io_lsu_exe_0_iresp_bits_uop_address_num(core_io_lsu_exe_0_iresp_bits_uop_address_num),
    .io_lsu_exe_0_iresp_bits_uop_uopc(core_io_lsu_exe_0_iresp_bits_uop_uopc),
    .io_lsu_exe_0_iresp_bits_uop_inst(core_io_lsu_exe_0_iresp_bits_uop_inst),
    .io_lsu_exe_0_iresp_bits_uop_debug_inst(core_io_lsu_exe_0_iresp_bits_uop_debug_inst),
    .io_lsu_exe_0_iresp_bits_uop_is_rvc(core_io_lsu_exe_0_iresp_bits_uop_is_rvc),
    .io_lsu_exe_0_iresp_bits_uop_debug_pc(core_io_lsu_exe_0_iresp_bits_uop_debug_pc),
    .io_lsu_exe_0_iresp_bits_uop_iq_type(core_io_lsu_exe_0_iresp_bits_uop_iq_type),
    .io_lsu_exe_0_iresp_bits_uop_fu_code(core_io_lsu_exe_0_iresp_bits_uop_fu_code),
    .io_lsu_exe_0_iresp_bits_uop_ctrl_br_type(core_io_lsu_exe_0_iresp_bits_uop_ctrl_br_type),
    .io_lsu_exe_0_iresp_bits_uop_ctrl_op1_sel(core_io_lsu_exe_0_iresp_bits_uop_ctrl_op1_sel),
    .io_lsu_exe_0_iresp_bits_uop_ctrl_op2_sel(core_io_lsu_exe_0_iresp_bits_uop_ctrl_op2_sel),
    .io_lsu_exe_0_iresp_bits_uop_ctrl_imm_sel(core_io_lsu_exe_0_iresp_bits_uop_ctrl_imm_sel),
    .io_lsu_exe_0_iresp_bits_uop_ctrl_op_fcn(core_io_lsu_exe_0_iresp_bits_uop_ctrl_op_fcn),
    .io_lsu_exe_0_iresp_bits_uop_ctrl_fcn_dw(core_io_lsu_exe_0_iresp_bits_uop_ctrl_fcn_dw),
    .io_lsu_exe_0_iresp_bits_uop_ctrl_csr_cmd(core_io_lsu_exe_0_iresp_bits_uop_ctrl_csr_cmd),
    .io_lsu_exe_0_iresp_bits_uop_ctrl_is_load(core_io_lsu_exe_0_iresp_bits_uop_ctrl_is_load),
    .io_lsu_exe_0_iresp_bits_uop_ctrl_is_sta(core_io_lsu_exe_0_iresp_bits_uop_ctrl_is_sta),
    .io_lsu_exe_0_iresp_bits_uop_ctrl_is_std(core_io_lsu_exe_0_iresp_bits_uop_ctrl_is_std),
    .io_lsu_exe_0_iresp_bits_uop_ctrl_op3_sel(core_io_lsu_exe_0_iresp_bits_uop_ctrl_op3_sel),
    .io_lsu_exe_0_iresp_bits_uop_iw_state(core_io_lsu_exe_0_iresp_bits_uop_iw_state),
    .io_lsu_exe_0_iresp_bits_uop_iw_p1_poisoned(core_io_lsu_exe_0_iresp_bits_uop_iw_p1_poisoned),
    .io_lsu_exe_0_iresp_bits_uop_iw_p2_poisoned(core_io_lsu_exe_0_iresp_bits_uop_iw_p2_poisoned),
    .io_lsu_exe_0_iresp_bits_uop_is_br(core_io_lsu_exe_0_iresp_bits_uop_is_br),
    .io_lsu_exe_0_iresp_bits_uop_is_jalr(core_io_lsu_exe_0_iresp_bits_uop_is_jalr),
    .io_lsu_exe_0_iresp_bits_uop_is_jal(core_io_lsu_exe_0_iresp_bits_uop_is_jal),
    .io_lsu_exe_0_iresp_bits_uop_is_sfb(core_io_lsu_exe_0_iresp_bits_uop_is_sfb),
    .io_lsu_exe_0_iresp_bits_uop_br_mask(core_io_lsu_exe_0_iresp_bits_uop_br_mask),
    .io_lsu_exe_0_iresp_bits_uop_br_tag(core_io_lsu_exe_0_iresp_bits_uop_br_tag),
    .io_lsu_exe_0_iresp_bits_uop_ftq_idx(core_io_lsu_exe_0_iresp_bits_uop_ftq_idx),
    .io_lsu_exe_0_iresp_bits_uop_edge_inst(core_io_lsu_exe_0_iresp_bits_uop_edge_inst),
    .io_lsu_exe_0_iresp_bits_uop_pc_lob(core_io_lsu_exe_0_iresp_bits_uop_pc_lob),
    .io_lsu_exe_0_iresp_bits_uop_taken(core_io_lsu_exe_0_iresp_bits_uop_taken),
    .io_lsu_exe_0_iresp_bits_uop_imm_packed(core_io_lsu_exe_0_iresp_bits_uop_imm_packed),
    .io_lsu_exe_0_iresp_bits_uop_csr_addr(core_io_lsu_exe_0_iresp_bits_uop_csr_addr),
    .io_lsu_exe_0_iresp_bits_uop_rob_idx(core_io_lsu_exe_0_iresp_bits_uop_rob_idx),
    .io_lsu_exe_0_iresp_bits_uop_ldq_idx(core_io_lsu_exe_0_iresp_bits_uop_ldq_idx),
    .io_lsu_exe_0_iresp_bits_uop_stq_idx(core_io_lsu_exe_0_iresp_bits_uop_stq_idx),
    .io_lsu_exe_0_iresp_bits_uop_rxq_idx(core_io_lsu_exe_0_iresp_bits_uop_rxq_idx),
    .io_lsu_exe_0_iresp_bits_uop_pdst(core_io_lsu_exe_0_iresp_bits_uop_pdst),
    .io_lsu_exe_0_iresp_bits_uop_prs1(core_io_lsu_exe_0_iresp_bits_uop_prs1),
    .io_lsu_exe_0_iresp_bits_uop_prs2(core_io_lsu_exe_0_iresp_bits_uop_prs2),
    .io_lsu_exe_0_iresp_bits_uop_prs3(core_io_lsu_exe_0_iresp_bits_uop_prs3),
    .io_lsu_exe_0_iresp_bits_uop_ppred(core_io_lsu_exe_0_iresp_bits_uop_ppred),
    .io_lsu_exe_0_iresp_bits_uop_prs1_busy(core_io_lsu_exe_0_iresp_bits_uop_prs1_busy),
    .io_lsu_exe_0_iresp_bits_uop_prs2_busy(core_io_lsu_exe_0_iresp_bits_uop_prs2_busy),
    .io_lsu_exe_0_iresp_bits_uop_prs3_busy(core_io_lsu_exe_0_iresp_bits_uop_prs3_busy),
    .io_lsu_exe_0_iresp_bits_uop_ppred_busy(core_io_lsu_exe_0_iresp_bits_uop_ppred_busy),
    .io_lsu_exe_0_iresp_bits_uop_stale_pdst(core_io_lsu_exe_0_iresp_bits_uop_stale_pdst),
    .io_lsu_exe_0_iresp_bits_uop_exception(core_io_lsu_exe_0_iresp_bits_uop_exception),
    .io_lsu_exe_0_iresp_bits_uop_exc_cause(core_io_lsu_exe_0_iresp_bits_uop_exc_cause),
    .io_lsu_exe_0_iresp_bits_uop_bypassable(core_io_lsu_exe_0_iresp_bits_uop_bypassable),
    .io_lsu_exe_0_iresp_bits_uop_mem_cmd(core_io_lsu_exe_0_iresp_bits_uop_mem_cmd),
    .io_lsu_exe_0_iresp_bits_uop_mem_size(core_io_lsu_exe_0_iresp_bits_uop_mem_size),
    .io_lsu_exe_0_iresp_bits_uop_mem_signed(core_io_lsu_exe_0_iresp_bits_uop_mem_signed),
    .io_lsu_exe_0_iresp_bits_uop_is_fence(core_io_lsu_exe_0_iresp_bits_uop_is_fence),
    .io_lsu_exe_0_iresp_bits_uop_is_fencei(core_io_lsu_exe_0_iresp_bits_uop_is_fencei),
    .io_lsu_exe_0_iresp_bits_uop_is_amo(core_io_lsu_exe_0_iresp_bits_uop_is_amo),
    .io_lsu_exe_0_iresp_bits_uop_uses_ldq(core_io_lsu_exe_0_iresp_bits_uop_uses_ldq),
    .io_lsu_exe_0_iresp_bits_uop_uses_stq(core_io_lsu_exe_0_iresp_bits_uop_uses_stq),
    .io_lsu_exe_0_iresp_bits_uop_is_sys_pc2epc(core_io_lsu_exe_0_iresp_bits_uop_is_sys_pc2epc),
    .io_lsu_exe_0_iresp_bits_uop_is_unique(core_io_lsu_exe_0_iresp_bits_uop_is_unique),
    .io_lsu_exe_0_iresp_bits_uop_flush_on_commit(core_io_lsu_exe_0_iresp_bits_uop_flush_on_commit),
    .io_lsu_exe_0_iresp_bits_uop_ldst_is_rs1(core_io_lsu_exe_0_iresp_bits_uop_ldst_is_rs1),
    .io_lsu_exe_0_iresp_bits_uop_ldst(core_io_lsu_exe_0_iresp_bits_uop_ldst),
    .io_lsu_exe_0_iresp_bits_uop_lrs1(core_io_lsu_exe_0_iresp_bits_uop_lrs1),
    .io_lsu_exe_0_iresp_bits_uop_lrs2(core_io_lsu_exe_0_iresp_bits_uop_lrs2),
    .io_lsu_exe_0_iresp_bits_uop_lrs3(core_io_lsu_exe_0_iresp_bits_uop_lrs3),
    .io_lsu_exe_0_iresp_bits_uop_ldst_val(core_io_lsu_exe_0_iresp_bits_uop_ldst_val),
    .io_lsu_exe_0_iresp_bits_uop_dst_rtype(core_io_lsu_exe_0_iresp_bits_uop_dst_rtype),
    .io_lsu_exe_0_iresp_bits_uop_lrs1_rtype(core_io_lsu_exe_0_iresp_bits_uop_lrs1_rtype),
    .io_lsu_exe_0_iresp_bits_uop_lrs2_rtype(core_io_lsu_exe_0_iresp_bits_uop_lrs2_rtype),
    .io_lsu_exe_0_iresp_bits_uop_frs3_en(core_io_lsu_exe_0_iresp_bits_uop_frs3_en),
    .io_lsu_exe_0_iresp_bits_uop_fp_val(core_io_lsu_exe_0_iresp_bits_uop_fp_val),
    .io_lsu_exe_0_iresp_bits_uop_fp_single(core_io_lsu_exe_0_iresp_bits_uop_fp_single),
    .io_lsu_exe_0_iresp_bits_uop_xcpt_pf_if(core_io_lsu_exe_0_iresp_bits_uop_xcpt_pf_if),
    .io_lsu_exe_0_iresp_bits_uop_xcpt_ae_if(core_io_lsu_exe_0_iresp_bits_uop_xcpt_ae_if),
    .io_lsu_exe_0_iresp_bits_uop_xcpt_ma_if(core_io_lsu_exe_0_iresp_bits_uop_xcpt_ma_if),
    .io_lsu_exe_0_iresp_bits_uop_bp_debug_if(core_io_lsu_exe_0_iresp_bits_uop_bp_debug_if),
    .io_lsu_exe_0_iresp_bits_uop_bp_xcpt_if(core_io_lsu_exe_0_iresp_bits_uop_bp_xcpt_if),
    .io_lsu_exe_0_iresp_bits_uop_debug_fsrc(core_io_lsu_exe_0_iresp_bits_uop_debug_fsrc),
    .io_lsu_exe_0_iresp_bits_uop_debug_tsrc(core_io_lsu_exe_0_iresp_bits_uop_debug_tsrc),
    .io_lsu_exe_0_iresp_bits_data(core_io_lsu_exe_0_iresp_bits_data),
    .io_lsu_exe_0_iresp_bits_predicated(core_io_lsu_exe_0_iresp_bits_predicated),
    .io_lsu_exe_0_iresp_bits_fflags_valid(core_io_lsu_exe_0_iresp_bits_fflags_valid),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_switch(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_switch),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_switch_off(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_switch_off),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_unicore(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_unicore),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_shift(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_shift),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs3_rtype(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs3_rtype),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_rflag(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_rflag),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_wflag(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_wflag),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_prflag(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_prflag),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_pwflag(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_pwflag),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_pflag_busy(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_pflag_busy),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_stale_pflag(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_stale_pflag),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_op1_sel(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_op1_sel),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_op2_sel(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_op2_sel),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_split_num(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_split_num),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_self_index(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_self_index),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_rob_inst_idx(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_rob_inst_idx),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_address_num(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_address_num),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_uopc(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_uopc),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_inst(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_inst),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_debug_inst(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_debug_inst),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_rvc(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_rvc),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_debug_pc(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_debug_pc),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_iq_type(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_iq_type),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_fu_code(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_fu_code),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_br_type(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_br_type),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_op1_sel(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_op1_sel),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_op2_sel(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_op2_sel),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_imm_sel(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_imm_sel),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_op_fcn(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_op_fcn),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_fcn_dw(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_fcn_dw),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_csr_cmd(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_csr_cmd),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_load(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_load),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_sta(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_sta),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_std(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_std),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_op3_sel(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_op3_sel),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_iw_state(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_iw_state),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_iw_p1_poisoned(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_iw_p1_poisoned)
      ,
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_iw_p2_poisoned(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_iw_p2_poisoned)
      ,
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_br(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_br),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_jalr(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_jalr),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_jal(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_jal),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_sfb(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_sfb),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_br_mask(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_br_mask),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_br_tag(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_br_tag),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_ftq_idx(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ftq_idx),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_edge_inst(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_edge_inst),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_pc_lob(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_pc_lob),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_taken(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_taken),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_imm_packed(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_imm_packed),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_csr_addr(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_csr_addr),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_rob_idx(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_rob_idx),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_ldq_idx(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ldq_idx),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_stq_idx(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_stq_idx),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_rxq_idx(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_rxq_idx),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_pdst(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_pdst),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs1(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs1),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs2(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs2),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs3(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs3),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_ppred(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ppred),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs1_busy(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs1_busy),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs2_busy(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs2_busy),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs3_busy(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs3_busy),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_ppred_busy(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ppred_busy),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_stale_pdst(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_stale_pdst),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_exception(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_exception),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_exc_cause(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_exc_cause),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_bypassable(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_bypassable),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_mem_cmd(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_mem_cmd),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_mem_size(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_mem_size),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_mem_signed(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_mem_signed),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_fence(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_fence),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_fencei(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_fencei),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_amo(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_amo),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_uses_ldq(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_uses_ldq),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_uses_stq(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_uses_stq),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_sys_pc2epc(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_sys_pc2epc),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_unique(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_unique),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_flush_on_commit(
      core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_flush_on_commit),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_ldst_is_rs1(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ldst_is_rs1),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_ldst(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ldst),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs1(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs1),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs2(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs2),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs3(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs3),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_ldst_val(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ldst_val),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_dst_rtype(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_dst_rtype),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs1_rtype(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs1_rtype),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs2_rtype(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs2_rtype),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_frs3_en(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_frs3_en),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_fp_val(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_fp_val),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_fp_single(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_fp_single),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_xcpt_pf_if(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_xcpt_pf_if),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_xcpt_ae_if(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_xcpt_ae_if),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_xcpt_ma_if(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_xcpt_ma_if),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_bp_debug_if(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_bp_debug_if),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_bp_xcpt_if(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_bp_xcpt_if),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_debug_fsrc(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_debug_fsrc),
    .io_lsu_exe_0_iresp_bits_fflags_bits_uop_debug_tsrc(core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_debug_tsrc),
    .io_lsu_exe_0_iresp_bits_fflags_bits_flags(core_io_lsu_exe_0_iresp_bits_fflags_bits_flags),
    .io_lsu_exe_0_iresp_bits_flagdata(core_io_lsu_exe_0_iresp_bits_flagdata),
    .io_lsu_exe_0_iresp_bits_fflagdata_valid(core_io_lsu_exe_0_iresp_bits_fflagdata_valid),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_switch(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_switch),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_switch_off(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_switch_off),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_unicore(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_unicore),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_shift(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_shift),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs3_rtype(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs3_rtype),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_rflag(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_rflag),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_wflag(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_wflag),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prflag(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prflag),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_pwflag(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_pwflag),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_pflag_busy(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_pflag_busy),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_stale_pflag(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_stale_pflag)
      ,
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_op1_sel(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_op1_sel),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_op2_sel(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_op2_sel),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_split_num(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_split_num),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_self_index(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_self_index),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_rob_inst_idx(
      core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_rob_inst_idx),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_address_num(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_address_num)
      ,
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_uopc(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_uopc),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_inst(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_inst),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_debug_inst(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_debug_inst),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_rvc(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_rvc),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_debug_pc(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_debug_pc),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_iq_type(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_iq_type),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_fu_code(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_fu_code),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_br_type(
      core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_br_type),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op1_sel(
      core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op1_sel),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op2_sel(
      core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op2_sel),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_imm_sel(
      core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_imm_sel),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op_fcn(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op_fcn)
      ,
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_fcn_dw(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_fcn_dw)
      ,
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_csr_cmd(
      core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_csr_cmd),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_load(
      core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_load),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_sta(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_sta)
      ,
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_std(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_std)
      ,
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op3_sel(
      core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op3_sel),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_iw_state(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_iw_state),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_iw_p1_poisoned(
      core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_iw_p1_poisoned),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_iw_p2_poisoned(
      core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_iw_p2_poisoned),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_br(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_br),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_jalr(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_jalr),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_jal(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_jal),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_sfb(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_sfb),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_br_mask(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_br_mask),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_br_tag(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_br_tag),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ftq_idx(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ftq_idx),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_edge_inst(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_edge_inst),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_pc_lob(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_pc_lob),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_taken(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_taken),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_imm_packed(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_imm_packed),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_csr_addr(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_csr_addr),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_rob_idx(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_rob_idx),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ldq_idx(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ldq_idx),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_stq_idx(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_stq_idx),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_rxq_idx(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_rxq_idx),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_pdst(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_pdst),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs1(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs1),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs2(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs2),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs3(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs3),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ppred(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ppred),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs1_busy(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs1_busy),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs2_busy(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs2_busy),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs3_busy(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs3_busy),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ppred_busy(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ppred_busy),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_stale_pdst(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_stale_pdst),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_exception(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_exception),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_exc_cause(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_exc_cause),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_bypassable(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_bypassable),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_mem_cmd(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_mem_cmd),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_mem_size(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_mem_size),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_mem_signed(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_mem_signed),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_fence(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_fence),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_fencei(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_fencei),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_amo(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_amo),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_uses_ldq(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_uses_ldq),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_uses_stq(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_uses_stq),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_sys_pc2epc(
      core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_sys_pc2epc),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_unique(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_unique),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_flush_on_commit(
      core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_flush_on_commit),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ldst_is_rs1(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ldst_is_rs1)
      ,
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ldst(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ldst),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs1(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs1),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs2(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs2),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs3(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs3),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ldst_val(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ldst_val),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_dst_rtype(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_dst_rtype),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs1_rtype(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs1_rtype),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs2_rtype(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs2_rtype),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_frs3_en(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_frs3_en),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_fp_val(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_fp_val),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_fp_single(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_fp_single),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_pf_if(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_pf_if),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_ae_if(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_ae_if),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_ma_if(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_ma_if),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_bp_debug_if(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_bp_debug_if)
      ,
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_bp_xcpt_if(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_bp_xcpt_if),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_debug_fsrc(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_debug_fsrc),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_debug_tsrc(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_debug_tsrc),
    .io_lsu_exe_0_iresp_bits_fflagdata_bits_fflag(core_io_lsu_exe_0_iresp_bits_fflagdata_bits_fflag),
    .io_lsu_exe_0_fresp_ready(core_io_lsu_exe_0_fresp_ready),
    .io_lsu_exe_0_fresp_valid(core_io_lsu_exe_0_fresp_valid),
    .io_lsu_exe_0_fresp_bits_uop_switch(core_io_lsu_exe_0_fresp_bits_uop_switch),
    .io_lsu_exe_0_fresp_bits_uop_switch_off(core_io_lsu_exe_0_fresp_bits_uop_switch_off),
    .io_lsu_exe_0_fresp_bits_uop_is_unicore(core_io_lsu_exe_0_fresp_bits_uop_is_unicore),
    .io_lsu_exe_0_fresp_bits_uop_shift(core_io_lsu_exe_0_fresp_bits_uop_shift),
    .io_lsu_exe_0_fresp_bits_uop_lrs3_rtype(core_io_lsu_exe_0_fresp_bits_uop_lrs3_rtype),
    .io_lsu_exe_0_fresp_bits_uop_rflag(core_io_lsu_exe_0_fresp_bits_uop_rflag),
    .io_lsu_exe_0_fresp_bits_uop_wflag(core_io_lsu_exe_0_fresp_bits_uop_wflag),
    .io_lsu_exe_0_fresp_bits_uop_prflag(core_io_lsu_exe_0_fresp_bits_uop_prflag),
    .io_lsu_exe_0_fresp_bits_uop_pwflag(core_io_lsu_exe_0_fresp_bits_uop_pwflag),
    .io_lsu_exe_0_fresp_bits_uop_pflag_busy(core_io_lsu_exe_0_fresp_bits_uop_pflag_busy),
    .io_lsu_exe_0_fresp_bits_uop_stale_pflag(core_io_lsu_exe_0_fresp_bits_uop_stale_pflag),
    .io_lsu_exe_0_fresp_bits_uop_op1_sel(core_io_lsu_exe_0_fresp_bits_uop_op1_sel),
    .io_lsu_exe_0_fresp_bits_uop_op2_sel(core_io_lsu_exe_0_fresp_bits_uop_op2_sel),
    .io_lsu_exe_0_fresp_bits_uop_split_num(core_io_lsu_exe_0_fresp_bits_uop_split_num),
    .io_lsu_exe_0_fresp_bits_uop_self_index(core_io_lsu_exe_0_fresp_bits_uop_self_index),
    .io_lsu_exe_0_fresp_bits_uop_rob_inst_idx(core_io_lsu_exe_0_fresp_bits_uop_rob_inst_idx),
    .io_lsu_exe_0_fresp_bits_uop_address_num(core_io_lsu_exe_0_fresp_bits_uop_address_num),
    .io_lsu_exe_0_fresp_bits_uop_uopc(core_io_lsu_exe_0_fresp_bits_uop_uopc),
    .io_lsu_exe_0_fresp_bits_uop_inst(core_io_lsu_exe_0_fresp_bits_uop_inst),
    .io_lsu_exe_0_fresp_bits_uop_debug_inst(core_io_lsu_exe_0_fresp_bits_uop_debug_inst),
    .io_lsu_exe_0_fresp_bits_uop_is_rvc(core_io_lsu_exe_0_fresp_bits_uop_is_rvc),
    .io_lsu_exe_0_fresp_bits_uop_debug_pc(core_io_lsu_exe_0_fresp_bits_uop_debug_pc),
    .io_lsu_exe_0_fresp_bits_uop_iq_type(core_io_lsu_exe_0_fresp_bits_uop_iq_type),
    .io_lsu_exe_0_fresp_bits_uop_fu_code(core_io_lsu_exe_0_fresp_bits_uop_fu_code),
    .io_lsu_exe_0_fresp_bits_uop_ctrl_br_type(core_io_lsu_exe_0_fresp_bits_uop_ctrl_br_type),
    .io_lsu_exe_0_fresp_bits_uop_ctrl_op1_sel(core_io_lsu_exe_0_fresp_bits_uop_ctrl_op1_sel),
    .io_lsu_exe_0_fresp_bits_uop_ctrl_op2_sel(core_io_lsu_exe_0_fresp_bits_uop_ctrl_op2_sel),
    .io_lsu_exe_0_fresp_bits_uop_ctrl_imm_sel(core_io_lsu_exe_0_fresp_bits_uop_ctrl_imm_sel),
    .io_lsu_exe_0_fresp_bits_uop_ctrl_op_fcn(core_io_lsu_exe_0_fresp_bits_uop_ctrl_op_fcn),
    .io_lsu_exe_0_fresp_bits_uop_ctrl_fcn_dw(core_io_lsu_exe_0_fresp_bits_uop_ctrl_fcn_dw),
    .io_lsu_exe_0_fresp_bits_uop_ctrl_csr_cmd(core_io_lsu_exe_0_fresp_bits_uop_ctrl_csr_cmd),
    .io_lsu_exe_0_fresp_bits_uop_ctrl_is_load(core_io_lsu_exe_0_fresp_bits_uop_ctrl_is_load),
    .io_lsu_exe_0_fresp_bits_uop_ctrl_is_sta(core_io_lsu_exe_0_fresp_bits_uop_ctrl_is_sta),
    .io_lsu_exe_0_fresp_bits_uop_ctrl_is_std(core_io_lsu_exe_0_fresp_bits_uop_ctrl_is_std),
    .io_lsu_exe_0_fresp_bits_uop_ctrl_op3_sel(core_io_lsu_exe_0_fresp_bits_uop_ctrl_op3_sel),
    .io_lsu_exe_0_fresp_bits_uop_iw_state(core_io_lsu_exe_0_fresp_bits_uop_iw_state),
    .io_lsu_exe_0_fresp_bits_uop_iw_p1_poisoned(core_io_lsu_exe_0_fresp_bits_uop_iw_p1_poisoned),
    .io_lsu_exe_0_fresp_bits_uop_iw_p2_poisoned(core_io_lsu_exe_0_fresp_bits_uop_iw_p2_poisoned),
    .io_lsu_exe_0_fresp_bits_uop_is_br(core_io_lsu_exe_0_fresp_bits_uop_is_br),
    .io_lsu_exe_0_fresp_bits_uop_is_jalr(core_io_lsu_exe_0_fresp_bits_uop_is_jalr),
    .io_lsu_exe_0_fresp_bits_uop_is_jal(core_io_lsu_exe_0_fresp_bits_uop_is_jal),
    .io_lsu_exe_0_fresp_bits_uop_is_sfb(core_io_lsu_exe_0_fresp_bits_uop_is_sfb),
    .io_lsu_exe_0_fresp_bits_uop_br_mask(core_io_lsu_exe_0_fresp_bits_uop_br_mask),
    .io_lsu_exe_0_fresp_bits_uop_br_tag(core_io_lsu_exe_0_fresp_bits_uop_br_tag),
    .io_lsu_exe_0_fresp_bits_uop_ftq_idx(core_io_lsu_exe_0_fresp_bits_uop_ftq_idx),
    .io_lsu_exe_0_fresp_bits_uop_edge_inst(core_io_lsu_exe_0_fresp_bits_uop_edge_inst),
    .io_lsu_exe_0_fresp_bits_uop_pc_lob(core_io_lsu_exe_0_fresp_bits_uop_pc_lob),
    .io_lsu_exe_0_fresp_bits_uop_taken(core_io_lsu_exe_0_fresp_bits_uop_taken),
    .io_lsu_exe_0_fresp_bits_uop_imm_packed(core_io_lsu_exe_0_fresp_bits_uop_imm_packed),
    .io_lsu_exe_0_fresp_bits_uop_csr_addr(core_io_lsu_exe_0_fresp_bits_uop_csr_addr),
    .io_lsu_exe_0_fresp_bits_uop_rob_idx(core_io_lsu_exe_0_fresp_bits_uop_rob_idx),
    .io_lsu_exe_0_fresp_bits_uop_ldq_idx(core_io_lsu_exe_0_fresp_bits_uop_ldq_idx),
    .io_lsu_exe_0_fresp_bits_uop_stq_idx(core_io_lsu_exe_0_fresp_bits_uop_stq_idx),
    .io_lsu_exe_0_fresp_bits_uop_rxq_idx(core_io_lsu_exe_0_fresp_bits_uop_rxq_idx),
    .io_lsu_exe_0_fresp_bits_uop_pdst(core_io_lsu_exe_0_fresp_bits_uop_pdst),
    .io_lsu_exe_0_fresp_bits_uop_prs1(core_io_lsu_exe_0_fresp_bits_uop_prs1),
    .io_lsu_exe_0_fresp_bits_uop_prs2(core_io_lsu_exe_0_fresp_bits_uop_prs2),
    .io_lsu_exe_0_fresp_bits_uop_prs3(core_io_lsu_exe_0_fresp_bits_uop_prs3),
    .io_lsu_exe_0_fresp_bits_uop_ppred(core_io_lsu_exe_0_fresp_bits_uop_ppred),
    .io_lsu_exe_0_fresp_bits_uop_prs1_busy(core_io_lsu_exe_0_fresp_bits_uop_prs1_busy),
    .io_lsu_exe_0_fresp_bits_uop_prs2_busy(core_io_lsu_exe_0_fresp_bits_uop_prs2_busy),
    .io_lsu_exe_0_fresp_bits_uop_prs3_busy(core_io_lsu_exe_0_fresp_bits_uop_prs3_busy),
    .io_lsu_exe_0_fresp_bits_uop_ppred_busy(core_io_lsu_exe_0_fresp_bits_uop_ppred_busy),
    .io_lsu_exe_0_fresp_bits_uop_stale_pdst(core_io_lsu_exe_0_fresp_bits_uop_stale_pdst),
    .io_lsu_exe_0_fresp_bits_uop_exception(core_io_lsu_exe_0_fresp_bits_uop_exception),
    .io_lsu_exe_0_fresp_bits_uop_exc_cause(core_io_lsu_exe_0_fresp_bits_uop_exc_cause),
    .io_lsu_exe_0_fresp_bits_uop_bypassable(core_io_lsu_exe_0_fresp_bits_uop_bypassable),
    .io_lsu_exe_0_fresp_bits_uop_mem_cmd(core_io_lsu_exe_0_fresp_bits_uop_mem_cmd),
    .io_lsu_exe_0_fresp_bits_uop_mem_size(core_io_lsu_exe_0_fresp_bits_uop_mem_size),
    .io_lsu_exe_0_fresp_bits_uop_mem_signed(core_io_lsu_exe_0_fresp_bits_uop_mem_signed),
    .io_lsu_exe_0_fresp_bits_uop_is_fence(core_io_lsu_exe_0_fresp_bits_uop_is_fence),
    .io_lsu_exe_0_fresp_bits_uop_is_fencei(core_io_lsu_exe_0_fresp_bits_uop_is_fencei),
    .io_lsu_exe_0_fresp_bits_uop_is_amo(core_io_lsu_exe_0_fresp_bits_uop_is_amo),
    .io_lsu_exe_0_fresp_bits_uop_uses_ldq(core_io_lsu_exe_0_fresp_bits_uop_uses_ldq),
    .io_lsu_exe_0_fresp_bits_uop_uses_stq(core_io_lsu_exe_0_fresp_bits_uop_uses_stq),
    .io_lsu_exe_0_fresp_bits_uop_is_sys_pc2epc(core_io_lsu_exe_0_fresp_bits_uop_is_sys_pc2epc),
    .io_lsu_exe_0_fresp_bits_uop_is_unique(core_io_lsu_exe_0_fresp_bits_uop_is_unique),
    .io_lsu_exe_0_fresp_bits_uop_flush_on_commit(core_io_lsu_exe_0_fresp_bits_uop_flush_on_commit),
    .io_lsu_exe_0_fresp_bits_uop_ldst_is_rs1(core_io_lsu_exe_0_fresp_bits_uop_ldst_is_rs1),
    .io_lsu_exe_0_fresp_bits_uop_ldst(core_io_lsu_exe_0_fresp_bits_uop_ldst),
    .io_lsu_exe_0_fresp_bits_uop_lrs1(core_io_lsu_exe_0_fresp_bits_uop_lrs1),
    .io_lsu_exe_0_fresp_bits_uop_lrs2(core_io_lsu_exe_0_fresp_bits_uop_lrs2),
    .io_lsu_exe_0_fresp_bits_uop_lrs3(core_io_lsu_exe_0_fresp_bits_uop_lrs3),
    .io_lsu_exe_0_fresp_bits_uop_ldst_val(core_io_lsu_exe_0_fresp_bits_uop_ldst_val),
    .io_lsu_exe_0_fresp_bits_uop_dst_rtype(core_io_lsu_exe_0_fresp_bits_uop_dst_rtype),
    .io_lsu_exe_0_fresp_bits_uop_lrs1_rtype(core_io_lsu_exe_0_fresp_bits_uop_lrs1_rtype),
    .io_lsu_exe_0_fresp_bits_uop_lrs2_rtype(core_io_lsu_exe_0_fresp_bits_uop_lrs2_rtype),
    .io_lsu_exe_0_fresp_bits_uop_frs3_en(core_io_lsu_exe_0_fresp_bits_uop_frs3_en),
    .io_lsu_exe_0_fresp_bits_uop_fp_val(core_io_lsu_exe_0_fresp_bits_uop_fp_val),
    .io_lsu_exe_0_fresp_bits_uop_fp_single(core_io_lsu_exe_0_fresp_bits_uop_fp_single),
    .io_lsu_exe_0_fresp_bits_uop_xcpt_pf_if(core_io_lsu_exe_0_fresp_bits_uop_xcpt_pf_if),
    .io_lsu_exe_0_fresp_bits_uop_xcpt_ae_if(core_io_lsu_exe_0_fresp_bits_uop_xcpt_ae_if),
    .io_lsu_exe_0_fresp_bits_uop_xcpt_ma_if(core_io_lsu_exe_0_fresp_bits_uop_xcpt_ma_if),
    .io_lsu_exe_0_fresp_bits_uop_bp_debug_if(core_io_lsu_exe_0_fresp_bits_uop_bp_debug_if),
    .io_lsu_exe_0_fresp_bits_uop_bp_xcpt_if(core_io_lsu_exe_0_fresp_bits_uop_bp_xcpt_if),
    .io_lsu_exe_0_fresp_bits_uop_debug_fsrc(core_io_lsu_exe_0_fresp_bits_uop_debug_fsrc),
    .io_lsu_exe_0_fresp_bits_uop_debug_tsrc(core_io_lsu_exe_0_fresp_bits_uop_debug_tsrc),
    .io_lsu_exe_0_fresp_bits_data(core_io_lsu_exe_0_fresp_bits_data),
    .io_lsu_exe_0_fresp_bits_predicated(core_io_lsu_exe_0_fresp_bits_predicated),
    .io_lsu_exe_0_fresp_bits_fflags_valid(core_io_lsu_exe_0_fresp_bits_fflags_valid),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_switch(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_switch),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_switch_off(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_switch_off),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_unicore(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_unicore),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_shift(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_shift),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs3_rtype(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs3_rtype),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_rflag(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_rflag),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_wflag(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_wflag),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_prflag(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_prflag),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_pwflag(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_pwflag),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_pflag_busy(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_pflag_busy),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_stale_pflag(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_stale_pflag),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_op1_sel(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_op1_sel),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_op2_sel(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_op2_sel),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_split_num(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_split_num),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_self_index(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_self_index),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_rob_inst_idx(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_rob_inst_idx),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_address_num(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_address_num),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_uopc(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_uopc),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_inst(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_inst),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_debug_inst(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_debug_inst),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_rvc(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_rvc),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_debug_pc(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_debug_pc),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_iq_type(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_iq_type),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_fu_code(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_fu_code),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_br_type(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_br_type),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_op1_sel(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_op1_sel),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_op2_sel(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_op2_sel),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_imm_sel(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_imm_sel),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_op_fcn(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_op_fcn),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_fcn_dw(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_fcn_dw),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_csr_cmd(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_csr_cmd),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_load(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_load),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_sta(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_sta),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_std(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_std),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_op3_sel(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_op3_sel),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_iw_state(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_iw_state),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_iw_p1_poisoned(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_iw_p1_poisoned)
      ,
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_iw_p2_poisoned(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_iw_p2_poisoned)
      ,
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_br(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_br),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_jalr(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_jalr),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_jal(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_jal),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_sfb(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_sfb),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_br_mask(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_br_mask),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_br_tag(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_br_tag),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_ftq_idx(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ftq_idx),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_edge_inst(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_edge_inst),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_pc_lob(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_pc_lob),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_taken(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_taken),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_imm_packed(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_imm_packed),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_csr_addr(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_csr_addr),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_rob_idx(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_rob_idx),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_ldq_idx(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ldq_idx),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_stq_idx(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_stq_idx),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_rxq_idx(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_rxq_idx),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_pdst(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_pdst),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs1(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs1),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs2(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs2),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs3(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs3),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_ppred(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ppred),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs1_busy(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs1_busy),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs2_busy(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs2_busy),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs3_busy(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs3_busy),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_ppred_busy(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ppred_busy),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_stale_pdst(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_stale_pdst),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_exception(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_exception),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_exc_cause(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_exc_cause),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_bypassable(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_bypassable),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_mem_cmd(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_mem_cmd),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_mem_size(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_mem_size),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_mem_signed(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_mem_signed),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_fence(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_fence),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_fencei(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_fencei),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_amo(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_amo),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_uses_ldq(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_uses_ldq),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_uses_stq(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_uses_stq),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_sys_pc2epc(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_sys_pc2epc),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_unique(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_unique),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_flush_on_commit(
      core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_flush_on_commit),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_ldst_is_rs1(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ldst_is_rs1),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_ldst(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ldst),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs1(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs1),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs2(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs2),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs3(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs3),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_ldst_val(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ldst_val),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_dst_rtype(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_dst_rtype),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs1_rtype(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs1_rtype),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs2_rtype(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs2_rtype),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_frs3_en(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_frs3_en),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_fp_val(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_fp_val),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_fp_single(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_fp_single),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_xcpt_pf_if(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_xcpt_pf_if),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_xcpt_ae_if(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_xcpt_ae_if),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_xcpt_ma_if(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_xcpt_ma_if),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_bp_debug_if(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_bp_debug_if),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_bp_xcpt_if(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_bp_xcpt_if),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_debug_fsrc(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_debug_fsrc),
    .io_lsu_exe_0_fresp_bits_fflags_bits_uop_debug_tsrc(core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_debug_tsrc),
    .io_lsu_exe_0_fresp_bits_fflags_bits_flags(core_io_lsu_exe_0_fresp_bits_fflags_bits_flags),
    .io_lsu_exe_0_fresp_bits_flagdata(core_io_lsu_exe_0_fresp_bits_flagdata),
    .io_lsu_exe_0_fresp_bits_fflagdata_valid(core_io_lsu_exe_0_fresp_bits_fflagdata_valid),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_switch(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_switch),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_switch_off(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_switch_off),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_unicore(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_unicore),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_shift(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_shift),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs3_rtype(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs3_rtype),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_rflag(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_rflag),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_wflag(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_wflag),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prflag(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prflag),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_pwflag(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_pwflag),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_pflag_busy(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_pflag_busy),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_stale_pflag(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_stale_pflag)
      ,
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_op1_sel(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_op1_sel),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_op2_sel(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_op2_sel),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_split_num(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_split_num),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_self_index(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_self_index),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_rob_inst_idx(
      core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_rob_inst_idx),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_address_num(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_address_num)
      ,
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_uopc(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_uopc),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_inst(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_inst),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_debug_inst(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_debug_inst),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_rvc(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_rvc),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_debug_pc(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_debug_pc),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_iq_type(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_iq_type),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_fu_code(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_fu_code),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_br_type(
      core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_br_type),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op1_sel(
      core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op1_sel),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op2_sel(
      core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op2_sel),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_imm_sel(
      core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_imm_sel),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op_fcn(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op_fcn)
      ,
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_fcn_dw(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_fcn_dw)
      ,
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_csr_cmd(
      core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_csr_cmd),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_load(
      core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_load),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_sta(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_sta)
      ,
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_std(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_std)
      ,
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op3_sel(
      core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op3_sel),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_iw_state(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_iw_state),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_iw_p1_poisoned(
      core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_iw_p1_poisoned),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_iw_p2_poisoned(
      core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_iw_p2_poisoned),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_br(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_br),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_jalr(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_jalr),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_jal(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_jal),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_sfb(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_sfb),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_br_mask(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_br_mask),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_br_tag(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_br_tag),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ftq_idx(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ftq_idx),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_edge_inst(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_edge_inst),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_pc_lob(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_pc_lob),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_taken(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_taken),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_imm_packed(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_imm_packed),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_csr_addr(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_csr_addr),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_rob_idx(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_rob_idx),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ldq_idx(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ldq_idx),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_stq_idx(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_stq_idx),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_rxq_idx(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_rxq_idx),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_pdst(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_pdst),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs1(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs1),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs2(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs2),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs3(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs3),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ppred(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ppred),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs1_busy(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs1_busy),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs2_busy(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs2_busy),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs3_busy(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs3_busy),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ppred_busy(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ppred_busy),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_stale_pdst(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_stale_pdst),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_exception(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_exception),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_exc_cause(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_exc_cause),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_bypassable(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_bypassable),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_mem_cmd(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_mem_cmd),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_mem_size(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_mem_size),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_mem_signed(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_mem_signed),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_fence(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_fence),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_fencei(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_fencei),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_amo(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_amo),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_uses_ldq(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_uses_ldq),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_uses_stq(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_uses_stq),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_sys_pc2epc(
      core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_sys_pc2epc),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_unique(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_unique),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_flush_on_commit(
      core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_flush_on_commit),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ldst_is_rs1(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ldst_is_rs1)
      ,
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ldst(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ldst),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs1(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs1),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs2(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs2),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs3(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs3),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ldst_val(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ldst_val),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_dst_rtype(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_dst_rtype),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs1_rtype(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs1_rtype),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs2_rtype(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs2_rtype),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_frs3_en(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_frs3_en),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_fp_val(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_fp_val),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_fp_single(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_fp_single),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_pf_if(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_pf_if),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_ae_if(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_ae_if),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_ma_if(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_ma_if),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_bp_debug_if(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_bp_debug_if)
      ,
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_bp_xcpt_if(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_bp_xcpt_if),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_debug_fsrc(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_debug_fsrc),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_debug_tsrc(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_debug_tsrc),
    .io_lsu_exe_0_fresp_bits_fflagdata_bits_fflag(core_io_lsu_exe_0_fresp_bits_fflagdata_bits_fflag),
    .io_lsu_dis_uops_0_valid(core_io_lsu_dis_uops_0_valid),
    .io_lsu_dis_uops_0_bits_switch(core_io_lsu_dis_uops_0_bits_switch),
    .io_lsu_dis_uops_0_bits_switch_off(core_io_lsu_dis_uops_0_bits_switch_off),
    .io_lsu_dis_uops_0_bits_is_unicore(core_io_lsu_dis_uops_0_bits_is_unicore),
    .io_lsu_dis_uops_0_bits_shift(core_io_lsu_dis_uops_0_bits_shift),
    .io_lsu_dis_uops_0_bits_lrs3_rtype(core_io_lsu_dis_uops_0_bits_lrs3_rtype),
    .io_lsu_dis_uops_0_bits_rflag(core_io_lsu_dis_uops_0_bits_rflag),
    .io_lsu_dis_uops_0_bits_wflag(core_io_lsu_dis_uops_0_bits_wflag),
    .io_lsu_dis_uops_0_bits_prflag(core_io_lsu_dis_uops_0_bits_prflag),
    .io_lsu_dis_uops_0_bits_pwflag(core_io_lsu_dis_uops_0_bits_pwflag),
    .io_lsu_dis_uops_0_bits_pflag_busy(core_io_lsu_dis_uops_0_bits_pflag_busy),
    .io_lsu_dis_uops_0_bits_stale_pflag(core_io_lsu_dis_uops_0_bits_stale_pflag),
    .io_lsu_dis_uops_0_bits_op1_sel(core_io_lsu_dis_uops_0_bits_op1_sel),
    .io_lsu_dis_uops_0_bits_op2_sel(core_io_lsu_dis_uops_0_bits_op2_sel),
    .io_lsu_dis_uops_0_bits_split_num(core_io_lsu_dis_uops_0_bits_split_num),
    .io_lsu_dis_uops_0_bits_self_index(core_io_lsu_dis_uops_0_bits_self_index),
    .io_lsu_dis_uops_0_bits_rob_inst_idx(core_io_lsu_dis_uops_0_bits_rob_inst_idx),
    .io_lsu_dis_uops_0_bits_address_num(core_io_lsu_dis_uops_0_bits_address_num),
    .io_lsu_dis_uops_0_bits_uopc(core_io_lsu_dis_uops_0_bits_uopc),
    .io_lsu_dis_uops_0_bits_inst(core_io_lsu_dis_uops_0_bits_inst),
    .io_lsu_dis_uops_0_bits_debug_inst(core_io_lsu_dis_uops_0_bits_debug_inst),
    .io_lsu_dis_uops_0_bits_is_rvc(core_io_lsu_dis_uops_0_bits_is_rvc),
    .io_lsu_dis_uops_0_bits_debug_pc(core_io_lsu_dis_uops_0_bits_debug_pc),
    .io_lsu_dis_uops_0_bits_iq_type(core_io_lsu_dis_uops_0_bits_iq_type),
    .io_lsu_dis_uops_0_bits_fu_code(core_io_lsu_dis_uops_0_bits_fu_code),
    .io_lsu_dis_uops_0_bits_ctrl_br_type(core_io_lsu_dis_uops_0_bits_ctrl_br_type),
    .io_lsu_dis_uops_0_bits_ctrl_op1_sel(core_io_lsu_dis_uops_0_bits_ctrl_op1_sel),
    .io_lsu_dis_uops_0_bits_ctrl_op2_sel(core_io_lsu_dis_uops_0_bits_ctrl_op2_sel),
    .io_lsu_dis_uops_0_bits_ctrl_imm_sel(core_io_lsu_dis_uops_0_bits_ctrl_imm_sel),
    .io_lsu_dis_uops_0_bits_ctrl_op_fcn(core_io_lsu_dis_uops_0_bits_ctrl_op_fcn),
    .io_lsu_dis_uops_0_bits_ctrl_fcn_dw(core_io_lsu_dis_uops_0_bits_ctrl_fcn_dw),
    .io_lsu_dis_uops_0_bits_ctrl_csr_cmd(core_io_lsu_dis_uops_0_bits_ctrl_csr_cmd),
    .io_lsu_dis_uops_0_bits_ctrl_is_load(core_io_lsu_dis_uops_0_bits_ctrl_is_load),
    .io_lsu_dis_uops_0_bits_ctrl_is_sta(core_io_lsu_dis_uops_0_bits_ctrl_is_sta),
    .io_lsu_dis_uops_0_bits_ctrl_is_std(core_io_lsu_dis_uops_0_bits_ctrl_is_std),
    .io_lsu_dis_uops_0_bits_ctrl_op3_sel(core_io_lsu_dis_uops_0_bits_ctrl_op3_sel),
    .io_lsu_dis_uops_0_bits_iw_state(core_io_lsu_dis_uops_0_bits_iw_state),
    .io_lsu_dis_uops_0_bits_iw_p1_poisoned(core_io_lsu_dis_uops_0_bits_iw_p1_poisoned),
    .io_lsu_dis_uops_0_bits_iw_p2_poisoned(core_io_lsu_dis_uops_0_bits_iw_p2_poisoned),
    .io_lsu_dis_uops_0_bits_is_br(core_io_lsu_dis_uops_0_bits_is_br),
    .io_lsu_dis_uops_0_bits_is_jalr(core_io_lsu_dis_uops_0_bits_is_jalr),
    .io_lsu_dis_uops_0_bits_is_jal(core_io_lsu_dis_uops_0_bits_is_jal),
    .io_lsu_dis_uops_0_bits_is_sfb(core_io_lsu_dis_uops_0_bits_is_sfb),
    .io_lsu_dis_uops_0_bits_br_mask(core_io_lsu_dis_uops_0_bits_br_mask),
    .io_lsu_dis_uops_0_bits_br_tag(core_io_lsu_dis_uops_0_bits_br_tag),
    .io_lsu_dis_uops_0_bits_ftq_idx(core_io_lsu_dis_uops_0_bits_ftq_idx),
    .io_lsu_dis_uops_0_bits_edge_inst(core_io_lsu_dis_uops_0_bits_edge_inst),
    .io_lsu_dis_uops_0_bits_pc_lob(core_io_lsu_dis_uops_0_bits_pc_lob),
    .io_lsu_dis_uops_0_bits_taken(core_io_lsu_dis_uops_0_bits_taken),
    .io_lsu_dis_uops_0_bits_imm_packed(core_io_lsu_dis_uops_0_bits_imm_packed),
    .io_lsu_dis_uops_0_bits_csr_addr(core_io_lsu_dis_uops_0_bits_csr_addr),
    .io_lsu_dis_uops_0_bits_rob_idx(core_io_lsu_dis_uops_0_bits_rob_idx),
    .io_lsu_dis_uops_0_bits_ldq_idx(core_io_lsu_dis_uops_0_bits_ldq_idx),
    .io_lsu_dis_uops_0_bits_stq_idx(core_io_lsu_dis_uops_0_bits_stq_idx),
    .io_lsu_dis_uops_0_bits_rxq_idx(core_io_lsu_dis_uops_0_bits_rxq_idx),
    .io_lsu_dis_uops_0_bits_pdst(core_io_lsu_dis_uops_0_bits_pdst),
    .io_lsu_dis_uops_0_bits_prs1(core_io_lsu_dis_uops_0_bits_prs1),
    .io_lsu_dis_uops_0_bits_prs2(core_io_lsu_dis_uops_0_bits_prs2),
    .io_lsu_dis_uops_0_bits_prs3(core_io_lsu_dis_uops_0_bits_prs3),
    .io_lsu_dis_uops_0_bits_ppred(core_io_lsu_dis_uops_0_bits_ppred),
    .io_lsu_dis_uops_0_bits_prs1_busy(core_io_lsu_dis_uops_0_bits_prs1_busy),
    .io_lsu_dis_uops_0_bits_prs2_busy(core_io_lsu_dis_uops_0_bits_prs2_busy),
    .io_lsu_dis_uops_0_bits_prs3_busy(core_io_lsu_dis_uops_0_bits_prs3_busy),
    .io_lsu_dis_uops_0_bits_ppred_busy(core_io_lsu_dis_uops_0_bits_ppred_busy),
    .io_lsu_dis_uops_0_bits_stale_pdst(core_io_lsu_dis_uops_0_bits_stale_pdst),
    .io_lsu_dis_uops_0_bits_exception(core_io_lsu_dis_uops_0_bits_exception),
    .io_lsu_dis_uops_0_bits_exc_cause(core_io_lsu_dis_uops_0_bits_exc_cause),
    .io_lsu_dis_uops_0_bits_bypassable(core_io_lsu_dis_uops_0_bits_bypassable),
    .io_lsu_dis_uops_0_bits_mem_cmd(core_io_lsu_dis_uops_0_bits_mem_cmd),
    .io_lsu_dis_uops_0_bits_mem_size(core_io_lsu_dis_uops_0_bits_mem_size),
    .io_lsu_dis_uops_0_bits_mem_signed(core_io_lsu_dis_uops_0_bits_mem_signed),
    .io_lsu_dis_uops_0_bits_is_fence(core_io_lsu_dis_uops_0_bits_is_fence),
    .io_lsu_dis_uops_0_bits_is_fencei(core_io_lsu_dis_uops_0_bits_is_fencei),
    .io_lsu_dis_uops_0_bits_is_amo(core_io_lsu_dis_uops_0_bits_is_amo),
    .io_lsu_dis_uops_0_bits_uses_ldq(core_io_lsu_dis_uops_0_bits_uses_ldq),
    .io_lsu_dis_uops_0_bits_uses_stq(core_io_lsu_dis_uops_0_bits_uses_stq),
    .io_lsu_dis_uops_0_bits_is_sys_pc2epc(core_io_lsu_dis_uops_0_bits_is_sys_pc2epc),
    .io_lsu_dis_uops_0_bits_is_unique(core_io_lsu_dis_uops_0_bits_is_unique),
    .io_lsu_dis_uops_0_bits_flush_on_commit(core_io_lsu_dis_uops_0_bits_flush_on_commit),
    .io_lsu_dis_uops_0_bits_ldst_is_rs1(core_io_lsu_dis_uops_0_bits_ldst_is_rs1),
    .io_lsu_dis_uops_0_bits_ldst(core_io_lsu_dis_uops_0_bits_ldst),
    .io_lsu_dis_uops_0_bits_lrs1(core_io_lsu_dis_uops_0_bits_lrs1),
    .io_lsu_dis_uops_0_bits_lrs2(core_io_lsu_dis_uops_0_bits_lrs2),
    .io_lsu_dis_uops_0_bits_lrs3(core_io_lsu_dis_uops_0_bits_lrs3),
    .io_lsu_dis_uops_0_bits_ldst_val(core_io_lsu_dis_uops_0_bits_ldst_val),
    .io_lsu_dis_uops_0_bits_dst_rtype(core_io_lsu_dis_uops_0_bits_dst_rtype),
    .io_lsu_dis_uops_0_bits_lrs1_rtype(core_io_lsu_dis_uops_0_bits_lrs1_rtype),
    .io_lsu_dis_uops_0_bits_lrs2_rtype(core_io_lsu_dis_uops_0_bits_lrs2_rtype),
    .io_lsu_dis_uops_0_bits_frs3_en(core_io_lsu_dis_uops_0_bits_frs3_en),
    .io_lsu_dis_uops_0_bits_fp_val(core_io_lsu_dis_uops_0_bits_fp_val),
    .io_lsu_dis_uops_0_bits_fp_single(core_io_lsu_dis_uops_0_bits_fp_single),
    .io_lsu_dis_uops_0_bits_xcpt_pf_if(core_io_lsu_dis_uops_0_bits_xcpt_pf_if),
    .io_lsu_dis_uops_0_bits_xcpt_ae_if(core_io_lsu_dis_uops_0_bits_xcpt_ae_if),
    .io_lsu_dis_uops_0_bits_xcpt_ma_if(core_io_lsu_dis_uops_0_bits_xcpt_ma_if),
    .io_lsu_dis_uops_0_bits_bp_debug_if(core_io_lsu_dis_uops_0_bits_bp_debug_if),
    .io_lsu_dis_uops_0_bits_bp_xcpt_if(core_io_lsu_dis_uops_0_bits_bp_xcpt_if),
    .io_lsu_dis_uops_0_bits_debug_fsrc(core_io_lsu_dis_uops_0_bits_debug_fsrc),
    .io_lsu_dis_uops_0_bits_debug_tsrc(core_io_lsu_dis_uops_0_bits_debug_tsrc),
    .io_lsu_dis_uops_1_valid(core_io_lsu_dis_uops_1_valid),
    .io_lsu_dis_uops_1_bits_switch(core_io_lsu_dis_uops_1_bits_switch),
    .io_lsu_dis_uops_1_bits_switch_off(core_io_lsu_dis_uops_1_bits_switch_off),
    .io_lsu_dis_uops_1_bits_is_unicore(core_io_lsu_dis_uops_1_bits_is_unicore),
    .io_lsu_dis_uops_1_bits_shift(core_io_lsu_dis_uops_1_bits_shift),
    .io_lsu_dis_uops_1_bits_lrs3_rtype(core_io_lsu_dis_uops_1_bits_lrs3_rtype),
    .io_lsu_dis_uops_1_bits_rflag(core_io_lsu_dis_uops_1_bits_rflag),
    .io_lsu_dis_uops_1_bits_wflag(core_io_lsu_dis_uops_1_bits_wflag),
    .io_lsu_dis_uops_1_bits_prflag(core_io_lsu_dis_uops_1_bits_prflag),
    .io_lsu_dis_uops_1_bits_pwflag(core_io_lsu_dis_uops_1_bits_pwflag),
    .io_lsu_dis_uops_1_bits_pflag_busy(core_io_lsu_dis_uops_1_bits_pflag_busy),
    .io_lsu_dis_uops_1_bits_stale_pflag(core_io_lsu_dis_uops_1_bits_stale_pflag),
    .io_lsu_dis_uops_1_bits_op1_sel(core_io_lsu_dis_uops_1_bits_op1_sel),
    .io_lsu_dis_uops_1_bits_op2_sel(core_io_lsu_dis_uops_1_bits_op2_sel),
    .io_lsu_dis_uops_1_bits_split_num(core_io_lsu_dis_uops_1_bits_split_num),
    .io_lsu_dis_uops_1_bits_self_index(core_io_lsu_dis_uops_1_bits_self_index),
    .io_lsu_dis_uops_1_bits_rob_inst_idx(core_io_lsu_dis_uops_1_bits_rob_inst_idx),
    .io_lsu_dis_uops_1_bits_address_num(core_io_lsu_dis_uops_1_bits_address_num),
    .io_lsu_dis_uops_1_bits_uopc(core_io_lsu_dis_uops_1_bits_uopc),
    .io_lsu_dis_uops_1_bits_inst(core_io_lsu_dis_uops_1_bits_inst),
    .io_lsu_dis_uops_1_bits_debug_inst(core_io_lsu_dis_uops_1_bits_debug_inst),
    .io_lsu_dis_uops_1_bits_is_rvc(core_io_lsu_dis_uops_1_bits_is_rvc),
    .io_lsu_dis_uops_1_bits_debug_pc(core_io_lsu_dis_uops_1_bits_debug_pc),
    .io_lsu_dis_uops_1_bits_iq_type(core_io_lsu_dis_uops_1_bits_iq_type),
    .io_lsu_dis_uops_1_bits_fu_code(core_io_lsu_dis_uops_1_bits_fu_code),
    .io_lsu_dis_uops_1_bits_ctrl_br_type(core_io_lsu_dis_uops_1_bits_ctrl_br_type),
    .io_lsu_dis_uops_1_bits_ctrl_op1_sel(core_io_lsu_dis_uops_1_bits_ctrl_op1_sel),
    .io_lsu_dis_uops_1_bits_ctrl_op2_sel(core_io_lsu_dis_uops_1_bits_ctrl_op2_sel),
    .io_lsu_dis_uops_1_bits_ctrl_imm_sel(core_io_lsu_dis_uops_1_bits_ctrl_imm_sel),
    .io_lsu_dis_uops_1_bits_ctrl_op_fcn(core_io_lsu_dis_uops_1_bits_ctrl_op_fcn),
    .io_lsu_dis_uops_1_bits_ctrl_fcn_dw(core_io_lsu_dis_uops_1_bits_ctrl_fcn_dw),
    .io_lsu_dis_uops_1_bits_ctrl_csr_cmd(core_io_lsu_dis_uops_1_bits_ctrl_csr_cmd),
    .io_lsu_dis_uops_1_bits_ctrl_is_load(core_io_lsu_dis_uops_1_bits_ctrl_is_load),
    .io_lsu_dis_uops_1_bits_ctrl_is_sta(core_io_lsu_dis_uops_1_bits_ctrl_is_sta),
    .io_lsu_dis_uops_1_bits_ctrl_is_std(core_io_lsu_dis_uops_1_bits_ctrl_is_std),
    .io_lsu_dis_uops_1_bits_ctrl_op3_sel(core_io_lsu_dis_uops_1_bits_ctrl_op3_sel),
    .io_lsu_dis_uops_1_bits_iw_state(core_io_lsu_dis_uops_1_bits_iw_state),
    .io_lsu_dis_uops_1_bits_iw_p1_poisoned(core_io_lsu_dis_uops_1_bits_iw_p1_poisoned),
    .io_lsu_dis_uops_1_bits_iw_p2_poisoned(core_io_lsu_dis_uops_1_bits_iw_p2_poisoned),
    .io_lsu_dis_uops_1_bits_is_br(core_io_lsu_dis_uops_1_bits_is_br),
    .io_lsu_dis_uops_1_bits_is_jalr(core_io_lsu_dis_uops_1_bits_is_jalr),
    .io_lsu_dis_uops_1_bits_is_jal(core_io_lsu_dis_uops_1_bits_is_jal),
    .io_lsu_dis_uops_1_bits_is_sfb(core_io_lsu_dis_uops_1_bits_is_sfb),
    .io_lsu_dis_uops_1_bits_br_mask(core_io_lsu_dis_uops_1_bits_br_mask),
    .io_lsu_dis_uops_1_bits_br_tag(core_io_lsu_dis_uops_1_bits_br_tag),
    .io_lsu_dis_uops_1_bits_ftq_idx(core_io_lsu_dis_uops_1_bits_ftq_idx),
    .io_lsu_dis_uops_1_bits_edge_inst(core_io_lsu_dis_uops_1_bits_edge_inst),
    .io_lsu_dis_uops_1_bits_pc_lob(core_io_lsu_dis_uops_1_bits_pc_lob),
    .io_lsu_dis_uops_1_bits_taken(core_io_lsu_dis_uops_1_bits_taken),
    .io_lsu_dis_uops_1_bits_imm_packed(core_io_lsu_dis_uops_1_bits_imm_packed),
    .io_lsu_dis_uops_1_bits_csr_addr(core_io_lsu_dis_uops_1_bits_csr_addr),
    .io_lsu_dis_uops_1_bits_rob_idx(core_io_lsu_dis_uops_1_bits_rob_idx),
    .io_lsu_dis_uops_1_bits_ldq_idx(core_io_lsu_dis_uops_1_bits_ldq_idx),
    .io_lsu_dis_uops_1_bits_stq_idx(core_io_lsu_dis_uops_1_bits_stq_idx),
    .io_lsu_dis_uops_1_bits_rxq_idx(core_io_lsu_dis_uops_1_bits_rxq_idx),
    .io_lsu_dis_uops_1_bits_pdst(core_io_lsu_dis_uops_1_bits_pdst),
    .io_lsu_dis_uops_1_bits_prs1(core_io_lsu_dis_uops_1_bits_prs1),
    .io_lsu_dis_uops_1_bits_prs2(core_io_lsu_dis_uops_1_bits_prs2),
    .io_lsu_dis_uops_1_bits_prs3(core_io_lsu_dis_uops_1_bits_prs3),
    .io_lsu_dis_uops_1_bits_ppred(core_io_lsu_dis_uops_1_bits_ppred),
    .io_lsu_dis_uops_1_bits_prs1_busy(core_io_lsu_dis_uops_1_bits_prs1_busy),
    .io_lsu_dis_uops_1_bits_prs2_busy(core_io_lsu_dis_uops_1_bits_prs2_busy),
    .io_lsu_dis_uops_1_bits_prs3_busy(core_io_lsu_dis_uops_1_bits_prs3_busy),
    .io_lsu_dis_uops_1_bits_ppred_busy(core_io_lsu_dis_uops_1_bits_ppred_busy),
    .io_lsu_dis_uops_1_bits_stale_pdst(core_io_lsu_dis_uops_1_bits_stale_pdst),
    .io_lsu_dis_uops_1_bits_exception(core_io_lsu_dis_uops_1_bits_exception),
    .io_lsu_dis_uops_1_bits_exc_cause(core_io_lsu_dis_uops_1_bits_exc_cause),
    .io_lsu_dis_uops_1_bits_bypassable(core_io_lsu_dis_uops_1_bits_bypassable),
    .io_lsu_dis_uops_1_bits_mem_cmd(core_io_lsu_dis_uops_1_bits_mem_cmd),
    .io_lsu_dis_uops_1_bits_mem_size(core_io_lsu_dis_uops_1_bits_mem_size),
    .io_lsu_dis_uops_1_bits_mem_signed(core_io_lsu_dis_uops_1_bits_mem_signed),
    .io_lsu_dis_uops_1_bits_is_fence(core_io_lsu_dis_uops_1_bits_is_fence),
    .io_lsu_dis_uops_1_bits_is_fencei(core_io_lsu_dis_uops_1_bits_is_fencei),
    .io_lsu_dis_uops_1_bits_is_amo(core_io_lsu_dis_uops_1_bits_is_amo),
    .io_lsu_dis_uops_1_bits_uses_ldq(core_io_lsu_dis_uops_1_bits_uses_ldq),
    .io_lsu_dis_uops_1_bits_uses_stq(core_io_lsu_dis_uops_1_bits_uses_stq),
    .io_lsu_dis_uops_1_bits_is_sys_pc2epc(core_io_lsu_dis_uops_1_bits_is_sys_pc2epc),
    .io_lsu_dis_uops_1_bits_is_unique(core_io_lsu_dis_uops_1_bits_is_unique),
    .io_lsu_dis_uops_1_bits_flush_on_commit(core_io_lsu_dis_uops_1_bits_flush_on_commit),
    .io_lsu_dis_uops_1_bits_ldst_is_rs1(core_io_lsu_dis_uops_1_bits_ldst_is_rs1),
    .io_lsu_dis_uops_1_bits_ldst(core_io_lsu_dis_uops_1_bits_ldst),
    .io_lsu_dis_uops_1_bits_lrs1(core_io_lsu_dis_uops_1_bits_lrs1),
    .io_lsu_dis_uops_1_bits_lrs2(core_io_lsu_dis_uops_1_bits_lrs2),
    .io_lsu_dis_uops_1_bits_lrs3(core_io_lsu_dis_uops_1_bits_lrs3),
    .io_lsu_dis_uops_1_bits_ldst_val(core_io_lsu_dis_uops_1_bits_ldst_val),
    .io_lsu_dis_uops_1_bits_dst_rtype(core_io_lsu_dis_uops_1_bits_dst_rtype),
    .io_lsu_dis_uops_1_bits_lrs1_rtype(core_io_lsu_dis_uops_1_bits_lrs1_rtype),
    .io_lsu_dis_uops_1_bits_lrs2_rtype(core_io_lsu_dis_uops_1_bits_lrs2_rtype),
    .io_lsu_dis_uops_1_bits_frs3_en(core_io_lsu_dis_uops_1_bits_frs3_en),
    .io_lsu_dis_uops_1_bits_fp_val(core_io_lsu_dis_uops_1_bits_fp_val),
    .io_lsu_dis_uops_1_bits_fp_single(core_io_lsu_dis_uops_1_bits_fp_single),
    .io_lsu_dis_uops_1_bits_xcpt_pf_if(core_io_lsu_dis_uops_1_bits_xcpt_pf_if),
    .io_lsu_dis_uops_1_bits_xcpt_ae_if(core_io_lsu_dis_uops_1_bits_xcpt_ae_if),
    .io_lsu_dis_uops_1_bits_xcpt_ma_if(core_io_lsu_dis_uops_1_bits_xcpt_ma_if),
    .io_lsu_dis_uops_1_bits_bp_debug_if(core_io_lsu_dis_uops_1_bits_bp_debug_if),
    .io_lsu_dis_uops_1_bits_bp_xcpt_if(core_io_lsu_dis_uops_1_bits_bp_xcpt_if),
    .io_lsu_dis_uops_1_bits_debug_fsrc(core_io_lsu_dis_uops_1_bits_debug_fsrc),
    .io_lsu_dis_uops_1_bits_debug_tsrc(core_io_lsu_dis_uops_1_bits_debug_tsrc),
    .io_lsu_dis_ldq_idx_0(core_io_lsu_dis_ldq_idx_0),
    .io_lsu_dis_ldq_idx_1(core_io_lsu_dis_ldq_idx_1),
    .io_lsu_dis_stq_idx_0(core_io_lsu_dis_stq_idx_0),
    .io_lsu_dis_stq_idx_1(core_io_lsu_dis_stq_idx_1),
    .io_lsu_ldq_full_0(core_io_lsu_ldq_full_0),
    .io_lsu_ldq_full_1(core_io_lsu_ldq_full_1),
    .io_lsu_stq_full_0(core_io_lsu_stq_full_0),
    .io_lsu_stq_full_1(core_io_lsu_stq_full_1),
    .io_lsu_fp_stdata_ready(core_io_lsu_fp_stdata_ready),
    .io_lsu_fp_stdata_valid(core_io_lsu_fp_stdata_valid),
    .io_lsu_fp_stdata_bits_uop_switch(core_io_lsu_fp_stdata_bits_uop_switch),
    .io_lsu_fp_stdata_bits_uop_switch_off(core_io_lsu_fp_stdata_bits_uop_switch_off),
    .io_lsu_fp_stdata_bits_uop_is_unicore(core_io_lsu_fp_stdata_bits_uop_is_unicore),
    .io_lsu_fp_stdata_bits_uop_shift(core_io_lsu_fp_stdata_bits_uop_shift),
    .io_lsu_fp_stdata_bits_uop_lrs3_rtype(core_io_lsu_fp_stdata_bits_uop_lrs3_rtype),
    .io_lsu_fp_stdata_bits_uop_rflag(core_io_lsu_fp_stdata_bits_uop_rflag),
    .io_lsu_fp_stdata_bits_uop_wflag(core_io_lsu_fp_stdata_bits_uop_wflag),
    .io_lsu_fp_stdata_bits_uop_prflag(core_io_lsu_fp_stdata_bits_uop_prflag),
    .io_lsu_fp_stdata_bits_uop_pwflag(core_io_lsu_fp_stdata_bits_uop_pwflag),
    .io_lsu_fp_stdata_bits_uop_pflag_busy(core_io_lsu_fp_stdata_bits_uop_pflag_busy),
    .io_lsu_fp_stdata_bits_uop_stale_pflag(core_io_lsu_fp_stdata_bits_uop_stale_pflag),
    .io_lsu_fp_stdata_bits_uop_op1_sel(core_io_lsu_fp_stdata_bits_uop_op1_sel),
    .io_lsu_fp_stdata_bits_uop_op2_sel(core_io_lsu_fp_stdata_bits_uop_op2_sel),
    .io_lsu_fp_stdata_bits_uop_split_num(core_io_lsu_fp_stdata_bits_uop_split_num),
    .io_lsu_fp_stdata_bits_uop_self_index(core_io_lsu_fp_stdata_bits_uop_self_index),
    .io_lsu_fp_stdata_bits_uop_rob_inst_idx(core_io_lsu_fp_stdata_bits_uop_rob_inst_idx),
    .io_lsu_fp_stdata_bits_uop_address_num(core_io_lsu_fp_stdata_bits_uop_address_num),
    .io_lsu_fp_stdata_bits_uop_uopc(core_io_lsu_fp_stdata_bits_uop_uopc),
    .io_lsu_fp_stdata_bits_uop_inst(core_io_lsu_fp_stdata_bits_uop_inst),
    .io_lsu_fp_stdata_bits_uop_debug_inst(core_io_lsu_fp_stdata_bits_uop_debug_inst),
    .io_lsu_fp_stdata_bits_uop_is_rvc(core_io_lsu_fp_stdata_bits_uop_is_rvc),
    .io_lsu_fp_stdata_bits_uop_debug_pc(core_io_lsu_fp_stdata_bits_uop_debug_pc),
    .io_lsu_fp_stdata_bits_uop_iq_type(core_io_lsu_fp_stdata_bits_uop_iq_type),
    .io_lsu_fp_stdata_bits_uop_fu_code(core_io_lsu_fp_stdata_bits_uop_fu_code),
    .io_lsu_fp_stdata_bits_uop_ctrl_br_type(core_io_lsu_fp_stdata_bits_uop_ctrl_br_type),
    .io_lsu_fp_stdata_bits_uop_ctrl_op1_sel(core_io_lsu_fp_stdata_bits_uop_ctrl_op1_sel),
    .io_lsu_fp_stdata_bits_uop_ctrl_op2_sel(core_io_lsu_fp_stdata_bits_uop_ctrl_op2_sel),
    .io_lsu_fp_stdata_bits_uop_ctrl_imm_sel(core_io_lsu_fp_stdata_bits_uop_ctrl_imm_sel),
    .io_lsu_fp_stdata_bits_uop_ctrl_op_fcn(core_io_lsu_fp_stdata_bits_uop_ctrl_op_fcn),
    .io_lsu_fp_stdata_bits_uop_ctrl_fcn_dw(core_io_lsu_fp_stdata_bits_uop_ctrl_fcn_dw),
    .io_lsu_fp_stdata_bits_uop_ctrl_csr_cmd(core_io_lsu_fp_stdata_bits_uop_ctrl_csr_cmd),
    .io_lsu_fp_stdata_bits_uop_ctrl_is_load(core_io_lsu_fp_stdata_bits_uop_ctrl_is_load),
    .io_lsu_fp_stdata_bits_uop_ctrl_is_sta(core_io_lsu_fp_stdata_bits_uop_ctrl_is_sta),
    .io_lsu_fp_stdata_bits_uop_ctrl_is_std(core_io_lsu_fp_stdata_bits_uop_ctrl_is_std),
    .io_lsu_fp_stdata_bits_uop_ctrl_op3_sel(core_io_lsu_fp_stdata_bits_uop_ctrl_op3_sel),
    .io_lsu_fp_stdata_bits_uop_iw_state(core_io_lsu_fp_stdata_bits_uop_iw_state),
    .io_lsu_fp_stdata_bits_uop_iw_p1_poisoned(core_io_lsu_fp_stdata_bits_uop_iw_p1_poisoned),
    .io_lsu_fp_stdata_bits_uop_iw_p2_poisoned(core_io_lsu_fp_stdata_bits_uop_iw_p2_poisoned),
    .io_lsu_fp_stdata_bits_uop_is_br(core_io_lsu_fp_stdata_bits_uop_is_br),
    .io_lsu_fp_stdata_bits_uop_is_jalr(core_io_lsu_fp_stdata_bits_uop_is_jalr),
    .io_lsu_fp_stdata_bits_uop_is_jal(core_io_lsu_fp_stdata_bits_uop_is_jal),
    .io_lsu_fp_stdata_bits_uop_is_sfb(core_io_lsu_fp_stdata_bits_uop_is_sfb),
    .io_lsu_fp_stdata_bits_uop_br_mask(core_io_lsu_fp_stdata_bits_uop_br_mask),
    .io_lsu_fp_stdata_bits_uop_br_tag(core_io_lsu_fp_stdata_bits_uop_br_tag),
    .io_lsu_fp_stdata_bits_uop_ftq_idx(core_io_lsu_fp_stdata_bits_uop_ftq_idx),
    .io_lsu_fp_stdata_bits_uop_edge_inst(core_io_lsu_fp_stdata_bits_uop_edge_inst),
    .io_lsu_fp_stdata_bits_uop_pc_lob(core_io_lsu_fp_stdata_bits_uop_pc_lob),
    .io_lsu_fp_stdata_bits_uop_taken(core_io_lsu_fp_stdata_bits_uop_taken),
    .io_lsu_fp_stdata_bits_uop_imm_packed(core_io_lsu_fp_stdata_bits_uop_imm_packed),
    .io_lsu_fp_stdata_bits_uop_csr_addr(core_io_lsu_fp_stdata_bits_uop_csr_addr),
    .io_lsu_fp_stdata_bits_uop_rob_idx(core_io_lsu_fp_stdata_bits_uop_rob_idx),
    .io_lsu_fp_stdata_bits_uop_ldq_idx(core_io_lsu_fp_stdata_bits_uop_ldq_idx),
    .io_lsu_fp_stdata_bits_uop_stq_idx(core_io_lsu_fp_stdata_bits_uop_stq_idx),
    .io_lsu_fp_stdata_bits_uop_rxq_idx(core_io_lsu_fp_stdata_bits_uop_rxq_idx),
    .io_lsu_fp_stdata_bits_uop_pdst(core_io_lsu_fp_stdata_bits_uop_pdst),
    .io_lsu_fp_stdata_bits_uop_prs1(core_io_lsu_fp_stdata_bits_uop_prs1),
    .io_lsu_fp_stdata_bits_uop_prs2(core_io_lsu_fp_stdata_bits_uop_prs2),
    .io_lsu_fp_stdata_bits_uop_prs3(core_io_lsu_fp_stdata_bits_uop_prs3),
    .io_lsu_fp_stdata_bits_uop_ppred(core_io_lsu_fp_stdata_bits_uop_ppred),
    .io_lsu_fp_stdata_bits_uop_prs1_busy(core_io_lsu_fp_stdata_bits_uop_prs1_busy),
    .io_lsu_fp_stdata_bits_uop_prs2_busy(core_io_lsu_fp_stdata_bits_uop_prs2_busy),
    .io_lsu_fp_stdata_bits_uop_prs3_busy(core_io_lsu_fp_stdata_bits_uop_prs3_busy),
    .io_lsu_fp_stdata_bits_uop_ppred_busy(core_io_lsu_fp_stdata_bits_uop_ppred_busy),
    .io_lsu_fp_stdata_bits_uop_stale_pdst(core_io_lsu_fp_stdata_bits_uop_stale_pdst),
    .io_lsu_fp_stdata_bits_uop_exception(core_io_lsu_fp_stdata_bits_uop_exception),
    .io_lsu_fp_stdata_bits_uop_exc_cause(core_io_lsu_fp_stdata_bits_uop_exc_cause),
    .io_lsu_fp_stdata_bits_uop_bypassable(core_io_lsu_fp_stdata_bits_uop_bypassable),
    .io_lsu_fp_stdata_bits_uop_mem_cmd(core_io_lsu_fp_stdata_bits_uop_mem_cmd),
    .io_lsu_fp_stdata_bits_uop_mem_size(core_io_lsu_fp_stdata_bits_uop_mem_size),
    .io_lsu_fp_stdata_bits_uop_mem_signed(core_io_lsu_fp_stdata_bits_uop_mem_signed),
    .io_lsu_fp_stdata_bits_uop_is_fence(core_io_lsu_fp_stdata_bits_uop_is_fence),
    .io_lsu_fp_stdata_bits_uop_is_fencei(core_io_lsu_fp_stdata_bits_uop_is_fencei),
    .io_lsu_fp_stdata_bits_uop_is_amo(core_io_lsu_fp_stdata_bits_uop_is_amo),
    .io_lsu_fp_stdata_bits_uop_uses_ldq(core_io_lsu_fp_stdata_bits_uop_uses_ldq),
    .io_lsu_fp_stdata_bits_uop_uses_stq(core_io_lsu_fp_stdata_bits_uop_uses_stq),
    .io_lsu_fp_stdata_bits_uop_is_sys_pc2epc(core_io_lsu_fp_stdata_bits_uop_is_sys_pc2epc),
    .io_lsu_fp_stdata_bits_uop_is_unique(core_io_lsu_fp_stdata_bits_uop_is_unique),
    .io_lsu_fp_stdata_bits_uop_flush_on_commit(core_io_lsu_fp_stdata_bits_uop_flush_on_commit),
    .io_lsu_fp_stdata_bits_uop_ldst_is_rs1(core_io_lsu_fp_stdata_bits_uop_ldst_is_rs1),
    .io_lsu_fp_stdata_bits_uop_ldst(core_io_lsu_fp_stdata_bits_uop_ldst),
    .io_lsu_fp_stdata_bits_uop_lrs1(core_io_lsu_fp_stdata_bits_uop_lrs1),
    .io_lsu_fp_stdata_bits_uop_lrs2(core_io_lsu_fp_stdata_bits_uop_lrs2),
    .io_lsu_fp_stdata_bits_uop_lrs3(core_io_lsu_fp_stdata_bits_uop_lrs3),
    .io_lsu_fp_stdata_bits_uop_ldst_val(core_io_lsu_fp_stdata_bits_uop_ldst_val),
    .io_lsu_fp_stdata_bits_uop_dst_rtype(core_io_lsu_fp_stdata_bits_uop_dst_rtype),
    .io_lsu_fp_stdata_bits_uop_lrs1_rtype(core_io_lsu_fp_stdata_bits_uop_lrs1_rtype),
    .io_lsu_fp_stdata_bits_uop_lrs2_rtype(core_io_lsu_fp_stdata_bits_uop_lrs2_rtype),
    .io_lsu_fp_stdata_bits_uop_frs3_en(core_io_lsu_fp_stdata_bits_uop_frs3_en),
    .io_lsu_fp_stdata_bits_uop_fp_val(core_io_lsu_fp_stdata_bits_uop_fp_val),
    .io_lsu_fp_stdata_bits_uop_fp_single(core_io_lsu_fp_stdata_bits_uop_fp_single),
    .io_lsu_fp_stdata_bits_uop_xcpt_pf_if(core_io_lsu_fp_stdata_bits_uop_xcpt_pf_if),
    .io_lsu_fp_stdata_bits_uop_xcpt_ae_if(core_io_lsu_fp_stdata_bits_uop_xcpt_ae_if),
    .io_lsu_fp_stdata_bits_uop_xcpt_ma_if(core_io_lsu_fp_stdata_bits_uop_xcpt_ma_if),
    .io_lsu_fp_stdata_bits_uop_bp_debug_if(core_io_lsu_fp_stdata_bits_uop_bp_debug_if),
    .io_lsu_fp_stdata_bits_uop_bp_xcpt_if(core_io_lsu_fp_stdata_bits_uop_bp_xcpt_if),
    .io_lsu_fp_stdata_bits_uop_debug_fsrc(core_io_lsu_fp_stdata_bits_uop_debug_fsrc),
    .io_lsu_fp_stdata_bits_uop_debug_tsrc(core_io_lsu_fp_stdata_bits_uop_debug_tsrc),
    .io_lsu_fp_stdata_bits_data(core_io_lsu_fp_stdata_bits_data),
    .io_lsu_fp_stdata_bits_predicated(core_io_lsu_fp_stdata_bits_predicated),
    .io_lsu_fp_stdata_bits_fflags_valid(core_io_lsu_fp_stdata_bits_fflags_valid),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_switch(core_io_lsu_fp_stdata_bits_fflags_bits_uop_switch),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_switch_off(core_io_lsu_fp_stdata_bits_fflags_bits_uop_switch_off),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_is_unicore(core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_unicore),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_shift(core_io_lsu_fp_stdata_bits_fflags_bits_uop_shift),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_lrs3_rtype(core_io_lsu_fp_stdata_bits_fflags_bits_uop_lrs3_rtype),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_rflag(core_io_lsu_fp_stdata_bits_fflags_bits_uop_rflag),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_wflag(core_io_lsu_fp_stdata_bits_fflags_bits_uop_wflag),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_prflag(core_io_lsu_fp_stdata_bits_fflags_bits_uop_prflag),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_pwflag(core_io_lsu_fp_stdata_bits_fflags_bits_uop_pwflag),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_pflag_busy(core_io_lsu_fp_stdata_bits_fflags_bits_uop_pflag_busy),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_stale_pflag(core_io_lsu_fp_stdata_bits_fflags_bits_uop_stale_pflag),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_op1_sel(core_io_lsu_fp_stdata_bits_fflags_bits_uop_op1_sel),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_op2_sel(core_io_lsu_fp_stdata_bits_fflags_bits_uop_op2_sel),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_split_num(core_io_lsu_fp_stdata_bits_fflags_bits_uop_split_num),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_self_index(core_io_lsu_fp_stdata_bits_fflags_bits_uop_self_index),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_rob_inst_idx(core_io_lsu_fp_stdata_bits_fflags_bits_uop_rob_inst_idx),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_address_num(core_io_lsu_fp_stdata_bits_fflags_bits_uop_address_num),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_uopc(core_io_lsu_fp_stdata_bits_fflags_bits_uop_uopc),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_inst(core_io_lsu_fp_stdata_bits_fflags_bits_uop_inst),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_debug_inst(core_io_lsu_fp_stdata_bits_fflags_bits_uop_debug_inst),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_is_rvc(core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_rvc),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_debug_pc(core_io_lsu_fp_stdata_bits_fflags_bits_uop_debug_pc),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_iq_type(core_io_lsu_fp_stdata_bits_fflags_bits_uop_iq_type),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_fu_code(core_io_lsu_fp_stdata_bits_fflags_bits_uop_fu_code),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_br_type(core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_br_type),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_op1_sel(core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_op1_sel),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_op2_sel(core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_op2_sel),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_imm_sel(core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_imm_sel),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_op_fcn(core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_op_fcn),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_fcn_dw(core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_fcn_dw),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_csr_cmd(core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_csr_cmd),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_is_load(core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_is_load),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_is_sta(core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_is_sta),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_is_std(core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_is_std),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_op3_sel(core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_op3_sel),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_iw_state(core_io_lsu_fp_stdata_bits_fflags_bits_uop_iw_state),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_iw_p1_poisoned(core_io_lsu_fp_stdata_bits_fflags_bits_uop_iw_p1_poisoned),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_iw_p2_poisoned(core_io_lsu_fp_stdata_bits_fflags_bits_uop_iw_p2_poisoned),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_is_br(core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_br),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_is_jalr(core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_jalr),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_is_jal(core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_jal),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_is_sfb(core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_sfb),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_br_mask(core_io_lsu_fp_stdata_bits_fflags_bits_uop_br_mask),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_br_tag(core_io_lsu_fp_stdata_bits_fflags_bits_uop_br_tag),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_ftq_idx(core_io_lsu_fp_stdata_bits_fflags_bits_uop_ftq_idx),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_edge_inst(core_io_lsu_fp_stdata_bits_fflags_bits_uop_edge_inst),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_pc_lob(core_io_lsu_fp_stdata_bits_fflags_bits_uop_pc_lob),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_taken(core_io_lsu_fp_stdata_bits_fflags_bits_uop_taken),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_imm_packed(core_io_lsu_fp_stdata_bits_fflags_bits_uop_imm_packed),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_csr_addr(core_io_lsu_fp_stdata_bits_fflags_bits_uop_csr_addr),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_rob_idx(core_io_lsu_fp_stdata_bits_fflags_bits_uop_rob_idx),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_ldq_idx(core_io_lsu_fp_stdata_bits_fflags_bits_uop_ldq_idx),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_stq_idx(core_io_lsu_fp_stdata_bits_fflags_bits_uop_stq_idx),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_rxq_idx(core_io_lsu_fp_stdata_bits_fflags_bits_uop_rxq_idx),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_pdst(core_io_lsu_fp_stdata_bits_fflags_bits_uop_pdst),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_prs1(core_io_lsu_fp_stdata_bits_fflags_bits_uop_prs1),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_prs2(core_io_lsu_fp_stdata_bits_fflags_bits_uop_prs2),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_prs3(core_io_lsu_fp_stdata_bits_fflags_bits_uop_prs3),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_ppred(core_io_lsu_fp_stdata_bits_fflags_bits_uop_ppred),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_prs1_busy(core_io_lsu_fp_stdata_bits_fflags_bits_uop_prs1_busy),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_prs2_busy(core_io_lsu_fp_stdata_bits_fflags_bits_uop_prs2_busy),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_prs3_busy(core_io_lsu_fp_stdata_bits_fflags_bits_uop_prs3_busy),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_ppred_busy(core_io_lsu_fp_stdata_bits_fflags_bits_uop_ppred_busy),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_stale_pdst(core_io_lsu_fp_stdata_bits_fflags_bits_uop_stale_pdst),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_exception(core_io_lsu_fp_stdata_bits_fflags_bits_uop_exception),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_exc_cause(core_io_lsu_fp_stdata_bits_fflags_bits_uop_exc_cause),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_bypassable(core_io_lsu_fp_stdata_bits_fflags_bits_uop_bypassable),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_mem_cmd(core_io_lsu_fp_stdata_bits_fflags_bits_uop_mem_cmd),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_mem_size(core_io_lsu_fp_stdata_bits_fflags_bits_uop_mem_size),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_mem_signed(core_io_lsu_fp_stdata_bits_fflags_bits_uop_mem_signed),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_is_fence(core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_fence),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_is_fencei(core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_fencei),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_is_amo(core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_amo),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_uses_ldq(core_io_lsu_fp_stdata_bits_fflags_bits_uop_uses_ldq),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_uses_stq(core_io_lsu_fp_stdata_bits_fflags_bits_uop_uses_stq),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_is_sys_pc2epc(core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_sys_pc2epc),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_is_unique(core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_unique),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_flush_on_commit(core_io_lsu_fp_stdata_bits_fflags_bits_uop_flush_on_commit),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_ldst_is_rs1(core_io_lsu_fp_stdata_bits_fflags_bits_uop_ldst_is_rs1),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_ldst(core_io_lsu_fp_stdata_bits_fflags_bits_uop_ldst),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_lrs1(core_io_lsu_fp_stdata_bits_fflags_bits_uop_lrs1),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_lrs2(core_io_lsu_fp_stdata_bits_fflags_bits_uop_lrs2),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_lrs3(core_io_lsu_fp_stdata_bits_fflags_bits_uop_lrs3),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_ldst_val(core_io_lsu_fp_stdata_bits_fflags_bits_uop_ldst_val),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_dst_rtype(core_io_lsu_fp_stdata_bits_fflags_bits_uop_dst_rtype),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_lrs1_rtype(core_io_lsu_fp_stdata_bits_fflags_bits_uop_lrs1_rtype),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_lrs2_rtype(core_io_lsu_fp_stdata_bits_fflags_bits_uop_lrs2_rtype),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_frs3_en(core_io_lsu_fp_stdata_bits_fflags_bits_uop_frs3_en),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_fp_val(core_io_lsu_fp_stdata_bits_fflags_bits_uop_fp_val),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_fp_single(core_io_lsu_fp_stdata_bits_fflags_bits_uop_fp_single),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_xcpt_pf_if(core_io_lsu_fp_stdata_bits_fflags_bits_uop_xcpt_pf_if),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_xcpt_ae_if(core_io_lsu_fp_stdata_bits_fflags_bits_uop_xcpt_ae_if),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_xcpt_ma_if(core_io_lsu_fp_stdata_bits_fflags_bits_uop_xcpt_ma_if),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_bp_debug_if(core_io_lsu_fp_stdata_bits_fflags_bits_uop_bp_debug_if),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_bp_xcpt_if(core_io_lsu_fp_stdata_bits_fflags_bits_uop_bp_xcpt_if),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_debug_fsrc(core_io_lsu_fp_stdata_bits_fflags_bits_uop_debug_fsrc),
    .io_lsu_fp_stdata_bits_fflags_bits_uop_debug_tsrc(core_io_lsu_fp_stdata_bits_fflags_bits_uop_debug_tsrc),
    .io_lsu_fp_stdata_bits_fflags_bits_flags(core_io_lsu_fp_stdata_bits_fflags_bits_flags),
    .io_lsu_fp_stdata_bits_flagdata(core_io_lsu_fp_stdata_bits_flagdata),
    .io_lsu_fp_stdata_bits_fflagdata_valid(core_io_lsu_fp_stdata_bits_fflagdata_valid),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_switch(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_switch),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_switch_off(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_switch_off),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_unicore(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_unicore),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_shift(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_shift),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs3_rtype(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs3_rtype),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_rflag(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_rflag),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_wflag(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_wflag),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_prflag(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_prflag),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_pwflag(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_pwflag),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_pflag_busy(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_pflag_busy),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_stale_pflag(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_stale_pflag),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_op1_sel(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_op1_sel),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_op2_sel(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_op2_sel),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_split_num(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_split_num),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_self_index(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_self_index),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_rob_inst_idx(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_rob_inst_idx),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_address_num(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_address_num),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_uopc(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_uopc),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_inst(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_inst),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_debug_inst(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_debug_inst),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_rvc(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_rvc),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_debug_pc(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_debug_pc),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_iq_type(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_iq_type),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_fu_code(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_fu_code),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_br_type(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_br_type),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_op1_sel(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_op1_sel),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_op2_sel(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_op2_sel),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_imm_sel(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_imm_sel),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_op_fcn(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_op_fcn),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_fcn_dw(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_fcn_dw),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_csr_cmd(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_csr_cmd),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_load(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_load),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_sta(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_sta),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_std(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_std),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_op3_sel(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_op3_sel),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_iw_state(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_iw_state),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_iw_p1_poisoned(
      core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_iw_p1_poisoned),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_iw_p2_poisoned(
      core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_iw_p2_poisoned),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_br(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_br),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_jalr(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_jalr),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_jal(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_jal),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_sfb(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_sfb),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_br_mask(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_br_mask),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_br_tag(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_br_tag),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_ftq_idx(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ftq_idx),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_edge_inst(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_edge_inst),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_pc_lob(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_pc_lob),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_taken(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_taken),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_imm_packed(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_imm_packed),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_csr_addr(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_csr_addr),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_rob_idx(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_rob_idx),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_ldq_idx(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ldq_idx),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_stq_idx(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_stq_idx),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_rxq_idx(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_rxq_idx),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_pdst(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_pdst),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs1(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs1),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs2(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs2),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs3(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs3),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_ppred(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ppred),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs1_busy(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs1_busy),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs2_busy(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs2_busy),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs3_busy(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs3_busy),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_ppred_busy(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ppred_busy),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_stale_pdst(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_stale_pdst),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_exception(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_exception),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_exc_cause(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_exc_cause),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_bypassable(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_bypassable),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_mem_cmd(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_mem_cmd),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_mem_size(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_mem_size),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_mem_signed(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_mem_signed),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_fence(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_fence),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_fencei(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_fencei),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_amo(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_amo),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_uses_ldq(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_uses_ldq),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_uses_stq(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_uses_stq),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_sys_pc2epc(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_sys_pc2epc)
      ,
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_unique(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_unique),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_flush_on_commit(
      core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_flush_on_commit),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_ldst_is_rs1(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ldst_is_rs1),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_ldst(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ldst),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs1(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs1),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs2(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs2),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs3(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs3),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_ldst_val(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ldst_val),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_dst_rtype(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_dst_rtype),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs1_rtype(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs1_rtype),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs2_rtype(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs2_rtype),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_frs3_en(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_frs3_en),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_fp_val(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_fp_val),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_fp_single(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_fp_single),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_xcpt_pf_if(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_xcpt_pf_if),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_xcpt_ae_if(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_xcpt_ae_if),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_xcpt_ma_if(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_xcpt_ma_if),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_bp_debug_if(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_bp_debug_if),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_bp_xcpt_if(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_bp_xcpt_if),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_debug_fsrc(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_debug_fsrc),
    .io_lsu_fp_stdata_bits_fflagdata_bits_uop_debug_tsrc(core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_debug_tsrc),
    .io_lsu_fp_stdata_bits_fflagdata_bits_fflag(core_io_lsu_fp_stdata_bits_fflagdata_bits_fflag),
    .io_lsu_commit_valids_0(core_io_lsu_commit_valids_0),
    .io_lsu_commit_valids_1(core_io_lsu_commit_valids_1),
    .io_lsu_commit_arch_valids_0(core_io_lsu_commit_arch_valids_0),
    .io_lsu_commit_arch_valids_1(core_io_lsu_commit_arch_valids_1),
    .io_lsu_commit_uops_0_switch(core_io_lsu_commit_uops_0_switch),
    .io_lsu_commit_uops_0_switch_off(core_io_lsu_commit_uops_0_switch_off),
    .io_lsu_commit_uops_0_is_unicore(core_io_lsu_commit_uops_0_is_unicore),
    .io_lsu_commit_uops_0_shift(core_io_lsu_commit_uops_0_shift),
    .io_lsu_commit_uops_0_lrs3_rtype(core_io_lsu_commit_uops_0_lrs3_rtype),
    .io_lsu_commit_uops_0_rflag(core_io_lsu_commit_uops_0_rflag),
    .io_lsu_commit_uops_0_wflag(core_io_lsu_commit_uops_0_wflag),
    .io_lsu_commit_uops_0_prflag(core_io_lsu_commit_uops_0_prflag),
    .io_lsu_commit_uops_0_pwflag(core_io_lsu_commit_uops_0_pwflag),
    .io_lsu_commit_uops_0_pflag_busy(core_io_lsu_commit_uops_0_pflag_busy),
    .io_lsu_commit_uops_0_stale_pflag(core_io_lsu_commit_uops_0_stale_pflag),
    .io_lsu_commit_uops_0_op1_sel(core_io_lsu_commit_uops_0_op1_sel),
    .io_lsu_commit_uops_0_op2_sel(core_io_lsu_commit_uops_0_op2_sel),
    .io_lsu_commit_uops_0_split_num(core_io_lsu_commit_uops_0_split_num),
    .io_lsu_commit_uops_0_self_index(core_io_lsu_commit_uops_0_self_index),
    .io_lsu_commit_uops_0_rob_inst_idx(core_io_lsu_commit_uops_0_rob_inst_idx),
    .io_lsu_commit_uops_0_address_num(core_io_lsu_commit_uops_0_address_num),
    .io_lsu_commit_uops_0_uopc(core_io_lsu_commit_uops_0_uopc),
    .io_lsu_commit_uops_0_inst(core_io_lsu_commit_uops_0_inst),
    .io_lsu_commit_uops_0_debug_inst(core_io_lsu_commit_uops_0_debug_inst),
    .io_lsu_commit_uops_0_is_rvc(core_io_lsu_commit_uops_0_is_rvc),
    .io_lsu_commit_uops_0_debug_pc(core_io_lsu_commit_uops_0_debug_pc),
    .io_lsu_commit_uops_0_iq_type(core_io_lsu_commit_uops_0_iq_type),
    .io_lsu_commit_uops_0_fu_code(core_io_lsu_commit_uops_0_fu_code),
    .io_lsu_commit_uops_0_ctrl_br_type(core_io_lsu_commit_uops_0_ctrl_br_type),
    .io_lsu_commit_uops_0_ctrl_op1_sel(core_io_lsu_commit_uops_0_ctrl_op1_sel),
    .io_lsu_commit_uops_0_ctrl_op2_sel(core_io_lsu_commit_uops_0_ctrl_op2_sel),
    .io_lsu_commit_uops_0_ctrl_imm_sel(core_io_lsu_commit_uops_0_ctrl_imm_sel),
    .io_lsu_commit_uops_0_ctrl_op_fcn(core_io_lsu_commit_uops_0_ctrl_op_fcn),
    .io_lsu_commit_uops_0_ctrl_fcn_dw(core_io_lsu_commit_uops_0_ctrl_fcn_dw),
    .io_lsu_commit_uops_0_ctrl_csr_cmd(core_io_lsu_commit_uops_0_ctrl_csr_cmd),
    .io_lsu_commit_uops_0_ctrl_is_load(core_io_lsu_commit_uops_0_ctrl_is_load),
    .io_lsu_commit_uops_0_ctrl_is_sta(core_io_lsu_commit_uops_0_ctrl_is_sta),
    .io_lsu_commit_uops_0_ctrl_is_std(core_io_lsu_commit_uops_0_ctrl_is_std),
    .io_lsu_commit_uops_0_ctrl_op3_sel(core_io_lsu_commit_uops_0_ctrl_op3_sel),
    .io_lsu_commit_uops_0_iw_state(core_io_lsu_commit_uops_0_iw_state),
    .io_lsu_commit_uops_0_iw_p1_poisoned(core_io_lsu_commit_uops_0_iw_p1_poisoned),
    .io_lsu_commit_uops_0_iw_p2_poisoned(core_io_lsu_commit_uops_0_iw_p2_poisoned),
    .io_lsu_commit_uops_0_is_br(core_io_lsu_commit_uops_0_is_br),
    .io_lsu_commit_uops_0_is_jalr(core_io_lsu_commit_uops_0_is_jalr),
    .io_lsu_commit_uops_0_is_jal(core_io_lsu_commit_uops_0_is_jal),
    .io_lsu_commit_uops_0_is_sfb(core_io_lsu_commit_uops_0_is_sfb),
    .io_lsu_commit_uops_0_br_mask(core_io_lsu_commit_uops_0_br_mask),
    .io_lsu_commit_uops_0_br_tag(core_io_lsu_commit_uops_0_br_tag),
    .io_lsu_commit_uops_0_ftq_idx(core_io_lsu_commit_uops_0_ftq_idx),
    .io_lsu_commit_uops_0_edge_inst(core_io_lsu_commit_uops_0_edge_inst),
    .io_lsu_commit_uops_0_pc_lob(core_io_lsu_commit_uops_0_pc_lob),
    .io_lsu_commit_uops_0_taken(core_io_lsu_commit_uops_0_taken),
    .io_lsu_commit_uops_0_imm_packed(core_io_lsu_commit_uops_0_imm_packed),
    .io_lsu_commit_uops_0_csr_addr(core_io_lsu_commit_uops_0_csr_addr),
    .io_lsu_commit_uops_0_rob_idx(core_io_lsu_commit_uops_0_rob_idx),
    .io_lsu_commit_uops_0_ldq_idx(core_io_lsu_commit_uops_0_ldq_idx),
    .io_lsu_commit_uops_0_stq_idx(core_io_lsu_commit_uops_0_stq_idx),
    .io_lsu_commit_uops_0_rxq_idx(core_io_lsu_commit_uops_0_rxq_idx),
    .io_lsu_commit_uops_0_pdst(core_io_lsu_commit_uops_0_pdst),
    .io_lsu_commit_uops_0_prs1(core_io_lsu_commit_uops_0_prs1),
    .io_lsu_commit_uops_0_prs2(core_io_lsu_commit_uops_0_prs2),
    .io_lsu_commit_uops_0_prs3(core_io_lsu_commit_uops_0_prs3),
    .io_lsu_commit_uops_0_ppred(core_io_lsu_commit_uops_0_ppred),
    .io_lsu_commit_uops_0_prs1_busy(core_io_lsu_commit_uops_0_prs1_busy),
    .io_lsu_commit_uops_0_prs2_busy(core_io_lsu_commit_uops_0_prs2_busy),
    .io_lsu_commit_uops_0_prs3_busy(core_io_lsu_commit_uops_0_prs3_busy),
    .io_lsu_commit_uops_0_ppred_busy(core_io_lsu_commit_uops_0_ppred_busy),
    .io_lsu_commit_uops_0_stale_pdst(core_io_lsu_commit_uops_0_stale_pdst),
    .io_lsu_commit_uops_0_exception(core_io_lsu_commit_uops_0_exception),
    .io_lsu_commit_uops_0_exc_cause(core_io_lsu_commit_uops_0_exc_cause),
    .io_lsu_commit_uops_0_bypassable(core_io_lsu_commit_uops_0_bypassable),
    .io_lsu_commit_uops_0_mem_cmd(core_io_lsu_commit_uops_0_mem_cmd),
    .io_lsu_commit_uops_0_mem_size(core_io_lsu_commit_uops_0_mem_size),
    .io_lsu_commit_uops_0_mem_signed(core_io_lsu_commit_uops_0_mem_signed),
    .io_lsu_commit_uops_0_is_fence(core_io_lsu_commit_uops_0_is_fence),
    .io_lsu_commit_uops_0_is_fencei(core_io_lsu_commit_uops_0_is_fencei),
    .io_lsu_commit_uops_0_is_amo(core_io_lsu_commit_uops_0_is_amo),
    .io_lsu_commit_uops_0_uses_ldq(core_io_lsu_commit_uops_0_uses_ldq),
    .io_lsu_commit_uops_0_uses_stq(core_io_lsu_commit_uops_0_uses_stq),
    .io_lsu_commit_uops_0_is_sys_pc2epc(core_io_lsu_commit_uops_0_is_sys_pc2epc),
    .io_lsu_commit_uops_0_is_unique(core_io_lsu_commit_uops_0_is_unique),
    .io_lsu_commit_uops_0_flush_on_commit(core_io_lsu_commit_uops_0_flush_on_commit),
    .io_lsu_commit_uops_0_ldst_is_rs1(core_io_lsu_commit_uops_0_ldst_is_rs1),
    .io_lsu_commit_uops_0_ldst(core_io_lsu_commit_uops_0_ldst),
    .io_lsu_commit_uops_0_lrs1(core_io_lsu_commit_uops_0_lrs1),
    .io_lsu_commit_uops_0_lrs2(core_io_lsu_commit_uops_0_lrs2),
    .io_lsu_commit_uops_0_lrs3(core_io_lsu_commit_uops_0_lrs3),
    .io_lsu_commit_uops_0_ldst_val(core_io_lsu_commit_uops_0_ldst_val),
    .io_lsu_commit_uops_0_dst_rtype(core_io_lsu_commit_uops_0_dst_rtype),
    .io_lsu_commit_uops_0_lrs1_rtype(core_io_lsu_commit_uops_0_lrs1_rtype),
    .io_lsu_commit_uops_0_lrs2_rtype(core_io_lsu_commit_uops_0_lrs2_rtype),
    .io_lsu_commit_uops_0_frs3_en(core_io_lsu_commit_uops_0_frs3_en),
    .io_lsu_commit_uops_0_fp_val(core_io_lsu_commit_uops_0_fp_val),
    .io_lsu_commit_uops_0_fp_single(core_io_lsu_commit_uops_0_fp_single),
    .io_lsu_commit_uops_0_xcpt_pf_if(core_io_lsu_commit_uops_0_xcpt_pf_if),
    .io_lsu_commit_uops_0_xcpt_ae_if(core_io_lsu_commit_uops_0_xcpt_ae_if),
    .io_lsu_commit_uops_0_xcpt_ma_if(core_io_lsu_commit_uops_0_xcpt_ma_if),
    .io_lsu_commit_uops_0_bp_debug_if(core_io_lsu_commit_uops_0_bp_debug_if),
    .io_lsu_commit_uops_0_bp_xcpt_if(core_io_lsu_commit_uops_0_bp_xcpt_if),
    .io_lsu_commit_uops_0_debug_fsrc(core_io_lsu_commit_uops_0_debug_fsrc),
    .io_lsu_commit_uops_0_debug_tsrc(core_io_lsu_commit_uops_0_debug_tsrc),
    .io_lsu_commit_uops_1_switch(core_io_lsu_commit_uops_1_switch),
    .io_lsu_commit_uops_1_switch_off(core_io_lsu_commit_uops_1_switch_off),
    .io_lsu_commit_uops_1_is_unicore(core_io_lsu_commit_uops_1_is_unicore),
    .io_lsu_commit_uops_1_shift(core_io_lsu_commit_uops_1_shift),
    .io_lsu_commit_uops_1_lrs3_rtype(core_io_lsu_commit_uops_1_lrs3_rtype),
    .io_lsu_commit_uops_1_rflag(core_io_lsu_commit_uops_1_rflag),
    .io_lsu_commit_uops_1_wflag(core_io_lsu_commit_uops_1_wflag),
    .io_lsu_commit_uops_1_prflag(core_io_lsu_commit_uops_1_prflag),
    .io_lsu_commit_uops_1_pwflag(core_io_lsu_commit_uops_1_pwflag),
    .io_lsu_commit_uops_1_pflag_busy(core_io_lsu_commit_uops_1_pflag_busy),
    .io_lsu_commit_uops_1_stale_pflag(core_io_lsu_commit_uops_1_stale_pflag),
    .io_lsu_commit_uops_1_op1_sel(core_io_lsu_commit_uops_1_op1_sel),
    .io_lsu_commit_uops_1_op2_sel(core_io_lsu_commit_uops_1_op2_sel),
    .io_lsu_commit_uops_1_split_num(core_io_lsu_commit_uops_1_split_num),
    .io_lsu_commit_uops_1_self_index(core_io_lsu_commit_uops_1_self_index),
    .io_lsu_commit_uops_1_rob_inst_idx(core_io_lsu_commit_uops_1_rob_inst_idx),
    .io_lsu_commit_uops_1_address_num(core_io_lsu_commit_uops_1_address_num),
    .io_lsu_commit_uops_1_uopc(core_io_lsu_commit_uops_1_uopc),
    .io_lsu_commit_uops_1_inst(core_io_lsu_commit_uops_1_inst),
    .io_lsu_commit_uops_1_debug_inst(core_io_lsu_commit_uops_1_debug_inst),
    .io_lsu_commit_uops_1_is_rvc(core_io_lsu_commit_uops_1_is_rvc),
    .io_lsu_commit_uops_1_debug_pc(core_io_lsu_commit_uops_1_debug_pc),
    .io_lsu_commit_uops_1_iq_type(core_io_lsu_commit_uops_1_iq_type),
    .io_lsu_commit_uops_1_fu_code(core_io_lsu_commit_uops_1_fu_code),
    .io_lsu_commit_uops_1_ctrl_br_type(core_io_lsu_commit_uops_1_ctrl_br_type),
    .io_lsu_commit_uops_1_ctrl_op1_sel(core_io_lsu_commit_uops_1_ctrl_op1_sel),
    .io_lsu_commit_uops_1_ctrl_op2_sel(core_io_lsu_commit_uops_1_ctrl_op2_sel),
    .io_lsu_commit_uops_1_ctrl_imm_sel(core_io_lsu_commit_uops_1_ctrl_imm_sel),
    .io_lsu_commit_uops_1_ctrl_op_fcn(core_io_lsu_commit_uops_1_ctrl_op_fcn),
    .io_lsu_commit_uops_1_ctrl_fcn_dw(core_io_lsu_commit_uops_1_ctrl_fcn_dw),
    .io_lsu_commit_uops_1_ctrl_csr_cmd(core_io_lsu_commit_uops_1_ctrl_csr_cmd),
    .io_lsu_commit_uops_1_ctrl_is_load(core_io_lsu_commit_uops_1_ctrl_is_load),
    .io_lsu_commit_uops_1_ctrl_is_sta(core_io_lsu_commit_uops_1_ctrl_is_sta),
    .io_lsu_commit_uops_1_ctrl_is_std(core_io_lsu_commit_uops_1_ctrl_is_std),
    .io_lsu_commit_uops_1_ctrl_op3_sel(core_io_lsu_commit_uops_1_ctrl_op3_sel),
    .io_lsu_commit_uops_1_iw_state(core_io_lsu_commit_uops_1_iw_state),
    .io_lsu_commit_uops_1_iw_p1_poisoned(core_io_lsu_commit_uops_1_iw_p1_poisoned),
    .io_lsu_commit_uops_1_iw_p2_poisoned(core_io_lsu_commit_uops_1_iw_p2_poisoned),
    .io_lsu_commit_uops_1_is_br(core_io_lsu_commit_uops_1_is_br),
    .io_lsu_commit_uops_1_is_jalr(core_io_lsu_commit_uops_1_is_jalr),
    .io_lsu_commit_uops_1_is_jal(core_io_lsu_commit_uops_1_is_jal),
    .io_lsu_commit_uops_1_is_sfb(core_io_lsu_commit_uops_1_is_sfb),
    .io_lsu_commit_uops_1_br_mask(core_io_lsu_commit_uops_1_br_mask),
    .io_lsu_commit_uops_1_br_tag(core_io_lsu_commit_uops_1_br_tag),
    .io_lsu_commit_uops_1_ftq_idx(core_io_lsu_commit_uops_1_ftq_idx),
    .io_lsu_commit_uops_1_edge_inst(core_io_lsu_commit_uops_1_edge_inst),
    .io_lsu_commit_uops_1_pc_lob(core_io_lsu_commit_uops_1_pc_lob),
    .io_lsu_commit_uops_1_taken(core_io_lsu_commit_uops_1_taken),
    .io_lsu_commit_uops_1_imm_packed(core_io_lsu_commit_uops_1_imm_packed),
    .io_lsu_commit_uops_1_csr_addr(core_io_lsu_commit_uops_1_csr_addr),
    .io_lsu_commit_uops_1_rob_idx(core_io_lsu_commit_uops_1_rob_idx),
    .io_lsu_commit_uops_1_ldq_idx(core_io_lsu_commit_uops_1_ldq_idx),
    .io_lsu_commit_uops_1_stq_idx(core_io_lsu_commit_uops_1_stq_idx),
    .io_lsu_commit_uops_1_rxq_idx(core_io_lsu_commit_uops_1_rxq_idx),
    .io_lsu_commit_uops_1_pdst(core_io_lsu_commit_uops_1_pdst),
    .io_lsu_commit_uops_1_prs1(core_io_lsu_commit_uops_1_prs1),
    .io_lsu_commit_uops_1_prs2(core_io_lsu_commit_uops_1_prs2),
    .io_lsu_commit_uops_1_prs3(core_io_lsu_commit_uops_1_prs3),
    .io_lsu_commit_uops_1_ppred(core_io_lsu_commit_uops_1_ppred),
    .io_lsu_commit_uops_1_prs1_busy(core_io_lsu_commit_uops_1_prs1_busy),
    .io_lsu_commit_uops_1_prs2_busy(core_io_lsu_commit_uops_1_prs2_busy),
    .io_lsu_commit_uops_1_prs3_busy(core_io_lsu_commit_uops_1_prs3_busy),
    .io_lsu_commit_uops_1_ppred_busy(core_io_lsu_commit_uops_1_ppred_busy),
    .io_lsu_commit_uops_1_stale_pdst(core_io_lsu_commit_uops_1_stale_pdst),
    .io_lsu_commit_uops_1_exception(core_io_lsu_commit_uops_1_exception),
    .io_lsu_commit_uops_1_exc_cause(core_io_lsu_commit_uops_1_exc_cause),
    .io_lsu_commit_uops_1_bypassable(core_io_lsu_commit_uops_1_bypassable),
    .io_lsu_commit_uops_1_mem_cmd(core_io_lsu_commit_uops_1_mem_cmd),
    .io_lsu_commit_uops_1_mem_size(core_io_lsu_commit_uops_1_mem_size),
    .io_lsu_commit_uops_1_mem_signed(core_io_lsu_commit_uops_1_mem_signed),
    .io_lsu_commit_uops_1_is_fence(core_io_lsu_commit_uops_1_is_fence),
    .io_lsu_commit_uops_1_is_fencei(core_io_lsu_commit_uops_1_is_fencei),
    .io_lsu_commit_uops_1_is_amo(core_io_lsu_commit_uops_1_is_amo),
    .io_lsu_commit_uops_1_uses_ldq(core_io_lsu_commit_uops_1_uses_ldq),
    .io_lsu_commit_uops_1_uses_stq(core_io_lsu_commit_uops_1_uses_stq),
    .io_lsu_commit_uops_1_is_sys_pc2epc(core_io_lsu_commit_uops_1_is_sys_pc2epc),
    .io_lsu_commit_uops_1_is_unique(core_io_lsu_commit_uops_1_is_unique),
    .io_lsu_commit_uops_1_flush_on_commit(core_io_lsu_commit_uops_1_flush_on_commit),
    .io_lsu_commit_uops_1_ldst_is_rs1(core_io_lsu_commit_uops_1_ldst_is_rs1),
    .io_lsu_commit_uops_1_ldst(core_io_lsu_commit_uops_1_ldst),
    .io_lsu_commit_uops_1_lrs1(core_io_lsu_commit_uops_1_lrs1),
    .io_lsu_commit_uops_1_lrs2(core_io_lsu_commit_uops_1_lrs2),
    .io_lsu_commit_uops_1_lrs3(core_io_lsu_commit_uops_1_lrs3),
    .io_lsu_commit_uops_1_ldst_val(core_io_lsu_commit_uops_1_ldst_val),
    .io_lsu_commit_uops_1_dst_rtype(core_io_lsu_commit_uops_1_dst_rtype),
    .io_lsu_commit_uops_1_lrs1_rtype(core_io_lsu_commit_uops_1_lrs1_rtype),
    .io_lsu_commit_uops_1_lrs2_rtype(core_io_lsu_commit_uops_1_lrs2_rtype),
    .io_lsu_commit_uops_1_frs3_en(core_io_lsu_commit_uops_1_frs3_en),
    .io_lsu_commit_uops_1_fp_val(core_io_lsu_commit_uops_1_fp_val),
    .io_lsu_commit_uops_1_fp_single(core_io_lsu_commit_uops_1_fp_single),
    .io_lsu_commit_uops_1_xcpt_pf_if(core_io_lsu_commit_uops_1_xcpt_pf_if),
    .io_lsu_commit_uops_1_xcpt_ae_if(core_io_lsu_commit_uops_1_xcpt_ae_if),
    .io_lsu_commit_uops_1_xcpt_ma_if(core_io_lsu_commit_uops_1_xcpt_ma_if),
    .io_lsu_commit_uops_1_bp_debug_if(core_io_lsu_commit_uops_1_bp_debug_if),
    .io_lsu_commit_uops_1_bp_xcpt_if(core_io_lsu_commit_uops_1_bp_xcpt_if),
    .io_lsu_commit_uops_1_debug_fsrc(core_io_lsu_commit_uops_1_debug_fsrc),
    .io_lsu_commit_uops_1_debug_tsrc(core_io_lsu_commit_uops_1_debug_tsrc),
    .io_lsu_commit_fflags_valid(core_io_lsu_commit_fflags_valid),
    .io_lsu_commit_fflags_bits(core_io_lsu_commit_fflags_bits),
    .io_lsu_commit_fflag_exception_valid(core_io_lsu_commit_fflag_exception_valid),
    .io_lsu_commit_fflag_exception_bits(core_io_lsu_commit_fflag_exception_bits),
    .io_lsu_commit_debug_insts_0(core_io_lsu_commit_debug_insts_0),
    .io_lsu_commit_debug_insts_1(core_io_lsu_commit_debug_insts_1),
    .io_lsu_commit_rbk_valids_0(core_io_lsu_commit_rbk_valids_0),
    .io_lsu_commit_rbk_valids_1(core_io_lsu_commit_rbk_valids_1),
    .io_lsu_commit_rollback(core_io_lsu_commit_rollback),
    .io_lsu_commit_debug_wdata_0(core_io_lsu_commit_debug_wdata_0),
    .io_lsu_commit_debug_wdata_1(core_io_lsu_commit_debug_wdata_1),
    .io_lsu_commit_debug_wflagdata_0(core_io_lsu_commit_debug_wflagdata_0),
    .io_lsu_commit_debug_wflagdata_1(core_io_lsu_commit_debug_wflagdata_1),
    .io_lsu_commit_load_at_rob_head(core_io_lsu_commit_load_at_rob_head),
    .io_lsu_clr_bsy_0_valid(core_io_lsu_clr_bsy_0_valid),
    .io_lsu_clr_bsy_0_bits(core_io_lsu_clr_bsy_0_bits),
    .io_lsu_clr_bsy_1_valid(core_io_lsu_clr_bsy_1_valid),
    .io_lsu_clr_bsy_1_bits(core_io_lsu_clr_bsy_1_bits),
    .io_lsu_clr_unsafe_0_valid(core_io_lsu_clr_unsafe_0_valid),
    .io_lsu_clr_unsafe_0_bits(core_io_lsu_clr_unsafe_0_bits),
    .io_lsu_clr_bsy_first_idx_0(core_io_lsu_clr_bsy_first_idx_0),
    .io_lsu_clr_bsy_first_idx_1(core_io_lsu_clr_bsy_first_idx_1),
    .io_lsu_clr_bsy_self_idx_0(core_io_lsu_clr_bsy_self_idx_0),
    .io_lsu_clr_bsy_self_idx_1(core_io_lsu_clr_bsy_self_idx_1),
    .io_lsu_fence_dmem(core_io_lsu_fence_dmem),
    .io_lsu_spec_ld_wakeup_0_valid(core_io_lsu_spec_ld_wakeup_0_valid),
    .io_lsu_spec_ld_wakeup_0_bits(core_io_lsu_spec_ld_wakeup_0_bits),
    .io_lsu_ld_miss(core_io_lsu_ld_miss),
    .io_lsu_brupdate_b1_resolve_mask(core_io_lsu_brupdate_b1_resolve_mask),
    .io_lsu_brupdate_b1_mispredict_mask(core_io_lsu_brupdate_b1_mispredict_mask),
    .io_lsu_brupdate_b2_uop_switch(core_io_lsu_brupdate_b2_uop_switch),
    .io_lsu_brupdate_b2_uop_switch_off(core_io_lsu_brupdate_b2_uop_switch_off),
    .io_lsu_brupdate_b2_uop_is_unicore(core_io_lsu_brupdate_b2_uop_is_unicore),
    .io_lsu_brupdate_b2_uop_shift(core_io_lsu_brupdate_b2_uop_shift),
    .io_lsu_brupdate_b2_uop_lrs3_rtype(core_io_lsu_brupdate_b2_uop_lrs3_rtype),
    .io_lsu_brupdate_b2_uop_rflag(core_io_lsu_brupdate_b2_uop_rflag),
    .io_lsu_brupdate_b2_uop_wflag(core_io_lsu_brupdate_b2_uop_wflag),
    .io_lsu_brupdate_b2_uop_prflag(core_io_lsu_brupdate_b2_uop_prflag),
    .io_lsu_brupdate_b2_uop_pwflag(core_io_lsu_brupdate_b2_uop_pwflag),
    .io_lsu_brupdate_b2_uop_pflag_busy(core_io_lsu_brupdate_b2_uop_pflag_busy),
    .io_lsu_brupdate_b2_uop_stale_pflag(core_io_lsu_brupdate_b2_uop_stale_pflag),
    .io_lsu_brupdate_b2_uop_op1_sel(core_io_lsu_brupdate_b2_uop_op1_sel),
    .io_lsu_brupdate_b2_uop_op2_sel(core_io_lsu_brupdate_b2_uop_op2_sel),
    .io_lsu_brupdate_b2_uop_split_num(core_io_lsu_brupdate_b2_uop_split_num),
    .io_lsu_brupdate_b2_uop_self_index(core_io_lsu_brupdate_b2_uop_self_index),
    .io_lsu_brupdate_b2_uop_rob_inst_idx(core_io_lsu_brupdate_b2_uop_rob_inst_idx),
    .io_lsu_brupdate_b2_uop_address_num(core_io_lsu_brupdate_b2_uop_address_num),
    .io_lsu_brupdate_b2_uop_uopc(core_io_lsu_brupdate_b2_uop_uopc),
    .io_lsu_brupdate_b2_uop_inst(core_io_lsu_brupdate_b2_uop_inst),
    .io_lsu_brupdate_b2_uop_debug_inst(core_io_lsu_brupdate_b2_uop_debug_inst),
    .io_lsu_brupdate_b2_uop_is_rvc(core_io_lsu_brupdate_b2_uop_is_rvc),
    .io_lsu_brupdate_b2_uop_debug_pc(core_io_lsu_brupdate_b2_uop_debug_pc),
    .io_lsu_brupdate_b2_uop_iq_type(core_io_lsu_brupdate_b2_uop_iq_type),
    .io_lsu_brupdate_b2_uop_fu_code(core_io_lsu_brupdate_b2_uop_fu_code),
    .io_lsu_brupdate_b2_uop_ctrl_br_type(core_io_lsu_brupdate_b2_uop_ctrl_br_type),
    .io_lsu_brupdate_b2_uop_ctrl_op1_sel(core_io_lsu_brupdate_b2_uop_ctrl_op1_sel),
    .io_lsu_brupdate_b2_uop_ctrl_op2_sel(core_io_lsu_brupdate_b2_uop_ctrl_op2_sel),
    .io_lsu_brupdate_b2_uop_ctrl_imm_sel(core_io_lsu_brupdate_b2_uop_ctrl_imm_sel),
    .io_lsu_brupdate_b2_uop_ctrl_op_fcn(core_io_lsu_brupdate_b2_uop_ctrl_op_fcn),
    .io_lsu_brupdate_b2_uop_ctrl_fcn_dw(core_io_lsu_brupdate_b2_uop_ctrl_fcn_dw),
    .io_lsu_brupdate_b2_uop_ctrl_csr_cmd(core_io_lsu_brupdate_b2_uop_ctrl_csr_cmd),
    .io_lsu_brupdate_b2_uop_ctrl_is_load(core_io_lsu_brupdate_b2_uop_ctrl_is_load),
    .io_lsu_brupdate_b2_uop_ctrl_is_sta(core_io_lsu_brupdate_b2_uop_ctrl_is_sta),
    .io_lsu_brupdate_b2_uop_ctrl_is_std(core_io_lsu_brupdate_b2_uop_ctrl_is_std),
    .io_lsu_brupdate_b2_uop_ctrl_op3_sel(core_io_lsu_brupdate_b2_uop_ctrl_op3_sel),
    .io_lsu_brupdate_b2_uop_iw_state(core_io_lsu_brupdate_b2_uop_iw_state),
    .io_lsu_brupdate_b2_uop_iw_p1_poisoned(core_io_lsu_brupdate_b2_uop_iw_p1_poisoned),
    .io_lsu_brupdate_b2_uop_iw_p2_poisoned(core_io_lsu_brupdate_b2_uop_iw_p2_poisoned),
    .io_lsu_brupdate_b2_uop_is_br(core_io_lsu_brupdate_b2_uop_is_br),
    .io_lsu_brupdate_b2_uop_is_jalr(core_io_lsu_brupdate_b2_uop_is_jalr),
    .io_lsu_brupdate_b2_uop_is_jal(core_io_lsu_brupdate_b2_uop_is_jal),
    .io_lsu_brupdate_b2_uop_is_sfb(core_io_lsu_brupdate_b2_uop_is_sfb),
    .io_lsu_brupdate_b2_uop_br_mask(core_io_lsu_brupdate_b2_uop_br_mask),
    .io_lsu_brupdate_b2_uop_br_tag(core_io_lsu_brupdate_b2_uop_br_tag),
    .io_lsu_brupdate_b2_uop_ftq_idx(core_io_lsu_brupdate_b2_uop_ftq_idx),
    .io_lsu_brupdate_b2_uop_edge_inst(core_io_lsu_brupdate_b2_uop_edge_inst),
    .io_lsu_brupdate_b2_uop_pc_lob(core_io_lsu_brupdate_b2_uop_pc_lob),
    .io_lsu_brupdate_b2_uop_taken(core_io_lsu_brupdate_b2_uop_taken),
    .io_lsu_brupdate_b2_uop_imm_packed(core_io_lsu_brupdate_b2_uop_imm_packed),
    .io_lsu_brupdate_b2_uop_csr_addr(core_io_lsu_brupdate_b2_uop_csr_addr),
    .io_lsu_brupdate_b2_uop_rob_idx(core_io_lsu_brupdate_b2_uop_rob_idx),
    .io_lsu_brupdate_b2_uop_ldq_idx(core_io_lsu_brupdate_b2_uop_ldq_idx),
    .io_lsu_brupdate_b2_uop_stq_idx(core_io_lsu_brupdate_b2_uop_stq_idx),
    .io_lsu_brupdate_b2_uop_rxq_idx(core_io_lsu_brupdate_b2_uop_rxq_idx),
    .io_lsu_brupdate_b2_uop_pdst(core_io_lsu_brupdate_b2_uop_pdst),
    .io_lsu_brupdate_b2_uop_prs1(core_io_lsu_brupdate_b2_uop_prs1),
    .io_lsu_brupdate_b2_uop_prs2(core_io_lsu_brupdate_b2_uop_prs2),
    .io_lsu_brupdate_b2_uop_prs3(core_io_lsu_brupdate_b2_uop_prs3),
    .io_lsu_brupdate_b2_uop_ppred(core_io_lsu_brupdate_b2_uop_ppred),
    .io_lsu_brupdate_b2_uop_prs1_busy(core_io_lsu_brupdate_b2_uop_prs1_busy),
    .io_lsu_brupdate_b2_uop_prs2_busy(core_io_lsu_brupdate_b2_uop_prs2_busy),
    .io_lsu_brupdate_b2_uop_prs3_busy(core_io_lsu_brupdate_b2_uop_prs3_busy),
    .io_lsu_brupdate_b2_uop_ppred_busy(core_io_lsu_brupdate_b2_uop_ppred_busy),
    .io_lsu_brupdate_b2_uop_stale_pdst(core_io_lsu_brupdate_b2_uop_stale_pdst),
    .io_lsu_brupdate_b2_uop_exception(core_io_lsu_brupdate_b2_uop_exception),
    .io_lsu_brupdate_b2_uop_exc_cause(core_io_lsu_brupdate_b2_uop_exc_cause),
    .io_lsu_brupdate_b2_uop_bypassable(core_io_lsu_brupdate_b2_uop_bypassable),
    .io_lsu_brupdate_b2_uop_mem_cmd(core_io_lsu_brupdate_b2_uop_mem_cmd),
    .io_lsu_brupdate_b2_uop_mem_size(core_io_lsu_brupdate_b2_uop_mem_size),
    .io_lsu_brupdate_b2_uop_mem_signed(core_io_lsu_brupdate_b2_uop_mem_signed),
    .io_lsu_brupdate_b2_uop_is_fence(core_io_lsu_brupdate_b2_uop_is_fence),
    .io_lsu_brupdate_b2_uop_is_fencei(core_io_lsu_brupdate_b2_uop_is_fencei),
    .io_lsu_brupdate_b2_uop_is_amo(core_io_lsu_brupdate_b2_uop_is_amo),
    .io_lsu_brupdate_b2_uop_uses_ldq(core_io_lsu_brupdate_b2_uop_uses_ldq),
    .io_lsu_brupdate_b2_uop_uses_stq(core_io_lsu_brupdate_b2_uop_uses_stq),
    .io_lsu_brupdate_b2_uop_is_sys_pc2epc(core_io_lsu_brupdate_b2_uop_is_sys_pc2epc),
    .io_lsu_brupdate_b2_uop_is_unique(core_io_lsu_brupdate_b2_uop_is_unique),
    .io_lsu_brupdate_b2_uop_flush_on_commit(core_io_lsu_brupdate_b2_uop_flush_on_commit),
    .io_lsu_brupdate_b2_uop_ldst_is_rs1(core_io_lsu_brupdate_b2_uop_ldst_is_rs1),
    .io_lsu_brupdate_b2_uop_ldst(core_io_lsu_brupdate_b2_uop_ldst),
    .io_lsu_brupdate_b2_uop_lrs1(core_io_lsu_brupdate_b2_uop_lrs1),
    .io_lsu_brupdate_b2_uop_lrs2(core_io_lsu_brupdate_b2_uop_lrs2),
    .io_lsu_brupdate_b2_uop_lrs3(core_io_lsu_brupdate_b2_uop_lrs3),
    .io_lsu_brupdate_b2_uop_ldst_val(core_io_lsu_brupdate_b2_uop_ldst_val),
    .io_lsu_brupdate_b2_uop_dst_rtype(core_io_lsu_brupdate_b2_uop_dst_rtype),
    .io_lsu_brupdate_b2_uop_lrs1_rtype(core_io_lsu_brupdate_b2_uop_lrs1_rtype),
    .io_lsu_brupdate_b2_uop_lrs2_rtype(core_io_lsu_brupdate_b2_uop_lrs2_rtype),
    .io_lsu_brupdate_b2_uop_frs3_en(core_io_lsu_brupdate_b2_uop_frs3_en),
    .io_lsu_brupdate_b2_uop_fp_val(core_io_lsu_brupdate_b2_uop_fp_val),
    .io_lsu_brupdate_b2_uop_fp_single(core_io_lsu_brupdate_b2_uop_fp_single),
    .io_lsu_brupdate_b2_uop_xcpt_pf_if(core_io_lsu_brupdate_b2_uop_xcpt_pf_if),
    .io_lsu_brupdate_b2_uop_xcpt_ae_if(core_io_lsu_brupdate_b2_uop_xcpt_ae_if),
    .io_lsu_brupdate_b2_uop_xcpt_ma_if(core_io_lsu_brupdate_b2_uop_xcpt_ma_if),
    .io_lsu_brupdate_b2_uop_bp_debug_if(core_io_lsu_brupdate_b2_uop_bp_debug_if),
    .io_lsu_brupdate_b2_uop_bp_xcpt_if(core_io_lsu_brupdate_b2_uop_bp_xcpt_if),
    .io_lsu_brupdate_b2_uop_debug_fsrc(core_io_lsu_brupdate_b2_uop_debug_fsrc),
    .io_lsu_brupdate_b2_uop_debug_tsrc(core_io_lsu_brupdate_b2_uop_debug_tsrc),
    .io_lsu_brupdate_b2_valid(core_io_lsu_brupdate_b2_valid),
    .io_lsu_brupdate_b2_mispredict(core_io_lsu_brupdate_b2_mispredict),
    .io_lsu_brupdate_b2_taken(core_io_lsu_brupdate_b2_taken),
    .io_lsu_brupdate_b2_cfi_type(core_io_lsu_brupdate_b2_cfi_type),
    .io_lsu_brupdate_b2_pc_sel(core_io_lsu_brupdate_b2_pc_sel),
    .io_lsu_brupdate_b2_jalr_target(core_io_lsu_brupdate_b2_jalr_target),
    .io_lsu_brupdate_b2_target_offset(core_io_lsu_brupdate_b2_target_offset),
    .io_lsu_rob_pnr_idx(core_io_lsu_rob_pnr_idx),
    .io_lsu_rob_head_idx(core_io_lsu_rob_head_idx),
    .io_lsu_exception(core_io_lsu_exception),
    .io_lsu_fencei_rdy(core_io_lsu_fencei_rdy),
    .io_lsu_lxcpt_valid(core_io_lsu_lxcpt_valid),
    .io_lsu_lxcpt_bits_uop_switch(core_io_lsu_lxcpt_bits_uop_switch),
    .io_lsu_lxcpt_bits_uop_switch_off(core_io_lsu_lxcpt_bits_uop_switch_off),
    .io_lsu_lxcpt_bits_uop_is_unicore(core_io_lsu_lxcpt_bits_uop_is_unicore),
    .io_lsu_lxcpt_bits_uop_shift(core_io_lsu_lxcpt_bits_uop_shift),
    .io_lsu_lxcpt_bits_uop_lrs3_rtype(core_io_lsu_lxcpt_bits_uop_lrs3_rtype),
    .io_lsu_lxcpt_bits_uop_rflag(core_io_lsu_lxcpt_bits_uop_rflag),
    .io_lsu_lxcpt_bits_uop_wflag(core_io_lsu_lxcpt_bits_uop_wflag),
    .io_lsu_lxcpt_bits_uop_prflag(core_io_lsu_lxcpt_bits_uop_prflag),
    .io_lsu_lxcpt_bits_uop_pwflag(core_io_lsu_lxcpt_bits_uop_pwflag),
    .io_lsu_lxcpt_bits_uop_pflag_busy(core_io_lsu_lxcpt_bits_uop_pflag_busy),
    .io_lsu_lxcpt_bits_uop_stale_pflag(core_io_lsu_lxcpt_bits_uop_stale_pflag),
    .io_lsu_lxcpt_bits_uop_op1_sel(core_io_lsu_lxcpt_bits_uop_op1_sel),
    .io_lsu_lxcpt_bits_uop_op2_sel(core_io_lsu_lxcpt_bits_uop_op2_sel),
    .io_lsu_lxcpt_bits_uop_split_num(core_io_lsu_lxcpt_bits_uop_split_num),
    .io_lsu_lxcpt_bits_uop_self_index(core_io_lsu_lxcpt_bits_uop_self_index),
    .io_lsu_lxcpt_bits_uop_rob_inst_idx(core_io_lsu_lxcpt_bits_uop_rob_inst_idx),
    .io_lsu_lxcpt_bits_uop_address_num(core_io_lsu_lxcpt_bits_uop_address_num),
    .io_lsu_lxcpt_bits_uop_uopc(core_io_lsu_lxcpt_bits_uop_uopc),
    .io_lsu_lxcpt_bits_uop_inst(core_io_lsu_lxcpt_bits_uop_inst),
    .io_lsu_lxcpt_bits_uop_debug_inst(core_io_lsu_lxcpt_bits_uop_debug_inst),
    .io_lsu_lxcpt_bits_uop_is_rvc(core_io_lsu_lxcpt_bits_uop_is_rvc),
    .io_lsu_lxcpt_bits_uop_debug_pc(core_io_lsu_lxcpt_bits_uop_debug_pc),
    .io_lsu_lxcpt_bits_uop_iq_type(core_io_lsu_lxcpt_bits_uop_iq_type),
    .io_lsu_lxcpt_bits_uop_fu_code(core_io_lsu_lxcpt_bits_uop_fu_code),
    .io_lsu_lxcpt_bits_uop_ctrl_br_type(core_io_lsu_lxcpt_bits_uop_ctrl_br_type),
    .io_lsu_lxcpt_bits_uop_ctrl_op1_sel(core_io_lsu_lxcpt_bits_uop_ctrl_op1_sel),
    .io_lsu_lxcpt_bits_uop_ctrl_op2_sel(core_io_lsu_lxcpt_bits_uop_ctrl_op2_sel),
    .io_lsu_lxcpt_bits_uop_ctrl_imm_sel(core_io_lsu_lxcpt_bits_uop_ctrl_imm_sel),
    .io_lsu_lxcpt_bits_uop_ctrl_op_fcn(core_io_lsu_lxcpt_bits_uop_ctrl_op_fcn),
    .io_lsu_lxcpt_bits_uop_ctrl_fcn_dw(core_io_lsu_lxcpt_bits_uop_ctrl_fcn_dw),
    .io_lsu_lxcpt_bits_uop_ctrl_csr_cmd(core_io_lsu_lxcpt_bits_uop_ctrl_csr_cmd),
    .io_lsu_lxcpt_bits_uop_ctrl_is_load(core_io_lsu_lxcpt_bits_uop_ctrl_is_load),
    .io_lsu_lxcpt_bits_uop_ctrl_is_sta(core_io_lsu_lxcpt_bits_uop_ctrl_is_sta),
    .io_lsu_lxcpt_bits_uop_ctrl_is_std(core_io_lsu_lxcpt_bits_uop_ctrl_is_std),
    .io_lsu_lxcpt_bits_uop_ctrl_op3_sel(core_io_lsu_lxcpt_bits_uop_ctrl_op3_sel),
    .io_lsu_lxcpt_bits_uop_iw_state(core_io_lsu_lxcpt_bits_uop_iw_state),
    .io_lsu_lxcpt_bits_uop_iw_p1_poisoned(core_io_lsu_lxcpt_bits_uop_iw_p1_poisoned),
    .io_lsu_lxcpt_bits_uop_iw_p2_poisoned(core_io_lsu_lxcpt_bits_uop_iw_p2_poisoned),
    .io_lsu_lxcpt_bits_uop_is_br(core_io_lsu_lxcpt_bits_uop_is_br),
    .io_lsu_lxcpt_bits_uop_is_jalr(core_io_lsu_lxcpt_bits_uop_is_jalr),
    .io_lsu_lxcpt_bits_uop_is_jal(core_io_lsu_lxcpt_bits_uop_is_jal),
    .io_lsu_lxcpt_bits_uop_is_sfb(core_io_lsu_lxcpt_bits_uop_is_sfb),
    .io_lsu_lxcpt_bits_uop_br_mask(core_io_lsu_lxcpt_bits_uop_br_mask),
    .io_lsu_lxcpt_bits_uop_br_tag(core_io_lsu_lxcpt_bits_uop_br_tag),
    .io_lsu_lxcpt_bits_uop_ftq_idx(core_io_lsu_lxcpt_bits_uop_ftq_idx),
    .io_lsu_lxcpt_bits_uop_edge_inst(core_io_lsu_lxcpt_bits_uop_edge_inst),
    .io_lsu_lxcpt_bits_uop_pc_lob(core_io_lsu_lxcpt_bits_uop_pc_lob),
    .io_lsu_lxcpt_bits_uop_taken(core_io_lsu_lxcpt_bits_uop_taken),
    .io_lsu_lxcpt_bits_uop_imm_packed(core_io_lsu_lxcpt_bits_uop_imm_packed),
    .io_lsu_lxcpt_bits_uop_csr_addr(core_io_lsu_lxcpt_bits_uop_csr_addr),
    .io_lsu_lxcpt_bits_uop_rob_idx(core_io_lsu_lxcpt_bits_uop_rob_idx),
    .io_lsu_lxcpt_bits_uop_ldq_idx(core_io_lsu_lxcpt_bits_uop_ldq_idx),
    .io_lsu_lxcpt_bits_uop_stq_idx(core_io_lsu_lxcpt_bits_uop_stq_idx),
    .io_lsu_lxcpt_bits_uop_rxq_idx(core_io_lsu_lxcpt_bits_uop_rxq_idx),
    .io_lsu_lxcpt_bits_uop_pdst(core_io_lsu_lxcpt_bits_uop_pdst),
    .io_lsu_lxcpt_bits_uop_prs1(core_io_lsu_lxcpt_bits_uop_prs1),
    .io_lsu_lxcpt_bits_uop_prs2(core_io_lsu_lxcpt_bits_uop_prs2),
    .io_lsu_lxcpt_bits_uop_prs3(core_io_lsu_lxcpt_bits_uop_prs3),
    .io_lsu_lxcpt_bits_uop_ppred(core_io_lsu_lxcpt_bits_uop_ppred),
    .io_lsu_lxcpt_bits_uop_prs1_busy(core_io_lsu_lxcpt_bits_uop_prs1_busy),
    .io_lsu_lxcpt_bits_uop_prs2_busy(core_io_lsu_lxcpt_bits_uop_prs2_busy),
    .io_lsu_lxcpt_bits_uop_prs3_busy(core_io_lsu_lxcpt_bits_uop_prs3_busy),
    .io_lsu_lxcpt_bits_uop_ppred_busy(core_io_lsu_lxcpt_bits_uop_ppred_busy),
    .io_lsu_lxcpt_bits_uop_stale_pdst(core_io_lsu_lxcpt_bits_uop_stale_pdst),
    .io_lsu_lxcpt_bits_uop_exception(core_io_lsu_lxcpt_bits_uop_exception),
    .io_lsu_lxcpt_bits_uop_exc_cause(core_io_lsu_lxcpt_bits_uop_exc_cause),
    .io_lsu_lxcpt_bits_uop_bypassable(core_io_lsu_lxcpt_bits_uop_bypassable),
    .io_lsu_lxcpt_bits_uop_mem_cmd(core_io_lsu_lxcpt_bits_uop_mem_cmd),
    .io_lsu_lxcpt_bits_uop_mem_size(core_io_lsu_lxcpt_bits_uop_mem_size),
    .io_lsu_lxcpt_bits_uop_mem_signed(core_io_lsu_lxcpt_bits_uop_mem_signed),
    .io_lsu_lxcpt_bits_uop_is_fence(core_io_lsu_lxcpt_bits_uop_is_fence),
    .io_lsu_lxcpt_bits_uop_is_fencei(core_io_lsu_lxcpt_bits_uop_is_fencei),
    .io_lsu_lxcpt_bits_uop_is_amo(core_io_lsu_lxcpt_bits_uop_is_amo),
    .io_lsu_lxcpt_bits_uop_uses_ldq(core_io_lsu_lxcpt_bits_uop_uses_ldq),
    .io_lsu_lxcpt_bits_uop_uses_stq(core_io_lsu_lxcpt_bits_uop_uses_stq),
    .io_lsu_lxcpt_bits_uop_is_sys_pc2epc(core_io_lsu_lxcpt_bits_uop_is_sys_pc2epc),
    .io_lsu_lxcpt_bits_uop_is_unique(core_io_lsu_lxcpt_bits_uop_is_unique),
    .io_lsu_lxcpt_bits_uop_flush_on_commit(core_io_lsu_lxcpt_bits_uop_flush_on_commit),
    .io_lsu_lxcpt_bits_uop_ldst_is_rs1(core_io_lsu_lxcpt_bits_uop_ldst_is_rs1),
    .io_lsu_lxcpt_bits_uop_ldst(core_io_lsu_lxcpt_bits_uop_ldst),
    .io_lsu_lxcpt_bits_uop_lrs1(core_io_lsu_lxcpt_bits_uop_lrs1),
    .io_lsu_lxcpt_bits_uop_lrs2(core_io_lsu_lxcpt_bits_uop_lrs2),
    .io_lsu_lxcpt_bits_uop_lrs3(core_io_lsu_lxcpt_bits_uop_lrs3),
    .io_lsu_lxcpt_bits_uop_ldst_val(core_io_lsu_lxcpt_bits_uop_ldst_val),
    .io_lsu_lxcpt_bits_uop_dst_rtype(core_io_lsu_lxcpt_bits_uop_dst_rtype),
    .io_lsu_lxcpt_bits_uop_lrs1_rtype(core_io_lsu_lxcpt_bits_uop_lrs1_rtype),
    .io_lsu_lxcpt_bits_uop_lrs2_rtype(core_io_lsu_lxcpt_bits_uop_lrs2_rtype),
    .io_lsu_lxcpt_bits_uop_frs3_en(core_io_lsu_lxcpt_bits_uop_frs3_en),
    .io_lsu_lxcpt_bits_uop_fp_val(core_io_lsu_lxcpt_bits_uop_fp_val),
    .io_lsu_lxcpt_bits_uop_fp_single(core_io_lsu_lxcpt_bits_uop_fp_single),
    .io_lsu_lxcpt_bits_uop_xcpt_pf_if(core_io_lsu_lxcpt_bits_uop_xcpt_pf_if),
    .io_lsu_lxcpt_bits_uop_xcpt_ae_if(core_io_lsu_lxcpt_bits_uop_xcpt_ae_if),
    .io_lsu_lxcpt_bits_uop_xcpt_ma_if(core_io_lsu_lxcpt_bits_uop_xcpt_ma_if),
    .io_lsu_lxcpt_bits_uop_bp_debug_if(core_io_lsu_lxcpt_bits_uop_bp_debug_if),
    .io_lsu_lxcpt_bits_uop_bp_xcpt_if(core_io_lsu_lxcpt_bits_uop_bp_xcpt_if),
    .io_lsu_lxcpt_bits_uop_debug_fsrc(core_io_lsu_lxcpt_bits_uop_debug_fsrc),
    .io_lsu_lxcpt_bits_uop_debug_tsrc(core_io_lsu_lxcpt_bits_uop_debug_tsrc),
    .io_lsu_lxcpt_bits_cause(core_io_lsu_lxcpt_bits_cause),
    .io_lsu_lxcpt_bits_badvaddr(core_io_lsu_lxcpt_bits_badvaddr),
    .io_lsu_tsc_reg(core_io_lsu_tsc_reg),
    .io_lsu_perf_acquire(core_io_lsu_perf_acquire),
    .io_lsu_perf_release(core_io_lsu_perf_release),
    .io_lsu_perf_tlbMiss(core_io_lsu_perf_tlbMiss),
    .io_ptw_tlb_req_ready(core_io_ptw_tlb_req_ready),
    .io_ptw_tlb_req_valid(core_io_ptw_tlb_req_valid),
    .io_ptw_tlb_req_bits_valid(core_io_ptw_tlb_req_bits_valid),
    .io_ptw_tlb_req_bits_bits_addr(core_io_ptw_tlb_req_bits_bits_addr),
    .io_ptw_tlb_resp_valid(core_io_ptw_tlb_resp_valid),
    .io_ptw_tlb_resp_bits_ae(core_io_ptw_tlb_resp_bits_ae),
    .io_ptw_tlb_resp_bits_pte_ppn(core_io_ptw_tlb_resp_bits_pte_ppn),
    .io_ptw_tlb_resp_bits_pte_reserved_for_software(core_io_ptw_tlb_resp_bits_pte_reserved_for_software),
    .io_ptw_tlb_resp_bits_pte_d(core_io_ptw_tlb_resp_bits_pte_d),
    .io_ptw_tlb_resp_bits_pte_a(core_io_ptw_tlb_resp_bits_pte_a),
    .io_ptw_tlb_resp_bits_pte_g(core_io_ptw_tlb_resp_bits_pte_g),
    .io_ptw_tlb_resp_bits_pte_u(core_io_ptw_tlb_resp_bits_pte_u),
    .io_ptw_tlb_resp_bits_pte_x(core_io_ptw_tlb_resp_bits_pte_x),
    .io_ptw_tlb_resp_bits_pte_w(core_io_ptw_tlb_resp_bits_pte_w),
    .io_ptw_tlb_resp_bits_pte_r(core_io_ptw_tlb_resp_bits_pte_r),
    .io_ptw_tlb_resp_bits_pte_v(core_io_ptw_tlb_resp_bits_pte_v),
    .io_ptw_tlb_resp_bits_level(core_io_ptw_tlb_resp_bits_level),
    .io_ptw_tlb_resp_bits_fragmented_superpage(core_io_ptw_tlb_resp_bits_fragmented_superpage),
    .io_ptw_tlb_resp_bits_homogeneous(core_io_ptw_tlb_resp_bits_homogeneous),
    .io_ptw_tlb_ptbr_mode(core_io_ptw_tlb_ptbr_mode),
    .io_ptw_tlb_ptbr_asid(core_io_ptw_tlb_ptbr_asid),
    .io_ptw_tlb_ptbr_ppn(core_io_ptw_tlb_ptbr_ppn),
    .io_ptw_tlb_status_debug(core_io_ptw_tlb_status_debug),
    .io_ptw_tlb_status_cease(core_io_ptw_tlb_status_cease),
    .io_ptw_tlb_status_wfi(core_io_ptw_tlb_status_wfi),
    .io_ptw_tlb_status_isa(core_io_ptw_tlb_status_isa),
    .io_ptw_tlb_status_dprv(core_io_ptw_tlb_status_dprv),
    .io_ptw_tlb_status_prv(core_io_ptw_tlb_status_prv),
    .io_ptw_tlb_status_sd(core_io_ptw_tlb_status_sd),
    .io_ptw_tlb_status_zero2(core_io_ptw_tlb_status_zero2),
    .io_ptw_tlb_status_sxl(core_io_ptw_tlb_status_sxl),
    .io_ptw_tlb_status_uxl(core_io_ptw_tlb_status_uxl),
    .io_ptw_tlb_status_sd_rv32(core_io_ptw_tlb_status_sd_rv32),
    .io_ptw_tlb_status_zero1(core_io_ptw_tlb_status_zero1),
    .io_ptw_tlb_status_tsr(core_io_ptw_tlb_status_tsr),
    .io_ptw_tlb_status_tw(core_io_ptw_tlb_status_tw),
    .io_ptw_tlb_status_tvm(core_io_ptw_tlb_status_tvm),
    .io_ptw_tlb_status_mxr(core_io_ptw_tlb_status_mxr),
    .io_ptw_tlb_status_sum(core_io_ptw_tlb_status_sum),
    .io_ptw_tlb_status_mprv(core_io_ptw_tlb_status_mprv),
    .io_ptw_tlb_status_xs(core_io_ptw_tlb_status_xs),
    .io_ptw_tlb_status_fs(core_io_ptw_tlb_status_fs),
    .io_ptw_tlb_status_mpp(core_io_ptw_tlb_status_mpp),
    .io_ptw_tlb_status_vs(core_io_ptw_tlb_status_vs),
    .io_ptw_tlb_status_spp(core_io_ptw_tlb_status_spp),
    .io_ptw_tlb_status_mpie(core_io_ptw_tlb_status_mpie),
    .io_ptw_tlb_status_hpie(core_io_ptw_tlb_status_hpie),
    .io_ptw_tlb_status_spie(core_io_ptw_tlb_status_spie),
    .io_ptw_tlb_status_upie(core_io_ptw_tlb_status_upie),
    .io_ptw_tlb_status_mie(core_io_ptw_tlb_status_mie),
    .io_ptw_tlb_status_hie(core_io_ptw_tlb_status_hie),
    .io_ptw_tlb_status_sie(core_io_ptw_tlb_status_sie),
    .io_ptw_tlb_status_uie(core_io_ptw_tlb_status_uie),
    .io_ptw_tlb_pmp_0_cfg_l(core_io_ptw_tlb_pmp_0_cfg_l),
    .io_ptw_tlb_pmp_0_cfg_res(core_io_ptw_tlb_pmp_0_cfg_res),
    .io_ptw_tlb_pmp_0_cfg_a(core_io_ptw_tlb_pmp_0_cfg_a),
    .io_ptw_tlb_pmp_0_cfg_x(core_io_ptw_tlb_pmp_0_cfg_x),
    .io_ptw_tlb_pmp_0_cfg_w(core_io_ptw_tlb_pmp_0_cfg_w),
    .io_ptw_tlb_pmp_0_cfg_r(core_io_ptw_tlb_pmp_0_cfg_r),
    .io_ptw_tlb_pmp_0_addr(core_io_ptw_tlb_pmp_0_addr),
    .io_ptw_tlb_pmp_0_mask(core_io_ptw_tlb_pmp_0_mask),
    .io_ptw_tlb_pmp_1_cfg_l(core_io_ptw_tlb_pmp_1_cfg_l),
    .io_ptw_tlb_pmp_1_cfg_res(core_io_ptw_tlb_pmp_1_cfg_res),
    .io_ptw_tlb_pmp_1_cfg_a(core_io_ptw_tlb_pmp_1_cfg_a),
    .io_ptw_tlb_pmp_1_cfg_x(core_io_ptw_tlb_pmp_1_cfg_x),
    .io_ptw_tlb_pmp_1_cfg_w(core_io_ptw_tlb_pmp_1_cfg_w),
    .io_ptw_tlb_pmp_1_cfg_r(core_io_ptw_tlb_pmp_1_cfg_r),
    .io_ptw_tlb_pmp_1_addr(core_io_ptw_tlb_pmp_1_addr),
    .io_ptw_tlb_pmp_1_mask(core_io_ptw_tlb_pmp_1_mask),
    .io_ptw_tlb_pmp_2_cfg_l(core_io_ptw_tlb_pmp_2_cfg_l),
    .io_ptw_tlb_pmp_2_cfg_res(core_io_ptw_tlb_pmp_2_cfg_res),
    .io_ptw_tlb_pmp_2_cfg_a(core_io_ptw_tlb_pmp_2_cfg_a),
    .io_ptw_tlb_pmp_2_cfg_x(core_io_ptw_tlb_pmp_2_cfg_x),
    .io_ptw_tlb_pmp_2_cfg_w(core_io_ptw_tlb_pmp_2_cfg_w),
    .io_ptw_tlb_pmp_2_cfg_r(core_io_ptw_tlb_pmp_2_cfg_r),
    .io_ptw_tlb_pmp_2_addr(core_io_ptw_tlb_pmp_2_addr),
    .io_ptw_tlb_pmp_2_mask(core_io_ptw_tlb_pmp_2_mask),
    .io_ptw_tlb_pmp_3_cfg_l(core_io_ptw_tlb_pmp_3_cfg_l),
    .io_ptw_tlb_pmp_3_cfg_res(core_io_ptw_tlb_pmp_3_cfg_res),
    .io_ptw_tlb_pmp_3_cfg_a(core_io_ptw_tlb_pmp_3_cfg_a),
    .io_ptw_tlb_pmp_3_cfg_x(core_io_ptw_tlb_pmp_3_cfg_x),
    .io_ptw_tlb_pmp_3_cfg_w(core_io_ptw_tlb_pmp_3_cfg_w),
    .io_ptw_tlb_pmp_3_cfg_r(core_io_ptw_tlb_pmp_3_cfg_r),
    .io_ptw_tlb_pmp_3_addr(core_io_ptw_tlb_pmp_3_addr),
    .io_ptw_tlb_pmp_3_mask(core_io_ptw_tlb_pmp_3_mask),
    .io_ptw_tlb_pmp_4_cfg_l(core_io_ptw_tlb_pmp_4_cfg_l),
    .io_ptw_tlb_pmp_4_cfg_res(core_io_ptw_tlb_pmp_4_cfg_res),
    .io_ptw_tlb_pmp_4_cfg_a(core_io_ptw_tlb_pmp_4_cfg_a),
    .io_ptw_tlb_pmp_4_cfg_x(core_io_ptw_tlb_pmp_4_cfg_x),
    .io_ptw_tlb_pmp_4_cfg_w(core_io_ptw_tlb_pmp_4_cfg_w),
    .io_ptw_tlb_pmp_4_cfg_r(core_io_ptw_tlb_pmp_4_cfg_r),
    .io_ptw_tlb_pmp_4_addr(core_io_ptw_tlb_pmp_4_addr),
    .io_ptw_tlb_pmp_4_mask(core_io_ptw_tlb_pmp_4_mask),
    .io_ptw_tlb_pmp_5_cfg_l(core_io_ptw_tlb_pmp_5_cfg_l),
    .io_ptw_tlb_pmp_5_cfg_res(core_io_ptw_tlb_pmp_5_cfg_res),
    .io_ptw_tlb_pmp_5_cfg_a(core_io_ptw_tlb_pmp_5_cfg_a),
    .io_ptw_tlb_pmp_5_cfg_x(core_io_ptw_tlb_pmp_5_cfg_x),
    .io_ptw_tlb_pmp_5_cfg_w(core_io_ptw_tlb_pmp_5_cfg_w),
    .io_ptw_tlb_pmp_5_cfg_r(core_io_ptw_tlb_pmp_5_cfg_r),
    .io_ptw_tlb_pmp_5_addr(core_io_ptw_tlb_pmp_5_addr),
    .io_ptw_tlb_pmp_5_mask(core_io_ptw_tlb_pmp_5_mask),
    .io_ptw_tlb_pmp_6_cfg_l(core_io_ptw_tlb_pmp_6_cfg_l),
    .io_ptw_tlb_pmp_6_cfg_res(core_io_ptw_tlb_pmp_6_cfg_res),
    .io_ptw_tlb_pmp_6_cfg_a(core_io_ptw_tlb_pmp_6_cfg_a),
    .io_ptw_tlb_pmp_6_cfg_x(core_io_ptw_tlb_pmp_6_cfg_x),
    .io_ptw_tlb_pmp_6_cfg_w(core_io_ptw_tlb_pmp_6_cfg_w),
    .io_ptw_tlb_pmp_6_cfg_r(core_io_ptw_tlb_pmp_6_cfg_r),
    .io_ptw_tlb_pmp_6_addr(core_io_ptw_tlb_pmp_6_addr),
    .io_ptw_tlb_pmp_6_mask(core_io_ptw_tlb_pmp_6_mask),
    .io_ptw_tlb_pmp_7_cfg_l(core_io_ptw_tlb_pmp_7_cfg_l),
    .io_ptw_tlb_pmp_7_cfg_res(core_io_ptw_tlb_pmp_7_cfg_res),
    .io_ptw_tlb_pmp_7_cfg_a(core_io_ptw_tlb_pmp_7_cfg_a),
    .io_ptw_tlb_pmp_7_cfg_x(core_io_ptw_tlb_pmp_7_cfg_x),
    .io_ptw_tlb_pmp_7_cfg_w(core_io_ptw_tlb_pmp_7_cfg_w),
    .io_ptw_tlb_pmp_7_cfg_r(core_io_ptw_tlb_pmp_7_cfg_r),
    .io_ptw_tlb_pmp_7_addr(core_io_ptw_tlb_pmp_7_addr),
    .io_ptw_tlb_pmp_7_mask(core_io_ptw_tlb_pmp_7_mask),
    .io_ptw_tlb_customCSRs_csrs_0_wen(core_io_ptw_tlb_customCSRs_csrs_0_wen),
    .io_ptw_tlb_customCSRs_csrs_0_wdata(core_io_ptw_tlb_customCSRs_csrs_0_wdata),
    .io_ptw_tlb_customCSRs_csrs_0_value(core_io_ptw_tlb_customCSRs_csrs_0_value),
    .io_trace_0_valid(core_io_trace_0_valid),
    .io_trace_0_iaddr(core_io_trace_0_iaddr),
    .io_trace_0_insn(core_io_trace_0_insn),
    .io_trace_0_priv(core_io_trace_0_priv),
    .io_trace_0_exception(core_io_trace_0_exception),
    .io_trace_0_interrupt(core_io_trace_0_interrupt),
    .io_trace_0_cause(core_io_trace_0_cause),
    .io_trace_0_tval(core_io_trace_0_tval),
    .io_trace_0_wdata(core_io_trace_0_wdata),
    .io_trace_1_valid(core_io_trace_1_valid),
    .io_trace_1_iaddr(core_io_trace_1_iaddr),
    .io_trace_1_insn(core_io_trace_1_insn),
    .io_trace_1_priv(core_io_trace_1_priv),
    .io_trace_1_exception(core_io_trace_1_exception),
    .io_trace_1_interrupt(core_io_trace_1_interrupt),
    .io_trace_1_cause(core_io_trace_1_cause),
    .io_trace_1_tval(core_io_trace_1_tval),
    .io_trace_1_wdata(core_io_trace_1_wdata),
    .io_fcsr_rm(core_io_fcsr_rm)
  );
  LSU lsu ( // @[tile.scala 160:20]
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io_ptw_req_ready(lsu_io_ptw_req_ready),
    .io_ptw_req_valid(lsu_io_ptw_req_valid),
    .io_ptw_req_bits_valid(lsu_io_ptw_req_bits_valid),
    .io_ptw_req_bits_bits_addr(lsu_io_ptw_req_bits_bits_addr),
    .io_ptw_resp_valid(lsu_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae(lsu_io_ptw_resp_bits_ae),
    .io_ptw_resp_bits_pte_ppn(lsu_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(lsu_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(lsu_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(lsu_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(lsu_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(lsu_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(lsu_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(lsu_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(lsu_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(lsu_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(lsu_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_fragmented_superpage(lsu_io_ptw_resp_bits_fragmented_superpage),
    .io_ptw_resp_bits_homogeneous(lsu_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(lsu_io_ptw_ptbr_mode),
    .io_ptw_ptbr_asid(lsu_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(lsu_io_ptw_ptbr_ppn),
    .io_ptw_status_debug(lsu_io_ptw_status_debug),
    .io_ptw_status_cease(lsu_io_ptw_status_cease),
    .io_ptw_status_wfi(lsu_io_ptw_status_wfi),
    .io_ptw_status_isa(lsu_io_ptw_status_isa),
    .io_ptw_status_dprv(lsu_io_ptw_status_dprv),
    .io_ptw_status_prv(lsu_io_ptw_status_prv),
    .io_ptw_status_sd(lsu_io_ptw_status_sd),
    .io_ptw_status_zero2(lsu_io_ptw_status_zero2),
    .io_ptw_status_sxl(lsu_io_ptw_status_sxl),
    .io_ptw_status_uxl(lsu_io_ptw_status_uxl),
    .io_ptw_status_sd_rv32(lsu_io_ptw_status_sd_rv32),
    .io_ptw_status_zero1(lsu_io_ptw_status_zero1),
    .io_ptw_status_tsr(lsu_io_ptw_status_tsr),
    .io_ptw_status_tw(lsu_io_ptw_status_tw),
    .io_ptw_status_tvm(lsu_io_ptw_status_tvm),
    .io_ptw_status_mxr(lsu_io_ptw_status_mxr),
    .io_ptw_status_sum(lsu_io_ptw_status_sum),
    .io_ptw_status_mprv(lsu_io_ptw_status_mprv),
    .io_ptw_status_xs(lsu_io_ptw_status_xs),
    .io_ptw_status_fs(lsu_io_ptw_status_fs),
    .io_ptw_status_mpp(lsu_io_ptw_status_mpp),
    .io_ptw_status_vs(lsu_io_ptw_status_vs),
    .io_ptw_status_spp(lsu_io_ptw_status_spp),
    .io_ptw_status_mpie(lsu_io_ptw_status_mpie),
    .io_ptw_status_hpie(lsu_io_ptw_status_hpie),
    .io_ptw_status_spie(lsu_io_ptw_status_spie),
    .io_ptw_status_upie(lsu_io_ptw_status_upie),
    .io_ptw_status_mie(lsu_io_ptw_status_mie),
    .io_ptw_status_hie(lsu_io_ptw_status_hie),
    .io_ptw_status_sie(lsu_io_ptw_status_sie),
    .io_ptw_status_uie(lsu_io_ptw_status_uie),
    .io_ptw_pmp_0_cfg_l(lsu_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_res(lsu_io_ptw_pmp_0_cfg_res),
    .io_ptw_pmp_0_cfg_a(lsu_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(lsu_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(lsu_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(lsu_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(lsu_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(lsu_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(lsu_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_res(lsu_io_ptw_pmp_1_cfg_res),
    .io_ptw_pmp_1_cfg_a(lsu_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(lsu_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(lsu_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(lsu_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(lsu_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(lsu_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(lsu_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_res(lsu_io_ptw_pmp_2_cfg_res),
    .io_ptw_pmp_2_cfg_a(lsu_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(lsu_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(lsu_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(lsu_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(lsu_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(lsu_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(lsu_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_res(lsu_io_ptw_pmp_3_cfg_res),
    .io_ptw_pmp_3_cfg_a(lsu_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(lsu_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(lsu_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(lsu_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(lsu_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(lsu_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(lsu_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_res(lsu_io_ptw_pmp_4_cfg_res),
    .io_ptw_pmp_4_cfg_a(lsu_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(lsu_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(lsu_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(lsu_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(lsu_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(lsu_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(lsu_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_res(lsu_io_ptw_pmp_5_cfg_res),
    .io_ptw_pmp_5_cfg_a(lsu_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(lsu_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(lsu_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(lsu_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(lsu_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(lsu_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(lsu_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_res(lsu_io_ptw_pmp_6_cfg_res),
    .io_ptw_pmp_6_cfg_a(lsu_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(lsu_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(lsu_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(lsu_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(lsu_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(lsu_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(lsu_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_res(lsu_io_ptw_pmp_7_cfg_res),
    .io_ptw_pmp_7_cfg_a(lsu_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(lsu_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(lsu_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(lsu_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(lsu_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(lsu_io_ptw_pmp_7_mask),
    .io_ptw_customCSRs_csrs_0_wen(lsu_io_ptw_customCSRs_csrs_0_wen),
    .io_ptw_customCSRs_csrs_0_wdata(lsu_io_ptw_customCSRs_csrs_0_wdata),
    .io_ptw_customCSRs_csrs_0_value(lsu_io_ptw_customCSRs_csrs_0_value),
    .io_core_exe_0_req_valid(lsu_io_core_exe_0_req_valid),
    .io_core_exe_0_req_bits_uop_switch(lsu_io_core_exe_0_req_bits_uop_switch),
    .io_core_exe_0_req_bits_uop_switch_off(lsu_io_core_exe_0_req_bits_uop_switch_off),
    .io_core_exe_0_req_bits_uop_is_unicore(lsu_io_core_exe_0_req_bits_uop_is_unicore),
    .io_core_exe_0_req_bits_uop_shift(lsu_io_core_exe_0_req_bits_uop_shift),
    .io_core_exe_0_req_bits_uop_lrs3_rtype(lsu_io_core_exe_0_req_bits_uop_lrs3_rtype),
    .io_core_exe_0_req_bits_uop_rflag(lsu_io_core_exe_0_req_bits_uop_rflag),
    .io_core_exe_0_req_bits_uop_wflag(lsu_io_core_exe_0_req_bits_uop_wflag),
    .io_core_exe_0_req_bits_uop_prflag(lsu_io_core_exe_0_req_bits_uop_prflag),
    .io_core_exe_0_req_bits_uop_pwflag(lsu_io_core_exe_0_req_bits_uop_pwflag),
    .io_core_exe_0_req_bits_uop_pflag_busy(lsu_io_core_exe_0_req_bits_uop_pflag_busy),
    .io_core_exe_0_req_bits_uop_stale_pflag(lsu_io_core_exe_0_req_bits_uop_stale_pflag),
    .io_core_exe_0_req_bits_uop_op1_sel(lsu_io_core_exe_0_req_bits_uop_op1_sel),
    .io_core_exe_0_req_bits_uop_op2_sel(lsu_io_core_exe_0_req_bits_uop_op2_sel),
    .io_core_exe_0_req_bits_uop_split_num(lsu_io_core_exe_0_req_bits_uop_split_num),
    .io_core_exe_0_req_bits_uop_self_index(lsu_io_core_exe_0_req_bits_uop_self_index),
    .io_core_exe_0_req_bits_uop_rob_inst_idx(lsu_io_core_exe_0_req_bits_uop_rob_inst_idx),
    .io_core_exe_0_req_bits_uop_address_num(lsu_io_core_exe_0_req_bits_uop_address_num),
    .io_core_exe_0_req_bits_uop_uopc(lsu_io_core_exe_0_req_bits_uop_uopc),
    .io_core_exe_0_req_bits_uop_inst(lsu_io_core_exe_0_req_bits_uop_inst),
    .io_core_exe_0_req_bits_uop_debug_inst(lsu_io_core_exe_0_req_bits_uop_debug_inst),
    .io_core_exe_0_req_bits_uop_is_rvc(lsu_io_core_exe_0_req_bits_uop_is_rvc),
    .io_core_exe_0_req_bits_uop_debug_pc(lsu_io_core_exe_0_req_bits_uop_debug_pc),
    .io_core_exe_0_req_bits_uop_iq_type(lsu_io_core_exe_0_req_bits_uop_iq_type),
    .io_core_exe_0_req_bits_uop_fu_code(lsu_io_core_exe_0_req_bits_uop_fu_code),
    .io_core_exe_0_req_bits_uop_ctrl_br_type(lsu_io_core_exe_0_req_bits_uop_ctrl_br_type),
    .io_core_exe_0_req_bits_uop_ctrl_op1_sel(lsu_io_core_exe_0_req_bits_uop_ctrl_op1_sel),
    .io_core_exe_0_req_bits_uop_ctrl_op2_sel(lsu_io_core_exe_0_req_bits_uop_ctrl_op2_sel),
    .io_core_exe_0_req_bits_uop_ctrl_imm_sel(lsu_io_core_exe_0_req_bits_uop_ctrl_imm_sel),
    .io_core_exe_0_req_bits_uop_ctrl_op_fcn(lsu_io_core_exe_0_req_bits_uop_ctrl_op_fcn),
    .io_core_exe_0_req_bits_uop_ctrl_fcn_dw(lsu_io_core_exe_0_req_bits_uop_ctrl_fcn_dw),
    .io_core_exe_0_req_bits_uop_ctrl_csr_cmd(lsu_io_core_exe_0_req_bits_uop_ctrl_csr_cmd),
    .io_core_exe_0_req_bits_uop_ctrl_is_load(lsu_io_core_exe_0_req_bits_uop_ctrl_is_load),
    .io_core_exe_0_req_bits_uop_ctrl_is_sta(lsu_io_core_exe_0_req_bits_uop_ctrl_is_sta),
    .io_core_exe_0_req_bits_uop_ctrl_is_std(lsu_io_core_exe_0_req_bits_uop_ctrl_is_std),
    .io_core_exe_0_req_bits_uop_ctrl_op3_sel(lsu_io_core_exe_0_req_bits_uop_ctrl_op3_sel),
    .io_core_exe_0_req_bits_uop_iw_state(lsu_io_core_exe_0_req_bits_uop_iw_state),
    .io_core_exe_0_req_bits_uop_iw_p1_poisoned(lsu_io_core_exe_0_req_bits_uop_iw_p1_poisoned),
    .io_core_exe_0_req_bits_uop_iw_p2_poisoned(lsu_io_core_exe_0_req_bits_uop_iw_p2_poisoned),
    .io_core_exe_0_req_bits_uop_is_br(lsu_io_core_exe_0_req_bits_uop_is_br),
    .io_core_exe_0_req_bits_uop_is_jalr(lsu_io_core_exe_0_req_bits_uop_is_jalr),
    .io_core_exe_0_req_bits_uop_is_jal(lsu_io_core_exe_0_req_bits_uop_is_jal),
    .io_core_exe_0_req_bits_uop_is_sfb(lsu_io_core_exe_0_req_bits_uop_is_sfb),
    .io_core_exe_0_req_bits_uop_br_mask(lsu_io_core_exe_0_req_bits_uop_br_mask),
    .io_core_exe_0_req_bits_uop_br_tag(lsu_io_core_exe_0_req_bits_uop_br_tag),
    .io_core_exe_0_req_bits_uop_ftq_idx(lsu_io_core_exe_0_req_bits_uop_ftq_idx),
    .io_core_exe_0_req_bits_uop_edge_inst(lsu_io_core_exe_0_req_bits_uop_edge_inst),
    .io_core_exe_0_req_bits_uop_pc_lob(lsu_io_core_exe_0_req_bits_uop_pc_lob),
    .io_core_exe_0_req_bits_uop_taken(lsu_io_core_exe_0_req_bits_uop_taken),
    .io_core_exe_0_req_bits_uop_imm_packed(lsu_io_core_exe_0_req_bits_uop_imm_packed),
    .io_core_exe_0_req_bits_uop_csr_addr(lsu_io_core_exe_0_req_bits_uop_csr_addr),
    .io_core_exe_0_req_bits_uop_rob_idx(lsu_io_core_exe_0_req_bits_uop_rob_idx),
    .io_core_exe_0_req_bits_uop_ldq_idx(lsu_io_core_exe_0_req_bits_uop_ldq_idx),
    .io_core_exe_0_req_bits_uop_stq_idx(lsu_io_core_exe_0_req_bits_uop_stq_idx),
    .io_core_exe_0_req_bits_uop_rxq_idx(lsu_io_core_exe_0_req_bits_uop_rxq_idx),
    .io_core_exe_0_req_bits_uop_pdst(lsu_io_core_exe_0_req_bits_uop_pdst),
    .io_core_exe_0_req_bits_uop_prs1(lsu_io_core_exe_0_req_bits_uop_prs1),
    .io_core_exe_0_req_bits_uop_prs2(lsu_io_core_exe_0_req_bits_uop_prs2),
    .io_core_exe_0_req_bits_uop_prs3(lsu_io_core_exe_0_req_bits_uop_prs3),
    .io_core_exe_0_req_bits_uop_ppred(lsu_io_core_exe_0_req_bits_uop_ppred),
    .io_core_exe_0_req_bits_uop_prs1_busy(lsu_io_core_exe_0_req_bits_uop_prs1_busy),
    .io_core_exe_0_req_bits_uop_prs2_busy(lsu_io_core_exe_0_req_bits_uop_prs2_busy),
    .io_core_exe_0_req_bits_uop_prs3_busy(lsu_io_core_exe_0_req_bits_uop_prs3_busy),
    .io_core_exe_0_req_bits_uop_ppred_busy(lsu_io_core_exe_0_req_bits_uop_ppred_busy),
    .io_core_exe_0_req_bits_uop_stale_pdst(lsu_io_core_exe_0_req_bits_uop_stale_pdst),
    .io_core_exe_0_req_bits_uop_exception(lsu_io_core_exe_0_req_bits_uop_exception),
    .io_core_exe_0_req_bits_uop_exc_cause(lsu_io_core_exe_0_req_bits_uop_exc_cause),
    .io_core_exe_0_req_bits_uop_bypassable(lsu_io_core_exe_0_req_bits_uop_bypassable),
    .io_core_exe_0_req_bits_uop_mem_cmd(lsu_io_core_exe_0_req_bits_uop_mem_cmd),
    .io_core_exe_0_req_bits_uop_mem_size(lsu_io_core_exe_0_req_bits_uop_mem_size),
    .io_core_exe_0_req_bits_uop_mem_signed(lsu_io_core_exe_0_req_bits_uop_mem_signed),
    .io_core_exe_0_req_bits_uop_is_fence(lsu_io_core_exe_0_req_bits_uop_is_fence),
    .io_core_exe_0_req_bits_uop_is_fencei(lsu_io_core_exe_0_req_bits_uop_is_fencei),
    .io_core_exe_0_req_bits_uop_is_amo(lsu_io_core_exe_0_req_bits_uop_is_amo),
    .io_core_exe_0_req_bits_uop_uses_ldq(lsu_io_core_exe_0_req_bits_uop_uses_ldq),
    .io_core_exe_0_req_bits_uop_uses_stq(lsu_io_core_exe_0_req_bits_uop_uses_stq),
    .io_core_exe_0_req_bits_uop_is_sys_pc2epc(lsu_io_core_exe_0_req_bits_uop_is_sys_pc2epc),
    .io_core_exe_0_req_bits_uop_is_unique(lsu_io_core_exe_0_req_bits_uop_is_unique),
    .io_core_exe_0_req_bits_uop_flush_on_commit(lsu_io_core_exe_0_req_bits_uop_flush_on_commit),
    .io_core_exe_0_req_bits_uop_ldst_is_rs1(lsu_io_core_exe_0_req_bits_uop_ldst_is_rs1),
    .io_core_exe_0_req_bits_uop_ldst(lsu_io_core_exe_0_req_bits_uop_ldst),
    .io_core_exe_0_req_bits_uop_lrs1(lsu_io_core_exe_0_req_bits_uop_lrs1),
    .io_core_exe_0_req_bits_uop_lrs2(lsu_io_core_exe_0_req_bits_uop_lrs2),
    .io_core_exe_0_req_bits_uop_lrs3(lsu_io_core_exe_0_req_bits_uop_lrs3),
    .io_core_exe_0_req_bits_uop_ldst_val(lsu_io_core_exe_0_req_bits_uop_ldst_val),
    .io_core_exe_0_req_bits_uop_dst_rtype(lsu_io_core_exe_0_req_bits_uop_dst_rtype),
    .io_core_exe_0_req_bits_uop_lrs1_rtype(lsu_io_core_exe_0_req_bits_uop_lrs1_rtype),
    .io_core_exe_0_req_bits_uop_lrs2_rtype(lsu_io_core_exe_0_req_bits_uop_lrs2_rtype),
    .io_core_exe_0_req_bits_uop_frs3_en(lsu_io_core_exe_0_req_bits_uop_frs3_en),
    .io_core_exe_0_req_bits_uop_fp_val(lsu_io_core_exe_0_req_bits_uop_fp_val),
    .io_core_exe_0_req_bits_uop_fp_single(lsu_io_core_exe_0_req_bits_uop_fp_single),
    .io_core_exe_0_req_bits_uop_xcpt_pf_if(lsu_io_core_exe_0_req_bits_uop_xcpt_pf_if),
    .io_core_exe_0_req_bits_uop_xcpt_ae_if(lsu_io_core_exe_0_req_bits_uop_xcpt_ae_if),
    .io_core_exe_0_req_bits_uop_xcpt_ma_if(lsu_io_core_exe_0_req_bits_uop_xcpt_ma_if),
    .io_core_exe_0_req_bits_uop_bp_debug_if(lsu_io_core_exe_0_req_bits_uop_bp_debug_if),
    .io_core_exe_0_req_bits_uop_bp_xcpt_if(lsu_io_core_exe_0_req_bits_uop_bp_xcpt_if),
    .io_core_exe_0_req_bits_uop_debug_fsrc(lsu_io_core_exe_0_req_bits_uop_debug_fsrc),
    .io_core_exe_0_req_bits_uop_debug_tsrc(lsu_io_core_exe_0_req_bits_uop_debug_tsrc),
    .io_core_exe_0_req_bits_predicated(lsu_io_core_exe_0_req_bits_predicated),
    .io_core_exe_0_req_bits_data(lsu_io_core_exe_0_req_bits_data),
    .io_core_exe_0_req_bits_fflags_valid(lsu_io_core_exe_0_req_bits_fflags_valid),
    .io_core_exe_0_req_bits_fflags_bits_uop_switch(lsu_io_core_exe_0_req_bits_fflags_bits_uop_switch),
    .io_core_exe_0_req_bits_fflags_bits_uop_switch_off(lsu_io_core_exe_0_req_bits_fflags_bits_uop_switch_off),
    .io_core_exe_0_req_bits_fflags_bits_uop_is_unicore(lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_unicore),
    .io_core_exe_0_req_bits_fflags_bits_uop_shift(lsu_io_core_exe_0_req_bits_fflags_bits_uop_shift),
    .io_core_exe_0_req_bits_fflags_bits_uop_lrs3_rtype(lsu_io_core_exe_0_req_bits_fflags_bits_uop_lrs3_rtype),
    .io_core_exe_0_req_bits_fflags_bits_uop_rflag(lsu_io_core_exe_0_req_bits_fflags_bits_uop_rflag),
    .io_core_exe_0_req_bits_fflags_bits_uop_wflag(lsu_io_core_exe_0_req_bits_fflags_bits_uop_wflag),
    .io_core_exe_0_req_bits_fflags_bits_uop_prflag(lsu_io_core_exe_0_req_bits_fflags_bits_uop_prflag),
    .io_core_exe_0_req_bits_fflags_bits_uop_pwflag(lsu_io_core_exe_0_req_bits_fflags_bits_uop_pwflag),
    .io_core_exe_0_req_bits_fflags_bits_uop_pflag_busy(lsu_io_core_exe_0_req_bits_fflags_bits_uop_pflag_busy),
    .io_core_exe_0_req_bits_fflags_bits_uop_stale_pflag(lsu_io_core_exe_0_req_bits_fflags_bits_uop_stale_pflag),
    .io_core_exe_0_req_bits_fflags_bits_uop_op1_sel(lsu_io_core_exe_0_req_bits_fflags_bits_uop_op1_sel),
    .io_core_exe_0_req_bits_fflags_bits_uop_op2_sel(lsu_io_core_exe_0_req_bits_fflags_bits_uop_op2_sel),
    .io_core_exe_0_req_bits_fflags_bits_uop_split_num(lsu_io_core_exe_0_req_bits_fflags_bits_uop_split_num),
    .io_core_exe_0_req_bits_fflags_bits_uop_self_index(lsu_io_core_exe_0_req_bits_fflags_bits_uop_self_index),
    .io_core_exe_0_req_bits_fflags_bits_uop_rob_inst_idx(lsu_io_core_exe_0_req_bits_fflags_bits_uop_rob_inst_idx),
    .io_core_exe_0_req_bits_fflags_bits_uop_address_num(lsu_io_core_exe_0_req_bits_fflags_bits_uop_address_num),
    .io_core_exe_0_req_bits_fflags_bits_uop_uopc(lsu_io_core_exe_0_req_bits_fflags_bits_uop_uopc),
    .io_core_exe_0_req_bits_fflags_bits_uop_inst(lsu_io_core_exe_0_req_bits_fflags_bits_uop_inst),
    .io_core_exe_0_req_bits_fflags_bits_uop_debug_inst(lsu_io_core_exe_0_req_bits_fflags_bits_uop_debug_inst),
    .io_core_exe_0_req_bits_fflags_bits_uop_is_rvc(lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_rvc),
    .io_core_exe_0_req_bits_fflags_bits_uop_debug_pc(lsu_io_core_exe_0_req_bits_fflags_bits_uop_debug_pc),
    .io_core_exe_0_req_bits_fflags_bits_uop_iq_type(lsu_io_core_exe_0_req_bits_fflags_bits_uop_iq_type),
    .io_core_exe_0_req_bits_fflags_bits_uop_fu_code(lsu_io_core_exe_0_req_bits_fflags_bits_uop_fu_code),
    .io_core_exe_0_req_bits_fflags_bits_uop_ctrl_br_type(lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_br_type),
    .io_core_exe_0_req_bits_fflags_bits_uop_ctrl_op1_sel(lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_op1_sel),
    .io_core_exe_0_req_bits_fflags_bits_uop_ctrl_op2_sel(lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_op2_sel),
    .io_core_exe_0_req_bits_fflags_bits_uop_ctrl_imm_sel(lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_imm_sel),
    .io_core_exe_0_req_bits_fflags_bits_uop_ctrl_op_fcn(lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_op_fcn),
    .io_core_exe_0_req_bits_fflags_bits_uop_ctrl_fcn_dw(lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_fcn_dw),
    .io_core_exe_0_req_bits_fflags_bits_uop_ctrl_csr_cmd(lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_csr_cmd),
    .io_core_exe_0_req_bits_fflags_bits_uop_ctrl_is_load(lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_is_load),
    .io_core_exe_0_req_bits_fflags_bits_uop_ctrl_is_sta(lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_is_sta),
    .io_core_exe_0_req_bits_fflags_bits_uop_ctrl_is_std(lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_is_std),
    .io_core_exe_0_req_bits_fflags_bits_uop_ctrl_op3_sel(lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_op3_sel),
    .io_core_exe_0_req_bits_fflags_bits_uop_iw_state(lsu_io_core_exe_0_req_bits_fflags_bits_uop_iw_state),
    .io_core_exe_0_req_bits_fflags_bits_uop_iw_p1_poisoned(lsu_io_core_exe_0_req_bits_fflags_bits_uop_iw_p1_poisoned),
    .io_core_exe_0_req_bits_fflags_bits_uop_iw_p2_poisoned(lsu_io_core_exe_0_req_bits_fflags_bits_uop_iw_p2_poisoned),
    .io_core_exe_0_req_bits_fflags_bits_uop_is_br(lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_br),
    .io_core_exe_0_req_bits_fflags_bits_uop_is_jalr(lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_jalr),
    .io_core_exe_0_req_bits_fflags_bits_uop_is_jal(lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_jal),
    .io_core_exe_0_req_bits_fflags_bits_uop_is_sfb(lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_sfb),
    .io_core_exe_0_req_bits_fflags_bits_uop_br_mask(lsu_io_core_exe_0_req_bits_fflags_bits_uop_br_mask),
    .io_core_exe_0_req_bits_fflags_bits_uop_br_tag(lsu_io_core_exe_0_req_bits_fflags_bits_uop_br_tag),
    .io_core_exe_0_req_bits_fflags_bits_uop_ftq_idx(lsu_io_core_exe_0_req_bits_fflags_bits_uop_ftq_idx),
    .io_core_exe_0_req_bits_fflags_bits_uop_edge_inst(lsu_io_core_exe_0_req_bits_fflags_bits_uop_edge_inst),
    .io_core_exe_0_req_bits_fflags_bits_uop_pc_lob(lsu_io_core_exe_0_req_bits_fflags_bits_uop_pc_lob),
    .io_core_exe_0_req_bits_fflags_bits_uop_taken(lsu_io_core_exe_0_req_bits_fflags_bits_uop_taken),
    .io_core_exe_0_req_bits_fflags_bits_uop_imm_packed(lsu_io_core_exe_0_req_bits_fflags_bits_uop_imm_packed),
    .io_core_exe_0_req_bits_fflags_bits_uop_csr_addr(lsu_io_core_exe_0_req_bits_fflags_bits_uop_csr_addr),
    .io_core_exe_0_req_bits_fflags_bits_uop_rob_idx(lsu_io_core_exe_0_req_bits_fflags_bits_uop_rob_idx),
    .io_core_exe_0_req_bits_fflags_bits_uop_ldq_idx(lsu_io_core_exe_0_req_bits_fflags_bits_uop_ldq_idx),
    .io_core_exe_0_req_bits_fflags_bits_uop_stq_idx(lsu_io_core_exe_0_req_bits_fflags_bits_uop_stq_idx),
    .io_core_exe_0_req_bits_fflags_bits_uop_rxq_idx(lsu_io_core_exe_0_req_bits_fflags_bits_uop_rxq_idx),
    .io_core_exe_0_req_bits_fflags_bits_uop_pdst(lsu_io_core_exe_0_req_bits_fflags_bits_uop_pdst),
    .io_core_exe_0_req_bits_fflags_bits_uop_prs1(lsu_io_core_exe_0_req_bits_fflags_bits_uop_prs1),
    .io_core_exe_0_req_bits_fflags_bits_uop_prs2(lsu_io_core_exe_0_req_bits_fflags_bits_uop_prs2),
    .io_core_exe_0_req_bits_fflags_bits_uop_prs3(lsu_io_core_exe_0_req_bits_fflags_bits_uop_prs3),
    .io_core_exe_0_req_bits_fflags_bits_uop_ppred(lsu_io_core_exe_0_req_bits_fflags_bits_uop_ppred),
    .io_core_exe_0_req_bits_fflags_bits_uop_prs1_busy(lsu_io_core_exe_0_req_bits_fflags_bits_uop_prs1_busy),
    .io_core_exe_0_req_bits_fflags_bits_uop_prs2_busy(lsu_io_core_exe_0_req_bits_fflags_bits_uop_prs2_busy),
    .io_core_exe_0_req_bits_fflags_bits_uop_prs3_busy(lsu_io_core_exe_0_req_bits_fflags_bits_uop_prs3_busy),
    .io_core_exe_0_req_bits_fflags_bits_uop_ppred_busy(lsu_io_core_exe_0_req_bits_fflags_bits_uop_ppred_busy),
    .io_core_exe_0_req_bits_fflags_bits_uop_stale_pdst(lsu_io_core_exe_0_req_bits_fflags_bits_uop_stale_pdst),
    .io_core_exe_0_req_bits_fflags_bits_uop_exception(lsu_io_core_exe_0_req_bits_fflags_bits_uop_exception),
    .io_core_exe_0_req_bits_fflags_bits_uop_exc_cause(lsu_io_core_exe_0_req_bits_fflags_bits_uop_exc_cause),
    .io_core_exe_0_req_bits_fflags_bits_uop_bypassable(lsu_io_core_exe_0_req_bits_fflags_bits_uop_bypassable),
    .io_core_exe_0_req_bits_fflags_bits_uop_mem_cmd(lsu_io_core_exe_0_req_bits_fflags_bits_uop_mem_cmd),
    .io_core_exe_0_req_bits_fflags_bits_uop_mem_size(lsu_io_core_exe_0_req_bits_fflags_bits_uop_mem_size),
    .io_core_exe_0_req_bits_fflags_bits_uop_mem_signed(lsu_io_core_exe_0_req_bits_fflags_bits_uop_mem_signed),
    .io_core_exe_0_req_bits_fflags_bits_uop_is_fence(lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_fence),
    .io_core_exe_0_req_bits_fflags_bits_uop_is_fencei(lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_fencei),
    .io_core_exe_0_req_bits_fflags_bits_uop_is_amo(lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_amo),
    .io_core_exe_0_req_bits_fflags_bits_uop_uses_ldq(lsu_io_core_exe_0_req_bits_fflags_bits_uop_uses_ldq),
    .io_core_exe_0_req_bits_fflags_bits_uop_uses_stq(lsu_io_core_exe_0_req_bits_fflags_bits_uop_uses_stq),
    .io_core_exe_0_req_bits_fflags_bits_uop_is_sys_pc2epc(lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_sys_pc2epc),
    .io_core_exe_0_req_bits_fflags_bits_uop_is_unique(lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_unique),
    .io_core_exe_0_req_bits_fflags_bits_uop_flush_on_commit(lsu_io_core_exe_0_req_bits_fflags_bits_uop_flush_on_commit),
    .io_core_exe_0_req_bits_fflags_bits_uop_ldst_is_rs1(lsu_io_core_exe_0_req_bits_fflags_bits_uop_ldst_is_rs1),
    .io_core_exe_0_req_bits_fflags_bits_uop_ldst(lsu_io_core_exe_0_req_bits_fflags_bits_uop_ldst),
    .io_core_exe_0_req_bits_fflags_bits_uop_lrs1(lsu_io_core_exe_0_req_bits_fflags_bits_uop_lrs1),
    .io_core_exe_0_req_bits_fflags_bits_uop_lrs2(lsu_io_core_exe_0_req_bits_fflags_bits_uop_lrs2),
    .io_core_exe_0_req_bits_fflags_bits_uop_lrs3(lsu_io_core_exe_0_req_bits_fflags_bits_uop_lrs3),
    .io_core_exe_0_req_bits_fflags_bits_uop_ldst_val(lsu_io_core_exe_0_req_bits_fflags_bits_uop_ldst_val),
    .io_core_exe_0_req_bits_fflags_bits_uop_dst_rtype(lsu_io_core_exe_0_req_bits_fflags_bits_uop_dst_rtype),
    .io_core_exe_0_req_bits_fflags_bits_uop_lrs1_rtype(lsu_io_core_exe_0_req_bits_fflags_bits_uop_lrs1_rtype),
    .io_core_exe_0_req_bits_fflags_bits_uop_lrs2_rtype(lsu_io_core_exe_0_req_bits_fflags_bits_uop_lrs2_rtype),
    .io_core_exe_0_req_bits_fflags_bits_uop_frs3_en(lsu_io_core_exe_0_req_bits_fflags_bits_uop_frs3_en),
    .io_core_exe_0_req_bits_fflags_bits_uop_fp_val(lsu_io_core_exe_0_req_bits_fflags_bits_uop_fp_val),
    .io_core_exe_0_req_bits_fflags_bits_uop_fp_single(lsu_io_core_exe_0_req_bits_fflags_bits_uop_fp_single),
    .io_core_exe_0_req_bits_fflags_bits_uop_xcpt_pf_if(lsu_io_core_exe_0_req_bits_fflags_bits_uop_xcpt_pf_if),
    .io_core_exe_0_req_bits_fflags_bits_uop_xcpt_ae_if(lsu_io_core_exe_0_req_bits_fflags_bits_uop_xcpt_ae_if),
    .io_core_exe_0_req_bits_fflags_bits_uop_xcpt_ma_if(lsu_io_core_exe_0_req_bits_fflags_bits_uop_xcpt_ma_if),
    .io_core_exe_0_req_bits_fflags_bits_uop_bp_debug_if(lsu_io_core_exe_0_req_bits_fflags_bits_uop_bp_debug_if),
    .io_core_exe_0_req_bits_fflags_bits_uop_bp_xcpt_if(lsu_io_core_exe_0_req_bits_fflags_bits_uop_bp_xcpt_if),
    .io_core_exe_0_req_bits_fflags_bits_uop_debug_fsrc(lsu_io_core_exe_0_req_bits_fflags_bits_uop_debug_fsrc),
    .io_core_exe_0_req_bits_fflags_bits_uop_debug_tsrc(lsu_io_core_exe_0_req_bits_fflags_bits_uop_debug_tsrc),
    .io_core_exe_0_req_bits_fflags_bits_flags(lsu_io_core_exe_0_req_bits_fflags_bits_flags),
    .io_core_exe_0_req_bits_addr(lsu_io_core_exe_0_req_bits_addr),
    .io_core_exe_0_req_bits_mxcpt_valid(lsu_io_core_exe_0_req_bits_mxcpt_valid),
    .io_core_exe_0_req_bits_mxcpt_bits(lsu_io_core_exe_0_req_bits_mxcpt_bits),
    .io_core_exe_0_req_bits_sfence_valid(lsu_io_core_exe_0_req_bits_sfence_valid),
    .io_core_exe_0_req_bits_sfence_bits_rs1(lsu_io_core_exe_0_req_bits_sfence_bits_rs1),
    .io_core_exe_0_req_bits_sfence_bits_rs2(lsu_io_core_exe_0_req_bits_sfence_bits_rs2),
    .io_core_exe_0_req_bits_sfence_bits_addr(lsu_io_core_exe_0_req_bits_sfence_bits_addr),
    .io_core_exe_0_req_bits_sfence_bits_asid(lsu_io_core_exe_0_req_bits_sfence_bits_asid),
    .io_core_exe_0_req_bits_flagdata(lsu_io_core_exe_0_req_bits_flagdata),
    .io_core_exe_0_req_bits_fflagdata_valid(lsu_io_core_exe_0_req_bits_fflagdata_valid),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_switch(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_switch),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_switch_off(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_switch_off),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_is_unicore(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_unicore),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_shift(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_shift),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_lrs3_rtype(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_lrs3_rtype),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_rflag(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_rflag),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_wflag(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_wflag),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_prflag(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_prflag),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_pwflag(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_pwflag),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_pflag_busy(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_pflag_busy),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_stale_pflag(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_stale_pflag),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_op1_sel(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_op1_sel),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_op2_sel(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_op2_sel),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_split_num(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_split_num),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_self_index(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_self_index),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_rob_inst_idx(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_rob_inst_idx),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_address_num(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_address_num),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_uopc(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_uopc),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_inst(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_inst),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_debug_inst(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_debug_inst),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_is_rvc(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_rvc),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_debug_pc(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_debug_pc),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_iq_type(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_iq_type),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_fu_code(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_fu_code),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_br_type(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_br_type),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_op1_sel(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_op1_sel),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_op2_sel(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_op2_sel),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_imm_sel(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_imm_sel),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_op_fcn(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_op_fcn),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_fcn_dw(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_fcn_dw),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_csr_cmd(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_csr_cmd),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_load(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_load),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_sta(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_sta),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_std(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_std),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_op3_sel(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_op3_sel),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_iw_state(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_iw_state),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_iw_p1_poisoned(
      lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_iw_p1_poisoned),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_iw_p2_poisoned(
      lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_iw_p2_poisoned),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_is_br(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_br),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_is_jalr(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_jalr),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_is_jal(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_jal),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_is_sfb(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_sfb),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_br_mask(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_br_mask),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_br_tag(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_br_tag),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_ftq_idx(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ftq_idx),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_edge_inst(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_edge_inst),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_pc_lob(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_pc_lob),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_taken(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_taken),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_imm_packed(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_imm_packed),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_csr_addr(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_csr_addr),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_rob_idx(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_rob_idx),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_ldq_idx(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ldq_idx),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_stq_idx(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_stq_idx),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_rxq_idx(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_rxq_idx),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_pdst(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_pdst),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_prs1(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_prs1),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_prs2(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_prs2),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_prs3(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_prs3),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_ppred(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ppred),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_prs1_busy(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_prs1_busy),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_prs2_busy(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_prs2_busy),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_prs3_busy(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_prs3_busy),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_ppred_busy(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ppred_busy),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_stale_pdst(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_stale_pdst),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_exception(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_exception),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_exc_cause(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_exc_cause),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_bypassable(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_bypassable),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_mem_cmd(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_mem_cmd),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_mem_size(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_mem_size),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_mem_signed(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_mem_signed),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_is_fence(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_fence),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_is_fencei(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_fencei),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_is_amo(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_amo),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_uses_ldq(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_uses_ldq),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_uses_stq(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_uses_stq),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_is_sys_pc2epc(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_sys_pc2epc
      ),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_is_unique(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_unique),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_flush_on_commit(
      lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_flush_on_commit),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_ldst_is_rs1(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ldst_is_rs1),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_ldst(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ldst),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_lrs1(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_lrs1),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_lrs2(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_lrs2),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_lrs3(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_lrs3),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_ldst_val(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ldst_val),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_dst_rtype(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_dst_rtype),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_lrs1_rtype(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_lrs1_rtype),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_lrs2_rtype(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_lrs2_rtype),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_frs3_en(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_frs3_en),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_fp_val(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_fp_val),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_fp_single(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_fp_single),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_xcpt_pf_if(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_xcpt_pf_if),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_xcpt_ae_if(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_xcpt_ae_if),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_xcpt_ma_if(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_xcpt_ma_if),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_bp_debug_if(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_bp_debug_if),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_bp_xcpt_if(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_bp_xcpt_if),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_debug_fsrc(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_debug_fsrc),
    .io_core_exe_0_req_bits_fflagdata_bits_uop_debug_tsrc(lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_debug_tsrc),
    .io_core_exe_0_req_bits_fflagdata_bits_fflag(lsu_io_core_exe_0_req_bits_fflagdata_bits_fflag),
    .io_core_exe_0_iresp_ready(lsu_io_core_exe_0_iresp_ready),
    .io_core_exe_0_iresp_valid(lsu_io_core_exe_0_iresp_valid),
    .io_core_exe_0_iresp_bits_uop_switch(lsu_io_core_exe_0_iresp_bits_uop_switch),
    .io_core_exe_0_iresp_bits_uop_switch_off(lsu_io_core_exe_0_iresp_bits_uop_switch_off),
    .io_core_exe_0_iresp_bits_uop_is_unicore(lsu_io_core_exe_0_iresp_bits_uop_is_unicore),
    .io_core_exe_0_iresp_bits_uop_shift(lsu_io_core_exe_0_iresp_bits_uop_shift),
    .io_core_exe_0_iresp_bits_uop_lrs3_rtype(lsu_io_core_exe_0_iresp_bits_uop_lrs3_rtype),
    .io_core_exe_0_iresp_bits_uop_rflag(lsu_io_core_exe_0_iresp_bits_uop_rflag),
    .io_core_exe_0_iresp_bits_uop_wflag(lsu_io_core_exe_0_iresp_bits_uop_wflag),
    .io_core_exe_0_iresp_bits_uop_prflag(lsu_io_core_exe_0_iresp_bits_uop_prflag),
    .io_core_exe_0_iresp_bits_uop_pwflag(lsu_io_core_exe_0_iresp_bits_uop_pwflag),
    .io_core_exe_0_iresp_bits_uop_pflag_busy(lsu_io_core_exe_0_iresp_bits_uop_pflag_busy),
    .io_core_exe_0_iresp_bits_uop_stale_pflag(lsu_io_core_exe_0_iresp_bits_uop_stale_pflag),
    .io_core_exe_0_iresp_bits_uop_op1_sel(lsu_io_core_exe_0_iresp_bits_uop_op1_sel),
    .io_core_exe_0_iresp_bits_uop_op2_sel(lsu_io_core_exe_0_iresp_bits_uop_op2_sel),
    .io_core_exe_0_iresp_bits_uop_split_num(lsu_io_core_exe_0_iresp_bits_uop_split_num),
    .io_core_exe_0_iresp_bits_uop_self_index(lsu_io_core_exe_0_iresp_bits_uop_self_index),
    .io_core_exe_0_iresp_bits_uop_rob_inst_idx(lsu_io_core_exe_0_iresp_bits_uop_rob_inst_idx),
    .io_core_exe_0_iresp_bits_uop_address_num(lsu_io_core_exe_0_iresp_bits_uop_address_num),
    .io_core_exe_0_iresp_bits_uop_uopc(lsu_io_core_exe_0_iresp_bits_uop_uopc),
    .io_core_exe_0_iresp_bits_uop_inst(lsu_io_core_exe_0_iresp_bits_uop_inst),
    .io_core_exe_0_iresp_bits_uop_debug_inst(lsu_io_core_exe_0_iresp_bits_uop_debug_inst),
    .io_core_exe_0_iresp_bits_uop_is_rvc(lsu_io_core_exe_0_iresp_bits_uop_is_rvc),
    .io_core_exe_0_iresp_bits_uop_debug_pc(lsu_io_core_exe_0_iresp_bits_uop_debug_pc),
    .io_core_exe_0_iresp_bits_uop_iq_type(lsu_io_core_exe_0_iresp_bits_uop_iq_type),
    .io_core_exe_0_iresp_bits_uop_fu_code(lsu_io_core_exe_0_iresp_bits_uop_fu_code),
    .io_core_exe_0_iresp_bits_uop_ctrl_br_type(lsu_io_core_exe_0_iresp_bits_uop_ctrl_br_type),
    .io_core_exe_0_iresp_bits_uop_ctrl_op1_sel(lsu_io_core_exe_0_iresp_bits_uop_ctrl_op1_sel),
    .io_core_exe_0_iresp_bits_uop_ctrl_op2_sel(lsu_io_core_exe_0_iresp_bits_uop_ctrl_op2_sel),
    .io_core_exe_0_iresp_bits_uop_ctrl_imm_sel(lsu_io_core_exe_0_iresp_bits_uop_ctrl_imm_sel),
    .io_core_exe_0_iresp_bits_uop_ctrl_op_fcn(lsu_io_core_exe_0_iresp_bits_uop_ctrl_op_fcn),
    .io_core_exe_0_iresp_bits_uop_ctrl_fcn_dw(lsu_io_core_exe_0_iresp_bits_uop_ctrl_fcn_dw),
    .io_core_exe_0_iresp_bits_uop_ctrl_csr_cmd(lsu_io_core_exe_0_iresp_bits_uop_ctrl_csr_cmd),
    .io_core_exe_0_iresp_bits_uop_ctrl_is_load(lsu_io_core_exe_0_iresp_bits_uop_ctrl_is_load),
    .io_core_exe_0_iresp_bits_uop_ctrl_is_sta(lsu_io_core_exe_0_iresp_bits_uop_ctrl_is_sta),
    .io_core_exe_0_iresp_bits_uop_ctrl_is_std(lsu_io_core_exe_0_iresp_bits_uop_ctrl_is_std),
    .io_core_exe_0_iresp_bits_uop_ctrl_op3_sel(lsu_io_core_exe_0_iresp_bits_uop_ctrl_op3_sel),
    .io_core_exe_0_iresp_bits_uop_iw_state(lsu_io_core_exe_0_iresp_bits_uop_iw_state),
    .io_core_exe_0_iresp_bits_uop_iw_p1_poisoned(lsu_io_core_exe_0_iresp_bits_uop_iw_p1_poisoned),
    .io_core_exe_0_iresp_bits_uop_iw_p2_poisoned(lsu_io_core_exe_0_iresp_bits_uop_iw_p2_poisoned),
    .io_core_exe_0_iresp_bits_uop_is_br(lsu_io_core_exe_0_iresp_bits_uop_is_br),
    .io_core_exe_0_iresp_bits_uop_is_jalr(lsu_io_core_exe_0_iresp_bits_uop_is_jalr),
    .io_core_exe_0_iresp_bits_uop_is_jal(lsu_io_core_exe_0_iresp_bits_uop_is_jal),
    .io_core_exe_0_iresp_bits_uop_is_sfb(lsu_io_core_exe_0_iresp_bits_uop_is_sfb),
    .io_core_exe_0_iresp_bits_uop_br_mask(lsu_io_core_exe_0_iresp_bits_uop_br_mask),
    .io_core_exe_0_iresp_bits_uop_br_tag(lsu_io_core_exe_0_iresp_bits_uop_br_tag),
    .io_core_exe_0_iresp_bits_uop_ftq_idx(lsu_io_core_exe_0_iresp_bits_uop_ftq_idx),
    .io_core_exe_0_iresp_bits_uop_edge_inst(lsu_io_core_exe_0_iresp_bits_uop_edge_inst),
    .io_core_exe_0_iresp_bits_uop_pc_lob(lsu_io_core_exe_0_iresp_bits_uop_pc_lob),
    .io_core_exe_0_iresp_bits_uop_taken(lsu_io_core_exe_0_iresp_bits_uop_taken),
    .io_core_exe_0_iresp_bits_uop_imm_packed(lsu_io_core_exe_0_iresp_bits_uop_imm_packed),
    .io_core_exe_0_iresp_bits_uop_csr_addr(lsu_io_core_exe_0_iresp_bits_uop_csr_addr),
    .io_core_exe_0_iresp_bits_uop_rob_idx(lsu_io_core_exe_0_iresp_bits_uop_rob_idx),
    .io_core_exe_0_iresp_bits_uop_ldq_idx(lsu_io_core_exe_0_iresp_bits_uop_ldq_idx),
    .io_core_exe_0_iresp_bits_uop_stq_idx(lsu_io_core_exe_0_iresp_bits_uop_stq_idx),
    .io_core_exe_0_iresp_bits_uop_rxq_idx(lsu_io_core_exe_0_iresp_bits_uop_rxq_idx),
    .io_core_exe_0_iresp_bits_uop_pdst(lsu_io_core_exe_0_iresp_bits_uop_pdst),
    .io_core_exe_0_iresp_bits_uop_prs1(lsu_io_core_exe_0_iresp_bits_uop_prs1),
    .io_core_exe_0_iresp_bits_uop_prs2(lsu_io_core_exe_0_iresp_bits_uop_prs2),
    .io_core_exe_0_iresp_bits_uop_prs3(lsu_io_core_exe_0_iresp_bits_uop_prs3),
    .io_core_exe_0_iresp_bits_uop_ppred(lsu_io_core_exe_0_iresp_bits_uop_ppred),
    .io_core_exe_0_iresp_bits_uop_prs1_busy(lsu_io_core_exe_0_iresp_bits_uop_prs1_busy),
    .io_core_exe_0_iresp_bits_uop_prs2_busy(lsu_io_core_exe_0_iresp_bits_uop_prs2_busy),
    .io_core_exe_0_iresp_bits_uop_prs3_busy(lsu_io_core_exe_0_iresp_bits_uop_prs3_busy),
    .io_core_exe_0_iresp_bits_uop_ppred_busy(lsu_io_core_exe_0_iresp_bits_uop_ppred_busy),
    .io_core_exe_0_iresp_bits_uop_stale_pdst(lsu_io_core_exe_0_iresp_bits_uop_stale_pdst),
    .io_core_exe_0_iresp_bits_uop_exception(lsu_io_core_exe_0_iresp_bits_uop_exception),
    .io_core_exe_0_iresp_bits_uop_exc_cause(lsu_io_core_exe_0_iresp_bits_uop_exc_cause),
    .io_core_exe_0_iresp_bits_uop_bypassable(lsu_io_core_exe_0_iresp_bits_uop_bypassable),
    .io_core_exe_0_iresp_bits_uop_mem_cmd(lsu_io_core_exe_0_iresp_bits_uop_mem_cmd),
    .io_core_exe_0_iresp_bits_uop_mem_size(lsu_io_core_exe_0_iresp_bits_uop_mem_size),
    .io_core_exe_0_iresp_bits_uop_mem_signed(lsu_io_core_exe_0_iresp_bits_uop_mem_signed),
    .io_core_exe_0_iresp_bits_uop_is_fence(lsu_io_core_exe_0_iresp_bits_uop_is_fence),
    .io_core_exe_0_iresp_bits_uop_is_fencei(lsu_io_core_exe_0_iresp_bits_uop_is_fencei),
    .io_core_exe_0_iresp_bits_uop_is_amo(lsu_io_core_exe_0_iresp_bits_uop_is_amo),
    .io_core_exe_0_iresp_bits_uop_uses_ldq(lsu_io_core_exe_0_iresp_bits_uop_uses_ldq),
    .io_core_exe_0_iresp_bits_uop_uses_stq(lsu_io_core_exe_0_iresp_bits_uop_uses_stq),
    .io_core_exe_0_iresp_bits_uop_is_sys_pc2epc(lsu_io_core_exe_0_iresp_bits_uop_is_sys_pc2epc),
    .io_core_exe_0_iresp_bits_uop_is_unique(lsu_io_core_exe_0_iresp_bits_uop_is_unique),
    .io_core_exe_0_iresp_bits_uop_flush_on_commit(lsu_io_core_exe_0_iresp_bits_uop_flush_on_commit),
    .io_core_exe_0_iresp_bits_uop_ldst_is_rs1(lsu_io_core_exe_0_iresp_bits_uop_ldst_is_rs1),
    .io_core_exe_0_iresp_bits_uop_ldst(lsu_io_core_exe_0_iresp_bits_uop_ldst),
    .io_core_exe_0_iresp_bits_uop_lrs1(lsu_io_core_exe_0_iresp_bits_uop_lrs1),
    .io_core_exe_0_iresp_bits_uop_lrs2(lsu_io_core_exe_0_iresp_bits_uop_lrs2),
    .io_core_exe_0_iresp_bits_uop_lrs3(lsu_io_core_exe_0_iresp_bits_uop_lrs3),
    .io_core_exe_0_iresp_bits_uop_ldst_val(lsu_io_core_exe_0_iresp_bits_uop_ldst_val),
    .io_core_exe_0_iresp_bits_uop_dst_rtype(lsu_io_core_exe_0_iresp_bits_uop_dst_rtype),
    .io_core_exe_0_iresp_bits_uop_lrs1_rtype(lsu_io_core_exe_0_iresp_bits_uop_lrs1_rtype),
    .io_core_exe_0_iresp_bits_uop_lrs2_rtype(lsu_io_core_exe_0_iresp_bits_uop_lrs2_rtype),
    .io_core_exe_0_iresp_bits_uop_frs3_en(lsu_io_core_exe_0_iresp_bits_uop_frs3_en),
    .io_core_exe_0_iresp_bits_uop_fp_val(lsu_io_core_exe_0_iresp_bits_uop_fp_val),
    .io_core_exe_0_iresp_bits_uop_fp_single(lsu_io_core_exe_0_iresp_bits_uop_fp_single),
    .io_core_exe_0_iresp_bits_uop_xcpt_pf_if(lsu_io_core_exe_0_iresp_bits_uop_xcpt_pf_if),
    .io_core_exe_0_iresp_bits_uop_xcpt_ae_if(lsu_io_core_exe_0_iresp_bits_uop_xcpt_ae_if),
    .io_core_exe_0_iresp_bits_uop_xcpt_ma_if(lsu_io_core_exe_0_iresp_bits_uop_xcpt_ma_if),
    .io_core_exe_0_iresp_bits_uop_bp_debug_if(lsu_io_core_exe_0_iresp_bits_uop_bp_debug_if),
    .io_core_exe_0_iresp_bits_uop_bp_xcpt_if(lsu_io_core_exe_0_iresp_bits_uop_bp_xcpt_if),
    .io_core_exe_0_iresp_bits_uop_debug_fsrc(lsu_io_core_exe_0_iresp_bits_uop_debug_fsrc),
    .io_core_exe_0_iresp_bits_uop_debug_tsrc(lsu_io_core_exe_0_iresp_bits_uop_debug_tsrc),
    .io_core_exe_0_iresp_bits_data(lsu_io_core_exe_0_iresp_bits_data),
    .io_core_exe_0_iresp_bits_predicated(lsu_io_core_exe_0_iresp_bits_predicated),
    .io_core_exe_0_iresp_bits_fflags_valid(lsu_io_core_exe_0_iresp_bits_fflags_valid),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_switch(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_switch),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_switch_off(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_switch_off),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_is_unicore(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_unicore),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_shift(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_shift),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_lrs3_rtype(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_lrs3_rtype),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_rflag(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_rflag),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_wflag(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_wflag),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_prflag(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_prflag),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_pwflag(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_pwflag),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_pflag_busy(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_pflag_busy),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_stale_pflag(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_stale_pflag),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_op1_sel(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_op1_sel),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_op2_sel(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_op2_sel),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_split_num(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_split_num),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_self_index(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_self_index),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_rob_inst_idx(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_rob_inst_idx),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_address_num(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_address_num),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_uopc(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_uopc),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_inst(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_inst),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_debug_inst(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_debug_inst),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_is_rvc(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_rvc),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_debug_pc(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_debug_pc),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_iq_type(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_iq_type),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_fu_code(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_fu_code),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_br_type(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_br_type),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_op1_sel(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_op1_sel),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_op2_sel(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_op2_sel),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_imm_sel(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_imm_sel),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_op_fcn(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_op_fcn),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_fcn_dw(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_fcn_dw),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_csr_cmd(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_csr_cmd),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_load(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_load),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_sta(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_sta),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_std(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_std),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_op3_sel(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_op3_sel),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_iw_state(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_iw_state),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_iw_p1_poisoned(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_iw_p1_poisoned
      ),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_iw_p2_poisoned(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_iw_p2_poisoned
      ),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_is_br(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_br),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_is_jalr(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_jalr),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_is_jal(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_jal),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_is_sfb(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_sfb),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_br_mask(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_br_mask),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_br_tag(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_br_tag),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_ftq_idx(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ftq_idx),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_edge_inst(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_edge_inst),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_pc_lob(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_pc_lob),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_taken(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_taken),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_imm_packed(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_imm_packed),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_csr_addr(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_csr_addr),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_rob_idx(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_rob_idx),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_ldq_idx(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ldq_idx),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_stq_idx(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_stq_idx),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_rxq_idx(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_rxq_idx),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_pdst(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_pdst),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_prs1(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_prs1),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_prs2(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_prs2),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_prs3(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_prs3),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_ppred(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ppred),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_prs1_busy(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_prs1_busy),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_prs2_busy(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_prs2_busy),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_prs3_busy(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_prs3_busy),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_ppred_busy(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ppred_busy),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_stale_pdst(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_stale_pdst),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_exception(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_exception),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_exc_cause(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_exc_cause),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_bypassable(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_bypassable),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_mem_cmd(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_mem_cmd),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_mem_size(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_mem_size),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_mem_signed(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_mem_signed),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_is_fence(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_fence),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_is_fencei(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_fencei),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_is_amo(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_amo),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_uses_ldq(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_uses_ldq),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_uses_stq(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_uses_stq),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_is_sys_pc2epc(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_sys_pc2epc),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_is_unique(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_unique),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_flush_on_commit(
      lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_flush_on_commit),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_ldst_is_rs1(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ldst_is_rs1),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_ldst(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ldst),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_lrs1(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_lrs1),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_lrs2(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_lrs2),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_lrs3(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_lrs3),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_ldst_val(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ldst_val),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_dst_rtype(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_dst_rtype),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_lrs1_rtype(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_lrs1_rtype),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_lrs2_rtype(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_lrs2_rtype),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_frs3_en(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_frs3_en),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_fp_val(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_fp_val),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_fp_single(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_fp_single),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_xcpt_pf_if(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_xcpt_pf_if),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_xcpt_ae_if(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_xcpt_ae_if),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_xcpt_ma_if(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_xcpt_ma_if),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_bp_debug_if(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_bp_debug_if),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_bp_xcpt_if(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_bp_xcpt_if),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_debug_fsrc(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_debug_fsrc),
    .io_core_exe_0_iresp_bits_fflags_bits_uop_debug_tsrc(lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_debug_tsrc),
    .io_core_exe_0_iresp_bits_fflags_bits_flags(lsu_io_core_exe_0_iresp_bits_fflags_bits_flags),
    .io_core_exe_0_iresp_bits_flagdata(lsu_io_core_exe_0_iresp_bits_flagdata),
    .io_core_exe_0_iresp_bits_fflagdata_valid(lsu_io_core_exe_0_iresp_bits_fflagdata_valid),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_switch(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_switch),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_switch_off(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_switch_off),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_unicore(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_unicore),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_shift(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_shift),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs3_rtype(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs3_rtype),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_rflag(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_rflag),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_wflag(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_wflag),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_prflag(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_prflag),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_pwflag(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_pwflag),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_pflag_busy(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_pflag_busy),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_stale_pflag(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_stale_pflag
      ),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_op1_sel(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_op1_sel),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_op2_sel(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_op2_sel),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_split_num(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_split_num),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_self_index(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_self_index),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_rob_inst_idx(
      lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_rob_inst_idx),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_address_num(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_address_num
      ),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_uopc(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_uopc),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_inst(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_inst),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_debug_inst(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_debug_inst),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_rvc(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_rvc),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_debug_pc(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_debug_pc),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_iq_type(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_iq_type),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_fu_code(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_fu_code),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_br_type(
      lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_br_type),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op1_sel(
      lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op1_sel),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op2_sel(
      lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op2_sel),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_imm_sel(
      lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_imm_sel),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op_fcn(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op_fcn
      ),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_fcn_dw(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_fcn_dw
      ),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_csr_cmd(
      lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_csr_cmd),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_load(
      lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_load),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_sta(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_sta
      ),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_std(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_std
      ),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op3_sel(
      lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op3_sel),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_iw_state(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_iw_state),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_iw_p1_poisoned(
      lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_iw_p1_poisoned),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_iw_p2_poisoned(
      lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_iw_p2_poisoned),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_br(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_br),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_jalr(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_jalr),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_jal(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_jal),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_sfb(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_sfb),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_br_mask(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_br_mask),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_br_tag(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_br_tag),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_ftq_idx(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ftq_idx),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_edge_inst(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_edge_inst),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_pc_lob(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_pc_lob),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_taken(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_taken),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_imm_packed(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_imm_packed),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_csr_addr(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_csr_addr),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_rob_idx(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_rob_idx),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_ldq_idx(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ldq_idx),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_stq_idx(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_stq_idx),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_rxq_idx(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_rxq_idx),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_pdst(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_pdst),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs1(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs1),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs2(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs2),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs3(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs3),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_ppred(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ppred),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs1_busy(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs1_busy),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs2_busy(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs2_busy),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs3_busy(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs3_busy),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_ppred_busy(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ppred_busy),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_stale_pdst(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_stale_pdst),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_exception(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_exception),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_exc_cause(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_exc_cause),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_bypassable(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_bypassable),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_mem_cmd(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_mem_cmd),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_mem_size(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_mem_size),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_mem_signed(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_mem_signed),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_fence(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_fence),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_fencei(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_fencei),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_amo(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_amo),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_uses_ldq(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_uses_ldq),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_uses_stq(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_uses_stq),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_sys_pc2epc(
      lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_sys_pc2epc),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_unique(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_unique),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_flush_on_commit(
      lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_flush_on_commit),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_ldst_is_rs1(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ldst_is_rs1
      ),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_ldst(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ldst),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs1(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs1),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs2(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs2),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs3(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs3),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_ldst_val(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ldst_val),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_dst_rtype(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_dst_rtype),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs1_rtype(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs1_rtype),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs2_rtype(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs2_rtype),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_frs3_en(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_frs3_en),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_fp_val(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_fp_val),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_fp_single(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_fp_single),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_pf_if(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_pf_if),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_ae_if(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_ae_if),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_ma_if(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_ma_if),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_bp_debug_if(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_bp_debug_if
      ),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_bp_xcpt_if(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_bp_xcpt_if),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_debug_fsrc(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_debug_fsrc),
    .io_core_exe_0_iresp_bits_fflagdata_bits_uop_debug_tsrc(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_debug_tsrc),
    .io_core_exe_0_iresp_bits_fflagdata_bits_fflag(lsu_io_core_exe_0_iresp_bits_fflagdata_bits_fflag),
    .io_core_exe_0_fresp_ready(lsu_io_core_exe_0_fresp_ready),
    .io_core_exe_0_fresp_valid(lsu_io_core_exe_0_fresp_valid),
    .io_core_exe_0_fresp_bits_uop_switch(lsu_io_core_exe_0_fresp_bits_uop_switch),
    .io_core_exe_0_fresp_bits_uop_switch_off(lsu_io_core_exe_0_fresp_bits_uop_switch_off),
    .io_core_exe_0_fresp_bits_uop_is_unicore(lsu_io_core_exe_0_fresp_bits_uop_is_unicore),
    .io_core_exe_0_fresp_bits_uop_shift(lsu_io_core_exe_0_fresp_bits_uop_shift),
    .io_core_exe_0_fresp_bits_uop_lrs3_rtype(lsu_io_core_exe_0_fresp_bits_uop_lrs3_rtype),
    .io_core_exe_0_fresp_bits_uop_rflag(lsu_io_core_exe_0_fresp_bits_uop_rflag),
    .io_core_exe_0_fresp_bits_uop_wflag(lsu_io_core_exe_0_fresp_bits_uop_wflag),
    .io_core_exe_0_fresp_bits_uop_prflag(lsu_io_core_exe_0_fresp_bits_uop_prflag),
    .io_core_exe_0_fresp_bits_uop_pwflag(lsu_io_core_exe_0_fresp_bits_uop_pwflag),
    .io_core_exe_0_fresp_bits_uop_pflag_busy(lsu_io_core_exe_0_fresp_bits_uop_pflag_busy),
    .io_core_exe_0_fresp_bits_uop_stale_pflag(lsu_io_core_exe_0_fresp_bits_uop_stale_pflag),
    .io_core_exe_0_fresp_bits_uop_op1_sel(lsu_io_core_exe_0_fresp_bits_uop_op1_sel),
    .io_core_exe_0_fresp_bits_uop_op2_sel(lsu_io_core_exe_0_fresp_bits_uop_op2_sel),
    .io_core_exe_0_fresp_bits_uop_split_num(lsu_io_core_exe_0_fresp_bits_uop_split_num),
    .io_core_exe_0_fresp_bits_uop_self_index(lsu_io_core_exe_0_fresp_bits_uop_self_index),
    .io_core_exe_0_fresp_bits_uop_rob_inst_idx(lsu_io_core_exe_0_fresp_bits_uop_rob_inst_idx),
    .io_core_exe_0_fresp_bits_uop_address_num(lsu_io_core_exe_0_fresp_bits_uop_address_num),
    .io_core_exe_0_fresp_bits_uop_uopc(lsu_io_core_exe_0_fresp_bits_uop_uopc),
    .io_core_exe_0_fresp_bits_uop_inst(lsu_io_core_exe_0_fresp_bits_uop_inst),
    .io_core_exe_0_fresp_bits_uop_debug_inst(lsu_io_core_exe_0_fresp_bits_uop_debug_inst),
    .io_core_exe_0_fresp_bits_uop_is_rvc(lsu_io_core_exe_0_fresp_bits_uop_is_rvc),
    .io_core_exe_0_fresp_bits_uop_debug_pc(lsu_io_core_exe_0_fresp_bits_uop_debug_pc),
    .io_core_exe_0_fresp_bits_uop_iq_type(lsu_io_core_exe_0_fresp_bits_uop_iq_type),
    .io_core_exe_0_fresp_bits_uop_fu_code(lsu_io_core_exe_0_fresp_bits_uop_fu_code),
    .io_core_exe_0_fresp_bits_uop_ctrl_br_type(lsu_io_core_exe_0_fresp_bits_uop_ctrl_br_type),
    .io_core_exe_0_fresp_bits_uop_ctrl_op1_sel(lsu_io_core_exe_0_fresp_bits_uop_ctrl_op1_sel),
    .io_core_exe_0_fresp_bits_uop_ctrl_op2_sel(lsu_io_core_exe_0_fresp_bits_uop_ctrl_op2_sel),
    .io_core_exe_0_fresp_bits_uop_ctrl_imm_sel(lsu_io_core_exe_0_fresp_bits_uop_ctrl_imm_sel),
    .io_core_exe_0_fresp_bits_uop_ctrl_op_fcn(lsu_io_core_exe_0_fresp_bits_uop_ctrl_op_fcn),
    .io_core_exe_0_fresp_bits_uop_ctrl_fcn_dw(lsu_io_core_exe_0_fresp_bits_uop_ctrl_fcn_dw),
    .io_core_exe_0_fresp_bits_uop_ctrl_csr_cmd(lsu_io_core_exe_0_fresp_bits_uop_ctrl_csr_cmd),
    .io_core_exe_0_fresp_bits_uop_ctrl_is_load(lsu_io_core_exe_0_fresp_bits_uop_ctrl_is_load),
    .io_core_exe_0_fresp_bits_uop_ctrl_is_sta(lsu_io_core_exe_0_fresp_bits_uop_ctrl_is_sta),
    .io_core_exe_0_fresp_bits_uop_ctrl_is_std(lsu_io_core_exe_0_fresp_bits_uop_ctrl_is_std),
    .io_core_exe_0_fresp_bits_uop_ctrl_op3_sel(lsu_io_core_exe_0_fresp_bits_uop_ctrl_op3_sel),
    .io_core_exe_0_fresp_bits_uop_iw_state(lsu_io_core_exe_0_fresp_bits_uop_iw_state),
    .io_core_exe_0_fresp_bits_uop_iw_p1_poisoned(lsu_io_core_exe_0_fresp_bits_uop_iw_p1_poisoned),
    .io_core_exe_0_fresp_bits_uop_iw_p2_poisoned(lsu_io_core_exe_0_fresp_bits_uop_iw_p2_poisoned),
    .io_core_exe_0_fresp_bits_uop_is_br(lsu_io_core_exe_0_fresp_bits_uop_is_br),
    .io_core_exe_0_fresp_bits_uop_is_jalr(lsu_io_core_exe_0_fresp_bits_uop_is_jalr),
    .io_core_exe_0_fresp_bits_uop_is_jal(lsu_io_core_exe_0_fresp_bits_uop_is_jal),
    .io_core_exe_0_fresp_bits_uop_is_sfb(lsu_io_core_exe_0_fresp_bits_uop_is_sfb),
    .io_core_exe_0_fresp_bits_uop_br_mask(lsu_io_core_exe_0_fresp_bits_uop_br_mask),
    .io_core_exe_0_fresp_bits_uop_br_tag(lsu_io_core_exe_0_fresp_bits_uop_br_tag),
    .io_core_exe_0_fresp_bits_uop_ftq_idx(lsu_io_core_exe_0_fresp_bits_uop_ftq_idx),
    .io_core_exe_0_fresp_bits_uop_edge_inst(lsu_io_core_exe_0_fresp_bits_uop_edge_inst),
    .io_core_exe_0_fresp_bits_uop_pc_lob(lsu_io_core_exe_0_fresp_bits_uop_pc_lob),
    .io_core_exe_0_fresp_bits_uop_taken(lsu_io_core_exe_0_fresp_bits_uop_taken),
    .io_core_exe_0_fresp_bits_uop_imm_packed(lsu_io_core_exe_0_fresp_bits_uop_imm_packed),
    .io_core_exe_0_fresp_bits_uop_csr_addr(lsu_io_core_exe_0_fresp_bits_uop_csr_addr),
    .io_core_exe_0_fresp_bits_uop_rob_idx(lsu_io_core_exe_0_fresp_bits_uop_rob_idx),
    .io_core_exe_0_fresp_bits_uop_ldq_idx(lsu_io_core_exe_0_fresp_bits_uop_ldq_idx),
    .io_core_exe_0_fresp_bits_uop_stq_idx(lsu_io_core_exe_0_fresp_bits_uop_stq_idx),
    .io_core_exe_0_fresp_bits_uop_rxq_idx(lsu_io_core_exe_0_fresp_bits_uop_rxq_idx),
    .io_core_exe_0_fresp_bits_uop_pdst(lsu_io_core_exe_0_fresp_bits_uop_pdst),
    .io_core_exe_0_fresp_bits_uop_prs1(lsu_io_core_exe_0_fresp_bits_uop_prs1),
    .io_core_exe_0_fresp_bits_uop_prs2(lsu_io_core_exe_0_fresp_bits_uop_prs2),
    .io_core_exe_0_fresp_bits_uop_prs3(lsu_io_core_exe_0_fresp_bits_uop_prs3),
    .io_core_exe_0_fresp_bits_uop_ppred(lsu_io_core_exe_0_fresp_bits_uop_ppred),
    .io_core_exe_0_fresp_bits_uop_prs1_busy(lsu_io_core_exe_0_fresp_bits_uop_prs1_busy),
    .io_core_exe_0_fresp_bits_uop_prs2_busy(lsu_io_core_exe_0_fresp_bits_uop_prs2_busy),
    .io_core_exe_0_fresp_bits_uop_prs3_busy(lsu_io_core_exe_0_fresp_bits_uop_prs3_busy),
    .io_core_exe_0_fresp_bits_uop_ppred_busy(lsu_io_core_exe_0_fresp_bits_uop_ppred_busy),
    .io_core_exe_0_fresp_bits_uop_stale_pdst(lsu_io_core_exe_0_fresp_bits_uop_stale_pdst),
    .io_core_exe_0_fresp_bits_uop_exception(lsu_io_core_exe_0_fresp_bits_uop_exception),
    .io_core_exe_0_fresp_bits_uop_exc_cause(lsu_io_core_exe_0_fresp_bits_uop_exc_cause),
    .io_core_exe_0_fresp_bits_uop_bypassable(lsu_io_core_exe_0_fresp_bits_uop_bypassable),
    .io_core_exe_0_fresp_bits_uop_mem_cmd(lsu_io_core_exe_0_fresp_bits_uop_mem_cmd),
    .io_core_exe_0_fresp_bits_uop_mem_size(lsu_io_core_exe_0_fresp_bits_uop_mem_size),
    .io_core_exe_0_fresp_bits_uop_mem_signed(lsu_io_core_exe_0_fresp_bits_uop_mem_signed),
    .io_core_exe_0_fresp_bits_uop_is_fence(lsu_io_core_exe_0_fresp_bits_uop_is_fence),
    .io_core_exe_0_fresp_bits_uop_is_fencei(lsu_io_core_exe_0_fresp_bits_uop_is_fencei),
    .io_core_exe_0_fresp_bits_uop_is_amo(lsu_io_core_exe_0_fresp_bits_uop_is_amo),
    .io_core_exe_0_fresp_bits_uop_uses_ldq(lsu_io_core_exe_0_fresp_bits_uop_uses_ldq),
    .io_core_exe_0_fresp_bits_uop_uses_stq(lsu_io_core_exe_0_fresp_bits_uop_uses_stq),
    .io_core_exe_0_fresp_bits_uop_is_sys_pc2epc(lsu_io_core_exe_0_fresp_bits_uop_is_sys_pc2epc),
    .io_core_exe_0_fresp_bits_uop_is_unique(lsu_io_core_exe_0_fresp_bits_uop_is_unique),
    .io_core_exe_0_fresp_bits_uop_flush_on_commit(lsu_io_core_exe_0_fresp_bits_uop_flush_on_commit),
    .io_core_exe_0_fresp_bits_uop_ldst_is_rs1(lsu_io_core_exe_0_fresp_bits_uop_ldst_is_rs1),
    .io_core_exe_0_fresp_bits_uop_ldst(lsu_io_core_exe_0_fresp_bits_uop_ldst),
    .io_core_exe_0_fresp_bits_uop_lrs1(lsu_io_core_exe_0_fresp_bits_uop_lrs1),
    .io_core_exe_0_fresp_bits_uop_lrs2(lsu_io_core_exe_0_fresp_bits_uop_lrs2),
    .io_core_exe_0_fresp_bits_uop_lrs3(lsu_io_core_exe_0_fresp_bits_uop_lrs3),
    .io_core_exe_0_fresp_bits_uop_ldst_val(lsu_io_core_exe_0_fresp_bits_uop_ldst_val),
    .io_core_exe_0_fresp_bits_uop_dst_rtype(lsu_io_core_exe_0_fresp_bits_uop_dst_rtype),
    .io_core_exe_0_fresp_bits_uop_lrs1_rtype(lsu_io_core_exe_0_fresp_bits_uop_lrs1_rtype),
    .io_core_exe_0_fresp_bits_uop_lrs2_rtype(lsu_io_core_exe_0_fresp_bits_uop_lrs2_rtype),
    .io_core_exe_0_fresp_bits_uop_frs3_en(lsu_io_core_exe_0_fresp_bits_uop_frs3_en),
    .io_core_exe_0_fresp_bits_uop_fp_val(lsu_io_core_exe_0_fresp_bits_uop_fp_val),
    .io_core_exe_0_fresp_bits_uop_fp_single(lsu_io_core_exe_0_fresp_bits_uop_fp_single),
    .io_core_exe_0_fresp_bits_uop_xcpt_pf_if(lsu_io_core_exe_0_fresp_bits_uop_xcpt_pf_if),
    .io_core_exe_0_fresp_bits_uop_xcpt_ae_if(lsu_io_core_exe_0_fresp_bits_uop_xcpt_ae_if),
    .io_core_exe_0_fresp_bits_uop_xcpt_ma_if(lsu_io_core_exe_0_fresp_bits_uop_xcpt_ma_if),
    .io_core_exe_0_fresp_bits_uop_bp_debug_if(lsu_io_core_exe_0_fresp_bits_uop_bp_debug_if),
    .io_core_exe_0_fresp_bits_uop_bp_xcpt_if(lsu_io_core_exe_0_fresp_bits_uop_bp_xcpt_if),
    .io_core_exe_0_fresp_bits_uop_debug_fsrc(lsu_io_core_exe_0_fresp_bits_uop_debug_fsrc),
    .io_core_exe_0_fresp_bits_uop_debug_tsrc(lsu_io_core_exe_0_fresp_bits_uop_debug_tsrc),
    .io_core_exe_0_fresp_bits_data(lsu_io_core_exe_0_fresp_bits_data),
    .io_core_exe_0_fresp_bits_predicated(lsu_io_core_exe_0_fresp_bits_predicated),
    .io_core_exe_0_fresp_bits_fflags_valid(lsu_io_core_exe_0_fresp_bits_fflags_valid),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_switch(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_switch),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_switch_off(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_switch_off),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_is_unicore(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_unicore),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_shift(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_shift),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_lrs3_rtype(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_lrs3_rtype),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_rflag(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_rflag),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_wflag(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_wflag),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_prflag(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_prflag),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_pwflag(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_pwflag),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_pflag_busy(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_pflag_busy),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_stale_pflag(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_stale_pflag),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_op1_sel(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_op1_sel),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_op2_sel(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_op2_sel),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_split_num(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_split_num),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_self_index(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_self_index),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_rob_inst_idx(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_rob_inst_idx),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_address_num(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_address_num),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_uopc(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_uopc),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_inst(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_inst),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_debug_inst(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_debug_inst),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_is_rvc(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_rvc),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_debug_pc(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_debug_pc),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_iq_type(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_iq_type),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_fu_code(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_fu_code),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_br_type(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_br_type),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_op1_sel(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_op1_sel),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_op2_sel(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_op2_sel),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_imm_sel(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_imm_sel),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_op_fcn(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_op_fcn),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_fcn_dw(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_fcn_dw),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_csr_cmd(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_csr_cmd),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_load(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_load),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_sta(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_sta),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_std(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_std),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_op3_sel(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_op3_sel),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_iw_state(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_iw_state),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_iw_p1_poisoned(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_iw_p1_poisoned
      ),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_iw_p2_poisoned(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_iw_p2_poisoned
      ),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_is_br(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_br),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_is_jalr(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_jalr),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_is_jal(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_jal),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_is_sfb(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_sfb),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_br_mask(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_br_mask),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_br_tag(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_br_tag),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_ftq_idx(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ftq_idx),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_edge_inst(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_edge_inst),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_pc_lob(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_pc_lob),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_taken(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_taken),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_imm_packed(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_imm_packed),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_csr_addr(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_csr_addr),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_rob_idx(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_rob_idx),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_ldq_idx(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ldq_idx),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_stq_idx(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_stq_idx),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_rxq_idx(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_rxq_idx),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_pdst(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_pdst),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_prs1(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_prs1),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_prs2(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_prs2),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_prs3(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_prs3),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_ppred(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ppred),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_prs1_busy(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_prs1_busy),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_prs2_busy(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_prs2_busy),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_prs3_busy(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_prs3_busy),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_ppred_busy(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ppred_busy),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_stale_pdst(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_stale_pdst),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_exception(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_exception),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_exc_cause(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_exc_cause),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_bypassable(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_bypassable),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_mem_cmd(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_mem_cmd),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_mem_size(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_mem_size),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_mem_signed(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_mem_signed),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_is_fence(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_fence),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_is_fencei(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_fencei),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_is_amo(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_amo),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_uses_ldq(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_uses_ldq),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_uses_stq(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_uses_stq),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_is_sys_pc2epc(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_sys_pc2epc),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_is_unique(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_unique),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_flush_on_commit(
      lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_flush_on_commit),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_ldst_is_rs1(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ldst_is_rs1),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_ldst(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ldst),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_lrs1(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_lrs1),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_lrs2(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_lrs2),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_lrs3(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_lrs3),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_ldst_val(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ldst_val),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_dst_rtype(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_dst_rtype),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_lrs1_rtype(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_lrs1_rtype),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_lrs2_rtype(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_lrs2_rtype),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_frs3_en(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_frs3_en),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_fp_val(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_fp_val),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_fp_single(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_fp_single),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_xcpt_pf_if(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_xcpt_pf_if),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_xcpt_ae_if(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_xcpt_ae_if),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_xcpt_ma_if(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_xcpt_ma_if),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_bp_debug_if(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_bp_debug_if),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_bp_xcpt_if(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_bp_xcpt_if),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_debug_fsrc(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_debug_fsrc),
    .io_core_exe_0_fresp_bits_fflags_bits_uop_debug_tsrc(lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_debug_tsrc),
    .io_core_exe_0_fresp_bits_fflags_bits_flags(lsu_io_core_exe_0_fresp_bits_fflags_bits_flags),
    .io_core_exe_0_fresp_bits_flagdata(lsu_io_core_exe_0_fresp_bits_flagdata),
    .io_core_exe_0_fresp_bits_fflagdata_valid(lsu_io_core_exe_0_fresp_bits_fflagdata_valid),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_switch(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_switch),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_switch_off(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_switch_off),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_unicore(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_unicore),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_shift(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_shift),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs3_rtype(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs3_rtype),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_rflag(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_rflag),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_wflag(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_wflag),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_prflag(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_prflag),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_pwflag(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_pwflag),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_pflag_busy(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_pflag_busy),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_stale_pflag(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_stale_pflag
      ),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_op1_sel(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_op1_sel),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_op2_sel(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_op2_sel),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_split_num(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_split_num),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_self_index(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_self_index),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_rob_inst_idx(
      lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_rob_inst_idx),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_address_num(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_address_num
      ),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_uopc(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_uopc),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_inst(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_inst),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_debug_inst(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_debug_inst),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_rvc(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_rvc),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_debug_pc(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_debug_pc),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_iq_type(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_iq_type),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_fu_code(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_fu_code),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_br_type(
      lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_br_type),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op1_sel(
      lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op1_sel),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op2_sel(
      lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op2_sel),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_imm_sel(
      lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_imm_sel),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op_fcn(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op_fcn
      ),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_fcn_dw(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_fcn_dw
      ),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_csr_cmd(
      lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_csr_cmd),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_load(
      lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_load),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_sta(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_sta
      ),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_std(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_std
      ),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op3_sel(
      lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op3_sel),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_iw_state(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_iw_state),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_iw_p1_poisoned(
      lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_iw_p1_poisoned),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_iw_p2_poisoned(
      lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_iw_p2_poisoned),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_br(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_br),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_jalr(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_jalr),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_jal(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_jal),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_sfb(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_sfb),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_br_mask(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_br_mask),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_br_tag(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_br_tag),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_ftq_idx(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ftq_idx),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_edge_inst(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_edge_inst),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_pc_lob(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_pc_lob),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_taken(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_taken),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_imm_packed(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_imm_packed),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_csr_addr(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_csr_addr),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_rob_idx(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_rob_idx),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_ldq_idx(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ldq_idx),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_stq_idx(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_stq_idx),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_rxq_idx(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_rxq_idx),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_pdst(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_pdst),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs1(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs1),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs2(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs2),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs3(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs3),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_ppred(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ppred),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs1_busy(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs1_busy),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs2_busy(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs2_busy),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs3_busy(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs3_busy),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_ppred_busy(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ppred_busy),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_stale_pdst(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_stale_pdst),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_exception(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_exception),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_exc_cause(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_exc_cause),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_bypassable(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_bypassable),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_mem_cmd(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_mem_cmd),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_mem_size(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_mem_size),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_mem_signed(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_mem_signed),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_fence(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_fence),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_fencei(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_fencei),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_amo(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_amo),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_uses_ldq(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_uses_ldq),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_uses_stq(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_uses_stq),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_sys_pc2epc(
      lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_sys_pc2epc),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_unique(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_unique),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_flush_on_commit(
      lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_flush_on_commit),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_ldst_is_rs1(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ldst_is_rs1
      ),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_ldst(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ldst),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs1(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs1),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs2(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs2),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs3(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs3),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_ldst_val(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ldst_val),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_dst_rtype(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_dst_rtype),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs1_rtype(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs1_rtype),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs2_rtype(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs2_rtype),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_frs3_en(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_frs3_en),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_fp_val(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_fp_val),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_fp_single(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_fp_single),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_pf_if(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_pf_if),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_ae_if(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_ae_if),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_ma_if(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_ma_if),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_bp_debug_if(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_bp_debug_if
      ),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_bp_xcpt_if(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_bp_xcpt_if),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_debug_fsrc(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_debug_fsrc),
    .io_core_exe_0_fresp_bits_fflagdata_bits_uop_debug_tsrc(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_debug_tsrc),
    .io_core_exe_0_fresp_bits_fflagdata_bits_fflag(lsu_io_core_exe_0_fresp_bits_fflagdata_bits_fflag),
    .io_core_dis_uops_0_valid(lsu_io_core_dis_uops_0_valid),
    .io_core_dis_uops_0_bits_switch(lsu_io_core_dis_uops_0_bits_switch),
    .io_core_dis_uops_0_bits_switch_off(lsu_io_core_dis_uops_0_bits_switch_off),
    .io_core_dis_uops_0_bits_is_unicore(lsu_io_core_dis_uops_0_bits_is_unicore),
    .io_core_dis_uops_0_bits_shift(lsu_io_core_dis_uops_0_bits_shift),
    .io_core_dis_uops_0_bits_lrs3_rtype(lsu_io_core_dis_uops_0_bits_lrs3_rtype),
    .io_core_dis_uops_0_bits_rflag(lsu_io_core_dis_uops_0_bits_rflag),
    .io_core_dis_uops_0_bits_wflag(lsu_io_core_dis_uops_0_bits_wflag),
    .io_core_dis_uops_0_bits_prflag(lsu_io_core_dis_uops_0_bits_prflag),
    .io_core_dis_uops_0_bits_pwflag(lsu_io_core_dis_uops_0_bits_pwflag),
    .io_core_dis_uops_0_bits_pflag_busy(lsu_io_core_dis_uops_0_bits_pflag_busy),
    .io_core_dis_uops_0_bits_stale_pflag(lsu_io_core_dis_uops_0_bits_stale_pflag),
    .io_core_dis_uops_0_bits_op1_sel(lsu_io_core_dis_uops_0_bits_op1_sel),
    .io_core_dis_uops_0_bits_op2_sel(lsu_io_core_dis_uops_0_bits_op2_sel),
    .io_core_dis_uops_0_bits_split_num(lsu_io_core_dis_uops_0_bits_split_num),
    .io_core_dis_uops_0_bits_self_index(lsu_io_core_dis_uops_0_bits_self_index),
    .io_core_dis_uops_0_bits_rob_inst_idx(lsu_io_core_dis_uops_0_bits_rob_inst_idx),
    .io_core_dis_uops_0_bits_address_num(lsu_io_core_dis_uops_0_bits_address_num),
    .io_core_dis_uops_0_bits_uopc(lsu_io_core_dis_uops_0_bits_uopc),
    .io_core_dis_uops_0_bits_inst(lsu_io_core_dis_uops_0_bits_inst),
    .io_core_dis_uops_0_bits_debug_inst(lsu_io_core_dis_uops_0_bits_debug_inst),
    .io_core_dis_uops_0_bits_is_rvc(lsu_io_core_dis_uops_0_bits_is_rvc),
    .io_core_dis_uops_0_bits_debug_pc(lsu_io_core_dis_uops_0_bits_debug_pc),
    .io_core_dis_uops_0_bits_iq_type(lsu_io_core_dis_uops_0_bits_iq_type),
    .io_core_dis_uops_0_bits_fu_code(lsu_io_core_dis_uops_0_bits_fu_code),
    .io_core_dis_uops_0_bits_ctrl_br_type(lsu_io_core_dis_uops_0_bits_ctrl_br_type),
    .io_core_dis_uops_0_bits_ctrl_op1_sel(lsu_io_core_dis_uops_0_bits_ctrl_op1_sel),
    .io_core_dis_uops_0_bits_ctrl_op2_sel(lsu_io_core_dis_uops_0_bits_ctrl_op2_sel),
    .io_core_dis_uops_0_bits_ctrl_imm_sel(lsu_io_core_dis_uops_0_bits_ctrl_imm_sel),
    .io_core_dis_uops_0_bits_ctrl_op_fcn(lsu_io_core_dis_uops_0_bits_ctrl_op_fcn),
    .io_core_dis_uops_0_bits_ctrl_fcn_dw(lsu_io_core_dis_uops_0_bits_ctrl_fcn_dw),
    .io_core_dis_uops_0_bits_ctrl_csr_cmd(lsu_io_core_dis_uops_0_bits_ctrl_csr_cmd),
    .io_core_dis_uops_0_bits_ctrl_is_load(lsu_io_core_dis_uops_0_bits_ctrl_is_load),
    .io_core_dis_uops_0_bits_ctrl_is_sta(lsu_io_core_dis_uops_0_bits_ctrl_is_sta),
    .io_core_dis_uops_0_bits_ctrl_is_std(lsu_io_core_dis_uops_0_bits_ctrl_is_std),
    .io_core_dis_uops_0_bits_ctrl_op3_sel(lsu_io_core_dis_uops_0_bits_ctrl_op3_sel),
    .io_core_dis_uops_0_bits_iw_state(lsu_io_core_dis_uops_0_bits_iw_state),
    .io_core_dis_uops_0_bits_iw_p1_poisoned(lsu_io_core_dis_uops_0_bits_iw_p1_poisoned),
    .io_core_dis_uops_0_bits_iw_p2_poisoned(lsu_io_core_dis_uops_0_bits_iw_p2_poisoned),
    .io_core_dis_uops_0_bits_is_br(lsu_io_core_dis_uops_0_bits_is_br),
    .io_core_dis_uops_0_bits_is_jalr(lsu_io_core_dis_uops_0_bits_is_jalr),
    .io_core_dis_uops_0_bits_is_jal(lsu_io_core_dis_uops_0_bits_is_jal),
    .io_core_dis_uops_0_bits_is_sfb(lsu_io_core_dis_uops_0_bits_is_sfb),
    .io_core_dis_uops_0_bits_br_mask(lsu_io_core_dis_uops_0_bits_br_mask),
    .io_core_dis_uops_0_bits_br_tag(lsu_io_core_dis_uops_0_bits_br_tag),
    .io_core_dis_uops_0_bits_ftq_idx(lsu_io_core_dis_uops_0_bits_ftq_idx),
    .io_core_dis_uops_0_bits_edge_inst(lsu_io_core_dis_uops_0_bits_edge_inst),
    .io_core_dis_uops_0_bits_pc_lob(lsu_io_core_dis_uops_0_bits_pc_lob),
    .io_core_dis_uops_0_bits_taken(lsu_io_core_dis_uops_0_bits_taken),
    .io_core_dis_uops_0_bits_imm_packed(lsu_io_core_dis_uops_0_bits_imm_packed),
    .io_core_dis_uops_0_bits_csr_addr(lsu_io_core_dis_uops_0_bits_csr_addr),
    .io_core_dis_uops_0_bits_rob_idx(lsu_io_core_dis_uops_0_bits_rob_idx),
    .io_core_dis_uops_0_bits_ldq_idx(lsu_io_core_dis_uops_0_bits_ldq_idx),
    .io_core_dis_uops_0_bits_stq_idx(lsu_io_core_dis_uops_0_bits_stq_idx),
    .io_core_dis_uops_0_bits_rxq_idx(lsu_io_core_dis_uops_0_bits_rxq_idx),
    .io_core_dis_uops_0_bits_pdst(lsu_io_core_dis_uops_0_bits_pdst),
    .io_core_dis_uops_0_bits_prs1(lsu_io_core_dis_uops_0_bits_prs1),
    .io_core_dis_uops_0_bits_prs2(lsu_io_core_dis_uops_0_bits_prs2),
    .io_core_dis_uops_0_bits_prs3(lsu_io_core_dis_uops_0_bits_prs3),
    .io_core_dis_uops_0_bits_ppred(lsu_io_core_dis_uops_0_bits_ppred),
    .io_core_dis_uops_0_bits_prs1_busy(lsu_io_core_dis_uops_0_bits_prs1_busy),
    .io_core_dis_uops_0_bits_prs2_busy(lsu_io_core_dis_uops_0_bits_prs2_busy),
    .io_core_dis_uops_0_bits_prs3_busy(lsu_io_core_dis_uops_0_bits_prs3_busy),
    .io_core_dis_uops_0_bits_ppred_busy(lsu_io_core_dis_uops_0_bits_ppred_busy),
    .io_core_dis_uops_0_bits_stale_pdst(lsu_io_core_dis_uops_0_bits_stale_pdst),
    .io_core_dis_uops_0_bits_exception(lsu_io_core_dis_uops_0_bits_exception),
    .io_core_dis_uops_0_bits_exc_cause(lsu_io_core_dis_uops_0_bits_exc_cause),
    .io_core_dis_uops_0_bits_bypassable(lsu_io_core_dis_uops_0_bits_bypassable),
    .io_core_dis_uops_0_bits_mem_cmd(lsu_io_core_dis_uops_0_bits_mem_cmd),
    .io_core_dis_uops_0_bits_mem_size(lsu_io_core_dis_uops_0_bits_mem_size),
    .io_core_dis_uops_0_bits_mem_signed(lsu_io_core_dis_uops_0_bits_mem_signed),
    .io_core_dis_uops_0_bits_is_fence(lsu_io_core_dis_uops_0_bits_is_fence),
    .io_core_dis_uops_0_bits_is_fencei(lsu_io_core_dis_uops_0_bits_is_fencei),
    .io_core_dis_uops_0_bits_is_amo(lsu_io_core_dis_uops_0_bits_is_amo),
    .io_core_dis_uops_0_bits_uses_ldq(lsu_io_core_dis_uops_0_bits_uses_ldq),
    .io_core_dis_uops_0_bits_uses_stq(lsu_io_core_dis_uops_0_bits_uses_stq),
    .io_core_dis_uops_0_bits_is_sys_pc2epc(lsu_io_core_dis_uops_0_bits_is_sys_pc2epc),
    .io_core_dis_uops_0_bits_is_unique(lsu_io_core_dis_uops_0_bits_is_unique),
    .io_core_dis_uops_0_bits_flush_on_commit(lsu_io_core_dis_uops_0_bits_flush_on_commit),
    .io_core_dis_uops_0_bits_ldst_is_rs1(lsu_io_core_dis_uops_0_bits_ldst_is_rs1),
    .io_core_dis_uops_0_bits_ldst(lsu_io_core_dis_uops_0_bits_ldst),
    .io_core_dis_uops_0_bits_lrs1(lsu_io_core_dis_uops_0_bits_lrs1),
    .io_core_dis_uops_0_bits_lrs2(lsu_io_core_dis_uops_0_bits_lrs2),
    .io_core_dis_uops_0_bits_lrs3(lsu_io_core_dis_uops_0_bits_lrs3),
    .io_core_dis_uops_0_bits_ldst_val(lsu_io_core_dis_uops_0_bits_ldst_val),
    .io_core_dis_uops_0_bits_dst_rtype(lsu_io_core_dis_uops_0_bits_dst_rtype),
    .io_core_dis_uops_0_bits_lrs1_rtype(lsu_io_core_dis_uops_0_bits_lrs1_rtype),
    .io_core_dis_uops_0_bits_lrs2_rtype(lsu_io_core_dis_uops_0_bits_lrs2_rtype),
    .io_core_dis_uops_0_bits_frs3_en(lsu_io_core_dis_uops_0_bits_frs3_en),
    .io_core_dis_uops_0_bits_fp_val(lsu_io_core_dis_uops_0_bits_fp_val),
    .io_core_dis_uops_0_bits_fp_single(lsu_io_core_dis_uops_0_bits_fp_single),
    .io_core_dis_uops_0_bits_xcpt_pf_if(lsu_io_core_dis_uops_0_bits_xcpt_pf_if),
    .io_core_dis_uops_0_bits_xcpt_ae_if(lsu_io_core_dis_uops_0_bits_xcpt_ae_if),
    .io_core_dis_uops_0_bits_xcpt_ma_if(lsu_io_core_dis_uops_0_bits_xcpt_ma_if),
    .io_core_dis_uops_0_bits_bp_debug_if(lsu_io_core_dis_uops_0_bits_bp_debug_if),
    .io_core_dis_uops_0_bits_bp_xcpt_if(lsu_io_core_dis_uops_0_bits_bp_xcpt_if),
    .io_core_dis_uops_0_bits_debug_fsrc(lsu_io_core_dis_uops_0_bits_debug_fsrc),
    .io_core_dis_uops_0_bits_debug_tsrc(lsu_io_core_dis_uops_0_bits_debug_tsrc),
    .io_core_dis_uops_1_valid(lsu_io_core_dis_uops_1_valid),
    .io_core_dis_uops_1_bits_switch(lsu_io_core_dis_uops_1_bits_switch),
    .io_core_dis_uops_1_bits_switch_off(lsu_io_core_dis_uops_1_bits_switch_off),
    .io_core_dis_uops_1_bits_is_unicore(lsu_io_core_dis_uops_1_bits_is_unicore),
    .io_core_dis_uops_1_bits_shift(lsu_io_core_dis_uops_1_bits_shift),
    .io_core_dis_uops_1_bits_lrs3_rtype(lsu_io_core_dis_uops_1_bits_lrs3_rtype),
    .io_core_dis_uops_1_bits_rflag(lsu_io_core_dis_uops_1_bits_rflag),
    .io_core_dis_uops_1_bits_wflag(lsu_io_core_dis_uops_1_bits_wflag),
    .io_core_dis_uops_1_bits_prflag(lsu_io_core_dis_uops_1_bits_prflag),
    .io_core_dis_uops_1_bits_pwflag(lsu_io_core_dis_uops_1_bits_pwflag),
    .io_core_dis_uops_1_bits_pflag_busy(lsu_io_core_dis_uops_1_bits_pflag_busy),
    .io_core_dis_uops_1_bits_stale_pflag(lsu_io_core_dis_uops_1_bits_stale_pflag),
    .io_core_dis_uops_1_bits_op1_sel(lsu_io_core_dis_uops_1_bits_op1_sel),
    .io_core_dis_uops_1_bits_op2_sel(lsu_io_core_dis_uops_1_bits_op2_sel),
    .io_core_dis_uops_1_bits_split_num(lsu_io_core_dis_uops_1_bits_split_num),
    .io_core_dis_uops_1_bits_self_index(lsu_io_core_dis_uops_1_bits_self_index),
    .io_core_dis_uops_1_bits_rob_inst_idx(lsu_io_core_dis_uops_1_bits_rob_inst_idx),
    .io_core_dis_uops_1_bits_address_num(lsu_io_core_dis_uops_1_bits_address_num),
    .io_core_dis_uops_1_bits_uopc(lsu_io_core_dis_uops_1_bits_uopc),
    .io_core_dis_uops_1_bits_inst(lsu_io_core_dis_uops_1_bits_inst),
    .io_core_dis_uops_1_bits_debug_inst(lsu_io_core_dis_uops_1_bits_debug_inst),
    .io_core_dis_uops_1_bits_is_rvc(lsu_io_core_dis_uops_1_bits_is_rvc),
    .io_core_dis_uops_1_bits_debug_pc(lsu_io_core_dis_uops_1_bits_debug_pc),
    .io_core_dis_uops_1_bits_iq_type(lsu_io_core_dis_uops_1_bits_iq_type),
    .io_core_dis_uops_1_bits_fu_code(lsu_io_core_dis_uops_1_bits_fu_code),
    .io_core_dis_uops_1_bits_ctrl_br_type(lsu_io_core_dis_uops_1_bits_ctrl_br_type),
    .io_core_dis_uops_1_bits_ctrl_op1_sel(lsu_io_core_dis_uops_1_bits_ctrl_op1_sel),
    .io_core_dis_uops_1_bits_ctrl_op2_sel(lsu_io_core_dis_uops_1_bits_ctrl_op2_sel),
    .io_core_dis_uops_1_bits_ctrl_imm_sel(lsu_io_core_dis_uops_1_bits_ctrl_imm_sel),
    .io_core_dis_uops_1_bits_ctrl_op_fcn(lsu_io_core_dis_uops_1_bits_ctrl_op_fcn),
    .io_core_dis_uops_1_bits_ctrl_fcn_dw(lsu_io_core_dis_uops_1_bits_ctrl_fcn_dw),
    .io_core_dis_uops_1_bits_ctrl_csr_cmd(lsu_io_core_dis_uops_1_bits_ctrl_csr_cmd),
    .io_core_dis_uops_1_bits_ctrl_is_load(lsu_io_core_dis_uops_1_bits_ctrl_is_load),
    .io_core_dis_uops_1_bits_ctrl_is_sta(lsu_io_core_dis_uops_1_bits_ctrl_is_sta),
    .io_core_dis_uops_1_bits_ctrl_is_std(lsu_io_core_dis_uops_1_bits_ctrl_is_std),
    .io_core_dis_uops_1_bits_ctrl_op3_sel(lsu_io_core_dis_uops_1_bits_ctrl_op3_sel),
    .io_core_dis_uops_1_bits_iw_state(lsu_io_core_dis_uops_1_bits_iw_state),
    .io_core_dis_uops_1_bits_iw_p1_poisoned(lsu_io_core_dis_uops_1_bits_iw_p1_poisoned),
    .io_core_dis_uops_1_bits_iw_p2_poisoned(lsu_io_core_dis_uops_1_bits_iw_p2_poisoned),
    .io_core_dis_uops_1_bits_is_br(lsu_io_core_dis_uops_1_bits_is_br),
    .io_core_dis_uops_1_bits_is_jalr(lsu_io_core_dis_uops_1_bits_is_jalr),
    .io_core_dis_uops_1_bits_is_jal(lsu_io_core_dis_uops_1_bits_is_jal),
    .io_core_dis_uops_1_bits_is_sfb(lsu_io_core_dis_uops_1_bits_is_sfb),
    .io_core_dis_uops_1_bits_br_mask(lsu_io_core_dis_uops_1_bits_br_mask),
    .io_core_dis_uops_1_bits_br_tag(lsu_io_core_dis_uops_1_bits_br_tag),
    .io_core_dis_uops_1_bits_ftq_idx(lsu_io_core_dis_uops_1_bits_ftq_idx),
    .io_core_dis_uops_1_bits_edge_inst(lsu_io_core_dis_uops_1_bits_edge_inst),
    .io_core_dis_uops_1_bits_pc_lob(lsu_io_core_dis_uops_1_bits_pc_lob),
    .io_core_dis_uops_1_bits_taken(lsu_io_core_dis_uops_1_bits_taken),
    .io_core_dis_uops_1_bits_imm_packed(lsu_io_core_dis_uops_1_bits_imm_packed),
    .io_core_dis_uops_1_bits_csr_addr(lsu_io_core_dis_uops_1_bits_csr_addr),
    .io_core_dis_uops_1_bits_rob_idx(lsu_io_core_dis_uops_1_bits_rob_idx),
    .io_core_dis_uops_1_bits_ldq_idx(lsu_io_core_dis_uops_1_bits_ldq_idx),
    .io_core_dis_uops_1_bits_stq_idx(lsu_io_core_dis_uops_1_bits_stq_idx),
    .io_core_dis_uops_1_bits_rxq_idx(lsu_io_core_dis_uops_1_bits_rxq_idx),
    .io_core_dis_uops_1_bits_pdst(lsu_io_core_dis_uops_1_bits_pdst),
    .io_core_dis_uops_1_bits_prs1(lsu_io_core_dis_uops_1_bits_prs1),
    .io_core_dis_uops_1_bits_prs2(lsu_io_core_dis_uops_1_bits_prs2),
    .io_core_dis_uops_1_bits_prs3(lsu_io_core_dis_uops_1_bits_prs3),
    .io_core_dis_uops_1_bits_ppred(lsu_io_core_dis_uops_1_bits_ppred),
    .io_core_dis_uops_1_bits_prs1_busy(lsu_io_core_dis_uops_1_bits_prs1_busy),
    .io_core_dis_uops_1_bits_prs2_busy(lsu_io_core_dis_uops_1_bits_prs2_busy),
    .io_core_dis_uops_1_bits_prs3_busy(lsu_io_core_dis_uops_1_bits_prs3_busy),
    .io_core_dis_uops_1_bits_ppred_busy(lsu_io_core_dis_uops_1_bits_ppred_busy),
    .io_core_dis_uops_1_bits_stale_pdst(lsu_io_core_dis_uops_1_bits_stale_pdst),
    .io_core_dis_uops_1_bits_exception(lsu_io_core_dis_uops_1_bits_exception),
    .io_core_dis_uops_1_bits_exc_cause(lsu_io_core_dis_uops_1_bits_exc_cause),
    .io_core_dis_uops_1_bits_bypassable(lsu_io_core_dis_uops_1_bits_bypassable),
    .io_core_dis_uops_1_bits_mem_cmd(lsu_io_core_dis_uops_1_bits_mem_cmd),
    .io_core_dis_uops_1_bits_mem_size(lsu_io_core_dis_uops_1_bits_mem_size),
    .io_core_dis_uops_1_bits_mem_signed(lsu_io_core_dis_uops_1_bits_mem_signed),
    .io_core_dis_uops_1_bits_is_fence(lsu_io_core_dis_uops_1_bits_is_fence),
    .io_core_dis_uops_1_bits_is_fencei(lsu_io_core_dis_uops_1_bits_is_fencei),
    .io_core_dis_uops_1_bits_is_amo(lsu_io_core_dis_uops_1_bits_is_amo),
    .io_core_dis_uops_1_bits_uses_ldq(lsu_io_core_dis_uops_1_bits_uses_ldq),
    .io_core_dis_uops_1_bits_uses_stq(lsu_io_core_dis_uops_1_bits_uses_stq),
    .io_core_dis_uops_1_bits_is_sys_pc2epc(lsu_io_core_dis_uops_1_bits_is_sys_pc2epc),
    .io_core_dis_uops_1_bits_is_unique(lsu_io_core_dis_uops_1_bits_is_unique),
    .io_core_dis_uops_1_bits_flush_on_commit(lsu_io_core_dis_uops_1_bits_flush_on_commit),
    .io_core_dis_uops_1_bits_ldst_is_rs1(lsu_io_core_dis_uops_1_bits_ldst_is_rs1),
    .io_core_dis_uops_1_bits_ldst(lsu_io_core_dis_uops_1_bits_ldst),
    .io_core_dis_uops_1_bits_lrs1(lsu_io_core_dis_uops_1_bits_lrs1),
    .io_core_dis_uops_1_bits_lrs2(lsu_io_core_dis_uops_1_bits_lrs2),
    .io_core_dis_uops_1_bits_lrs3(lsu_io_core_dis_uops_1_bits_lrs3),
    .io_core_dis_uops_1_bits_ldst_val(lsu_io_core_dis_uops_1_bits_ldst_val),
    .io_core_dis_uops_1_bits_dst_rtype(lsu_io_core_dis_uops_1_bits_dst_rtype),
    .io_core_dis_uops_1_bits_lrs1_rtype(lsu_io_core_dis_uops_1_bits_lrs1_rtype),
    .io_core_dis_uops_1_bits_lrs2_rtype(lsu_io_core_dis_uops_1_bits_lrs2_rtype),
    .io_core_dis_uops_1_bits_frs3_en(lsu_io_core_dis_uops_1_bits_frs3_en),
    .io_core_dis_uops_1_bits_fp_val(lsu_io_core_dis_uops_1_bits_fp_val),
    .io_core_dis_uops_1_bits_fp_single(lsu_io_core_dis_uops_1_bits_fp_single),
    .io_core_dis_uops_1_bits_xcpt_pf_if(lsu_io_core_dis_uops_1_bits_xcpt_pf_if),
    .io_core_dis_uops_1_bits_xcpt_ae_if(lsu_io_core_dis_uops_1_bits_xcpt_ae_if),
    .io_core_dis_uops_1_bits_xcpt_ma_if(lsu_io_core_dis_uops_1_bits_xcpt_ma_if),
    .io_core_dis_uops_1_bits_bp_debug_if(lsu_io_core_dis_uops_1_bits_bp_debug_if),
    .io_core_dis_uops_1_bits_bp_xcpt_if(lsu_io_core_dis_uops_1_bits_bp_xcpt_if),
    .io_core_dis_uops_1_bits_debug_fsrc(lsu_io_core_dis_uops_1_bits_debug_fsrc),
    .io_core_dis_uops_1_bits_debug_tsrc(lsu_io_core_dis_uops_1_bits_debug_tsrc),
    .io_core_dis_ldq_idx_0(lsu_io_core_dis_ldq_idx_0),
    .io_core_dis_ldq_idx_1(lsu_io_core_dis_ldq_idx_1),
    .io_core_dis_stq_idx_0(lsu_io_core_dis_stq_idx_0),
    .io_core_dis_stq_idx_1(lsu_io_core_dis_stq_idx_1),
    .io_core_ldq_full_0(lsu_io_core_ldq_full_0),
    .io_core_ldq_full_1(lsu_io_core_ldq_full_1),
    .io_core_stq_full_0(lsu_io_core_stq_full_0),
    .io_core_stq_full_1(lsu_io_core_stq_full_1),
    .io_core_fp_stdata_ready(lsu_io_core_fp_stdata_ready),
    .io_core_fp_stdata_valid(lsu_io_core_fp_stdata_valid),
    .io_core_fp_stdata_bits_uop_switch(lsu_io_core_fp_stdata_bits_uop_switch),
    .io_core_fp_stdata_bits_uop_switch_off(lsu_io_core_fp_stdata_bits_uop_switch_off),
    .io_core_fp_stdata_bits_uop_is_unicore(lsu_io_core_fp_stdata_bits_uop_is_unicore),
    .io_core_fp_stdata_bits_uop_shift(lsu_io_core_fp_stdata_bits_uop_shift),
    .io_core_fp_stdata_bits_uop_lrs3_rtype(lsu_io_core_fp_stdata_bits_uop_lrs3_rtype),
    .io_core_fp_stdata_bits_uop_rflag(lsu_io_core_fp_stdata_bits_uop_rflag),
    .io_core_fp_stdata_bits_uop_wflag(lsu_io_core_fp_stdata_bits_uop_wflag),
    .io_core_fp_stdata_bits_uop_prflag(lsu_io_core_fp_stdata_bits_uop_prflag),
    .io_core_fp_stdata_bits_uop_pwflag(lsu_io_core_fp_stdata_bits_uop_pwflag),
    .io_core_fp_stdata_bits_uop_pflag_busy(lsu_io_core_fp_stdata_bits_uop_pflag_busy),
    .io_core_fp_stdata_bits_uop_stale_pflag(lsu_io_core_fp_stdata_bits_uop_stale_pflag),
    .io_core_fp_stdata_bits_uop_op1_sel(lsu_io_core_fp_stdata_bits_uop_op1_sel),
    .io_core_fp_stdata_bits_uop_op2_sel(lsu_io_core_fp_stdata_bits_uop_op2_sel),
    .io_core_fp_stdata_bits_uop_split_num(lsu_io_core_fp_stdata_bits_uop_split_num),
    .io_core_fp_stdata_bits_uop_self_index(lsu_io_core_fp_stdata_bits_uop_self_index),
    .io_core_fp_stdata_bits_uop_rob_inst_idx(lsu_io_core_fp_stdata_bits_uop_rob_inst_idx),
    .io_core_fp_stdata_bits_uop_address_num(lsu_io_core_fp_stdata_bits_uop_address_num),
    .io_core_fp_stdata_bits_uop_uopc(lsu_io_core_fp_stdata_bits_uop_uopc),
    .io_core_fp_stdata_bits_uop_inst(lsu_io_core_fp_stdata_bits_uop_inst),
    .io_core_fp_stdata_bits_uop_debug_inst(lsu_io_core_fp_stdata_bits_uop_debug_inst),
    .io_core_fp_stdata_bits_uop_is_rvc(lsu_io_core_fp_stdata_bits_uop_is_rvc),
    .io_core_fp_stdata_bits_uop_debug_pc(lsu_io_core_fp_stdata_bits_uop_debug_pc),
    .io_core_fp_stdata_bits_uop_iq_type(lsu_io_core_fp_stdata_bits_uop_iq_type),
    .io_core_fp_stdata_bits_uop_fu_code(lsu_io_core_fp_stdata_bits_uop_fu_code),
    .io_core_fp_stdata_bits_uop_ctrl_br_type(lsu_io_core_fp_stdata_bits_uop_ctrl_br_type),
    .io_core_fp_stdata_bits_uop_ctrl_op1_sel(lsu_io_core_fp_stdata_bits_uop_ctrl_op1_sel),
    .io_core_fp_stdata_bits_uop_ctrl_op2_sel(lsu_io_core_fp_stdata_bits_uop_ctrl_op2_sel),
    .io_core_fp_stdata_bits_uop_ctrl_imm_sel(lsu_io_core_fp_stdata_bits_uop_ctrl_imm_sel),
    .io_core_fp_stdata_bits_uop_ctrl_op_fcn(lsu_io_core_fp_stdata_bits_uop_ctrl_op_fcn),
    .io_core_fp_stdata_bits_uop_ctrl_fcn_dw(lsu_io_core_fp_stdata_bits_uop_ctrl_fcn_dw),
    .io_core_fp_stdata_bits_uop_ctrl_csr_cmd(lsu_io_core_fp_stdata_bits_uop_ctrl_csr_cmd),
    .io_core_fp_stdata_bits_uop_ctrl_is_load(lsu_io_core_fp_stdata_bits_uop_ctrl_is_load),
    .io_core_fp_stdata_bits_uop_ctrl_is_sta(lsu_io_core_fp_stdata_bits_uop_ctrl_is_sta),
    .io_core_fp_stdata_bits_uop_ctrl_is_std(lsu_io_core_fp_stdata_bits_uop_ctrl_is_std),
    .io_core_fp_stdata_bits_uop_ctrl_op3_sel(lsu_io_core_fp_stdata_bits_uop_ctrl_op3_sel),
    .io_core_fp_stdata_bits_uop_iw_state(lsu_io_core_fp_stdata_bits_uop_iw_state),
    .io_core_fp_stdata_bits_uop_iw_p1_poisoned(lsu_io_core_fp_stdata_bits_uop_iw_p1_poisoned),
    .io_core_fp_stdata_bits_uop_iw_p2_poisoned(lsu_io_core_fp_stdata_bits_uop_iw_p2_poisoned),
    .io_core_fp_stdata_bits_uop_is_br(lsu_io_core_fp_stdata_bits_uop_is_br),
    .io_core_fp_stdata_bits_uop_is_jalr(lsu_io_core_fp_stdata_bits_uop_is_jalr),
    .io_core_fp_stdata_bits_uop_is_jal(lsu_io_core_fp_stdata_bits_uop_is_jal),
    .io_core_fp_stdata_bits_uop_is_sfb(lsu_io_core_fp_stdata_bits_uop_is_sfb),
    .io_core_fp_stdata_bits_uop_br_mask(lsu_io_core_fp_stdata_bits_uop_br_mask),
    .io_core_fp_stdata_bits_uop_br_tag(lsu_io_core_fp_stdata_bits_uop_br_tag),
    .io_core_fp_stdata_bits_uop_ftq_idx(lsu_io_core_fp_stdata_bits_uop_ftq_idx),
    .io_core_fp_stdata_bits_uop_edge_inst(lsu_io_core_fp_stdata_bits_uop_edge_inst),
    .io_core_fp_stdata_bits_uop_pc_lob(lsu_io_core_fp_stdata_bits_uop_pc_lob),
    .io_core_fp_stdata_bits_uop_taken(lsu_io_core_fp_stdata_bits_uop_taken),
    .io_core_fp_stdata_bits_uop_imm_packed(lsu_io_core_fp_stdata_bits_uop_imm_packed),
    .io_core_fp_stdata_bits_uop_csr_addr(lsu_io_core_fp_stdata_bits_uop_csr_addr),
    .io_core_fp_stdata_bits_uop_rob_idx(lsu_io_core_fp_stdata_bits_uop_rob_idx),
    .io_core_fp_stdata_bits_uop_ldq_idx(lsu_io_core_fp_stdata_bits_uop_ldq_idx),
    .io_core_fp_stdata_bits_uop_stq_idx(lsu_io_core_fp_stdata_bits_uop_stq_idx),
    .io_core_fp_stdata_bits_uop_rxq_idx(lsu_io_core_fp_stdata_bits_uop_rxq_idx),
    .io_core_fp_stdata_bits_uop_pdst(lsu_io_core_fp_stdata_bits_uop_pdst),
    .io_core_fp_stdata_bits_uop_prs1(lsu_io_core_fp_stdata_bits_uop_prs1),
    .io_core_fp_stdata_bits_uop_prs2(lsu_io_core_fp_stdata_bits_uop_prs2),
    .io_core_fp_stdata_bits_uop_prs3(lsu_io_core_fp_stdata_bits_uop_prs3),
    .io_core_fp_stdata_bits_uop_ppred(lsu_io_core_fp_stdata_bits_uop_ppred),
    .io_core_fp_stdata_bits_uop_prs1_busy(lsu_io_core_fp_stdata_bits_uop_prs1_busy),
    .io_core_fp_stdata_bits_uop_prs2_busy(lsu_io_core_fp_stdata_bits_uop_prs2_busy),
    .io_core_fp_stdata_bits_uop_prs3_busy(lsu_io_core_fp_stdata_bits_uop_prs3_busy),
    .io_core_fp_stdata_bits_uop_ppred_busy(lsu_io_core_fp_stdata_bits_uop_ppred_busy),
    .io_core_fp_stdata_bits_uop_stale_pdst(lsu_io_core_fp_stdata_bits_uop_stale_pdst),
    .io_core_fp_stdata_bits_uop_exception(lsu_io_core_fp_stdata_bits_uop_exception),
    .io_core_fp_stdata_bits_uop_exc_cause(lsu_io_core_fp_stdata_bits_uop_exc_cause),
    .io_core_fp_stdata_bits_uop_bypassable(lsu_io_core_fp_stdata_bits_uop_bypassable),
    .io_core_fp_stdata_bits_uop_mem_cmd(lsu_io_core_fp_stdata_bits_uop_mem_cmd),
    .io_core_fp_stdata_bits_uop_mem_size(lsu_io_core_fp_stdata_bits_uop_mem_size),
    .io_core_fp_stdata_bits_uop_mem_signed(lsu_io_core_fp_stdata_bits_uop_mem_signed),
    .io_core_fp_stdata_bits_uop_is_fence(lsu_io_core_fp_stdata_bits_uop_is_fence),
    .io_core_fp_stdata_bits_uop_is_fencei(lsu_io_core_fp_stdata_bits_uop_is_fencei),
    .io_core_fp_stdata_bits_uop_is_amo(lsu_io_core_fp_stdata_bits_uop_is_amo),
    .io_core_fp_stdata_bits_uop_uses_ldq(lsu_io_core_fp_stdata_bits_uop_uses_ldq),
    .io_core_fp_stdata_bits_uop_uses_stq(lsu_io_core_fp_stdata_bits_uop_uses_stq),
    .io_core_fp_stdata_bits_uop_is_sys_pc2epc(lsu_io_core_fp_stdata_bits_uop_is_sys_pc2epc),
    .io_core_fp_stdata_bits_uop_is_unique(lsu_io_core_fp_stdata_bits_uop_is_unique),
    .io_core_fp_stdata_bits_uop_flush_on_commit(lsu_io_core_fp_stdata_bits_uop_flush_on_commit),
    .io_core_fp_stdata_bits_uop_ldst_is_rs1(lsu_io_core_fp_stdata_bits_uop_ldst_is_rs1),
    .io_core_fp_stdata_bits_uop_ldst(lsu_io_core_fp_stdata_bits_uop_ldst),
    .io_core_fp_stdata_bits_uop_lrs1(lsu_io_core_fp_stdata_bits_uop_lrs1),
    .io_core_fp_stdata_bits_uop_lrs2(lsu_io_core_fp_stdata_bits_uop_lrs2),
    .io_core_fp_stdata_bits_uop_lrs3(lsu_io_core_fp_stdata_bits_uop_lrs3),
    .io_core_fp_stdata_bits_uop_ldst_val(lsu_io_core_fp_stdata_bits_uop_ldst_val),
    .io_core_fp_stdata_bits_uop_dst_rtype(lsu_io_core_fp_stdata_bits_uop_dst_rtype),
    .io_core_fp_stdata_bits_uop_lrs1_rtype(lsu_io_core_fp_stdata_bits_uop_lrs1_rtype),
    .io_core_fp_stdata_bits_uop_lrs2_rtype(lsu_io_core_fp_stdata_bits_uop_lrs2_rtype),
    .io_core_fp_stdata_bits_uop_frs3_en(lsu_io_core_fp_stdata_bits_uop_frs3_en),
    .io_core_fp_stdata_bits_uop_fp_val(lsu_io_core_fp_stdata_bits_uop_fp_val),
    .io_core_fp_stdata_bits_uop_fp_single(lsu_io_core_fp_stdata_bits_uop_fp_single),
    .io_core_fp_stdata_bits_uop_xcpt_pf_if(lsu_io_core_fp_stdata_bits_uop_xcpt_pf_if),
    .io_core_fp_stdata_bits_uop_xcpt_ae_if(lsu_io_core_fp_stdata_bits_uop_xcpt_ae_if),
    .io_core_fp_stdata_bits_uop_xcpt_ma_if(lsu_io_core_fp_stdata_bits_uop_xcpt_ma_if),
    .io_core_fp_stdata_bits_uop_bp_debug_if(lsu_io_core_fp_stdata_bits_uop_bp_debug_if),
    .io_core_fp_stdata_bits_uop_bp_xcpt_if(lsu_io_core_fp_stdata_bits_uop_bp_xcpt_if),
    .io_core_fp_stdata_bits_uop_debug_fsrc(lsu_io_core_fp_stdata_bits_uop_debug_fsrc),
    .io_core_fp_stdata_bits_uop_debug_tsrc(lsu_io_core_fp_stdata_bits_uop_debug_tsrc),
    .io_core_fp_stdata_bits_data(lsu_io_core_fp_stdata_bits_data),
    .io_core_fp_stdata_bits_predicated(lsu_io_core_fp_stdata_bits_predicated),
    .io_core_fp_stdata_bits_fflags_valid(lsu_io_core_fp_stdata_bits_fflags_valid),
    .io_core_fp_stdata_bits_fflags_bits_uop_switch(lsu_io_core_fp_stdata_bits_fflags_bits_uop_switch),
    .io_core_fp_stdata_bits_fflags_bits_uop_switch_off(lsu_io_core_fp_stdata_bits_fflags_bits_uop_switch_off),
    .io_core_fp_stdata_bits_fflags_bits_uop_is_unicore(lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_unicore),
    .io_core_fp_stdata_bits_fflags_bits_uop_shift(lsu_io_core_fp_stdata_bits_fflags_bits_uop_shift),
    .io_core_fp_stdata_bits_fflags_bits_uop_lrs3_rtype(lsu_io_core_fp_stdata_bits_fflags_bits_uop_lrs3_rtype),
    .io_core_fp_stdata_bits_fflags_bits_uop_rflag(lsu_io_core_fp_stdata_bits_fflags_bits_uop_rflag),
    .io_core_fp_stdata_bits_fflags_bits_uop_wflag(lsu_io_core_fp_stdata_bits_fflags_bits_uop_wflag),
    .io_core_fp_stdata_bits_fflags_bits_uop_prflag(lsu_io_core_fp_stdata_bits_fflags_bits_uop_prflag),
    .io_core_fp_stdata_bits_fflags_bits_uop_pwflag(lsu_io_core_fp_stdata_bits_fflags_bits_uop_pwflag),
    .io_core_fp_stdata_bits_fflags_bits_uop_pflag_busy(lsu_io_core_fp_stdata_bits_fflags_bits_uop_pflag_busy),
    .io_core_fp_stdata_bits_fflags_bits_uop_stale_pflag(lsu_io_core_fp_stdata_bits_fflags_bits_uop_stale_pflag),
    .io_core_fp_stdata_bits_fflags_bits_uop_op1_sel(lsu_io_core_fp_stdata_bits_fflags_bits_uop_op1_sel),
    .io_core_fp_stdata_bits_fflags_bits_uop_op2_sel(lsu_io_core_fp_stdata_bits_fflags_bits_uop_op2_sel),
    .io_core_fp_stdata_bits_fflags_bits_uop_split_num(lsu_io_core_fp_stdata_bits_fflags_bits_uop_split_num),
    .io_core_fp_stdata_bits_fflags_bits_uop_self_index(lsu_io_core_fp_stdata_bits_fflags_bits_uop_self_index),
    .io_core_fp_stdata_bits_fflags_bits_uop_rob_inst_idx(lsu_io_core_fp_stdata_bits_fflags_bits_uop_rob_inst_idx),
    .io_core_fp_stdata_bits_fflags_bits_uop_address_num(lsu_io_core_fp_stdata_bits_fflags_bits_uop_address_num),
    .io_core_fp_stdata_bits_fflags_bits_uop_uopc(lsu_io_core_fp_stdata_bits_fflags_bits_uop_uopc),
    .io_core_fp_stdata_bits_fflags_bits_uop_inst(lsu_io_core_fp_stdata_bits_fflags_bits_uop_inst),
    .io_core_fp_stdata_bits_fflags_bits_uop_debug_inst(lsu_io_core_fp_stdata_bits_fflags_bits_uop_debug_inst),
    .io_core_fp_stdata_bits_fflags_bits_uop_is_rvc(lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_rvc),
    .io_core_fp_stdata_bits_fflags_bits_uop_debug_pc(lsu_io_core_fp_stdata_bits_fflags_bits_uop_debug_pc),
    .io_core_fp_stdata_bits_fflags_bits_uop_iq_type(lsu_io_core_fp_stdata_bits_fflags_bits_uop_iq_type),
    .io_core_fp_stdata_bits_fflags_bits_uop_fu_code(lsu_io_core_fp_stdata_bits_fflags_bits_uop_fu_code),
    .io_core_fp_stdata_bits_fflags_bits_uop_ctrl_br_type(lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_br_type),
    .io_core_fp_stdata_bits_fflags_bits_uop_ctrl_op1_sel(lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_op1_sel),
    .io_core_fp_stdata_bits_fflags_bits_uop_ctrl_op2_sel(lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_op2_sel),
    .io_core_fp_stdata_bits_fflags_bits_uop_ctrl_imm_sel(lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_imm_sel),
    .io_core_fp_stdata_bits_fflags_bits_uop_ctrl_op_fcn(lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_op_fcn),
    .io_core_fp_stdata_bits_fflags_bits_uop_ctrl_fcn_dw(lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_fcn_dw),
    .io_core_fp_stdata_bits_fflags_bits_uop_ctrl_csr_cmd(lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_csr_cmd),
    .io_core_fp_stdata_bits_fflags_bits_uop_ctrl_is_load(lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_is_load),
    .io_core_fp_stdata_bits_fflags_bits_uop_ctrl_is_sta(lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_is_sta),
    .io_core_fp_stdata_bits_fflags_bits_uop_ctrl_is_std(lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_is_std),
    .io_core_fp_stdata_bits_fflags_bits_uop_ctrl_op3_sel(lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_op3_sel),
    .io_core_fp_stdata_bits_fflags_bits_uop_iw_state(lsu_io_core_fp_stdata_bits_fflags_bits_uop_iw_state),
    .io_core_fp_stdata_bits_fflags_bits_uop_iw_p1_poisoned(lsu_io_core_fp_stdata_bits_fflags_bits_uop_iw_p1_poisoned),
    .io_core_fp_stdata_bits_fflags_bits_uop_iw_p2_poisoned(lsu_io_core_fp_stdata_bits_fflags_bits_uop_iw_p2_poisoned),
    .io_core_fp_stdata_bits_fflags_bits_uop_is_br(lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_br),
    .io_core_fp_stdata_bits_fflags_bits_uop_is_jalr(lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_jalr),
    .io_core_fp_stdata_bits_fflags_bits_uop_is_jal(lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_jal),
    .io_core_fp_stdata_bits_fflags_bits_uop_is_sfb(lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_sfb),
    .io_core_fp_stdata_bits_fflags_bits_uop_br_mask(lsu_io_core_fp_stdata_bits_fflags_bits_uop_br_mask),
    .io_core_fp_stdata_bits_fflags_bits_uop_br_tag(lsu_io_core_fp_stdata_bits_fflags_bits_uop_br_tag),
    .io_core_fp_stdata_bits_fflags_bits_uop_ftq_idx(lsu_io_core_fp_stdata_bits_fflags_bits_uop_ftq_idx),
    .io_core_fp_stdata_bits_fflags_bits_uop_edge_inst(lsu_io_core_fp_stdata_bits_fflags_bits_uop_edge_inst),
    .io_core_fp_stdata_bits_fflags_bits_uop_pc_lob(lsu_io_core_fp_stdata_bits_fflags_bits_uop_pc_lob),
    .io_core_fp_stdata_bits_fflags_bits_uop_taken(lsu_io_core_fp_stdata_bits_fflags_bits_uop_taken),
    .io_core_fp_stdata_bits_fflags_bits_uop_imm_packed(lsu_io_core_fp_stdata_bits_fflags_bits_uop_imm_packed),
    .io_core_fp_stdata_bits_fflags_bits_uop_csr_addr(lsu_io_core_fp_stdata_bits_fflags_bits_uop_csr_addr),
    .io_core_fp_stdata_bits_fflags_bits_uop_rob_idx(lsu_io_core_fp_stdata_bits_fflags_bits_uop_rob_idx),
    .io_core_fp_stdata_bits_fflags_bits_uop_ldq_idx(lsu_io_core_fp_stdata_bits_fflags_bits_uop_ldq_idx),
    .io_core_fp_stdata_bits_fflags_bits_uop_stq_idx(lsu_io_core_fp_stdata_bits_fflags_bits_uop_stq_idx),
    .io_core_fp_stdata_bits_fflags_bits_uop_rxq_idx(lsu_io_core_fp_stdata_bits_fflags_bits_uop_rxq_idx),
    .io_core_fp_stdata_bits_fflags_bits_uop_pdst(lsu_io_core_fp_stdata_bits_fflags_bits_uop_pdst),
    .io_core_fp_stdata_bits_fflags_bits_uop_prs1(lsu_io_core_fp_stdata_bits_fflags_bits_uop_prs1),
    .io_core_fp_stdata_bits_fflags_bits_uop_prs2(lsu_io_core_fp_stdata_bits_fflags_bits_uop_prs2),
    .io_core_fp_stdata_bits_fflags_bits_uop_prs3(lsu_io_core_fp_stdata_bits_fflags_bits_uop_prs3),
    .io_core_fp_stdata_bits_fflags_bits_uop_ppred(lsu_io_core_fp_stdata_bits_fflags_bits_uop_ppred),
    .io_core_fp_stdata_bits_fflags_bits_uop_prs1_busy(lsu_io_core_fp_stdata_bits_fflags_bits_uop_prs1_busy),
    .io_core_fp_stdata_bits_fflags_bits_uop_prs2_busy(lsu_io_core_fp_stdata_bits_fflags_bits_uop_prs2_busy),
    .io_core_fp_stdata_bits_fflags_bits_uop_prs3_busy(lsu_io_core_fp_stdata_bits_fflags_bits_uop_prs3_busy),
    .io_core_fp_stdata_bits_fflags_bits_uop_ppred_busy(lsu_io_core_fp_stdata_bits_fflags_bits_uop_ppred_busy),
    .io_core_fp_stdata_bits_fflags_bits_uop_stale_pdst(lsu_io_core_fp_stdata_bits_fflags_bits_uop_stale_pdst),
    .io_core_fp_stdata_bits_fflags_bits_uop_exception(lsu_io_core_fp_stdata_bits_fflags_bits_uop_exception),
    .io_core_fp_stdata_bits_fflags_bits_uop_exc_cause(lsu_io_core_fp_stdata_bits_fflags_bits_uop_exc_cause),
    .io_core_fp_stdata_bits_fflags_bits_uop_bypassable(lsu_io_core_fp_stdata_bits_fflags_bits_uop_bypassable),
    .io_core_fp_stdata_bits_fflags_bits_uop_mem_cmd(lsu_io_core_fp_stdata_bits_fflags_bits_uop_mem_cmd),
    .io_core_fp_stdata_bits_fflags_bits_uop_mem_size(lsu_io_core_fp_stdata_bits_fflags_bits_uop_mem_size),
    .io_core_fp_stdata_bits_fflags_bits_uop_mem_signed(lsu_io_core_fp_stdata_bits_fflags_bits_uop_mem_signed),
    .io_core_fp_stdata_bits_fflags_bits_uop_is_fence(lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_fence),
    .io_core_fp_stdata_bits_fflags_bits_uop_is_fencei(lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_fencei),
    .io_core_fp_stdata_bits_fflags_bits_uop_is_amo(lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_amo),
    .io_core_fp_stdata_bits_fflags_bits_uop_uses_ldq(lsu_io_core_fp_stdata_bits_fflags_bits_uop_uses_ldq),
    .io_core_fp_stdata_bits_fflags_bits_uop_uses_stq(lsu_io_core_fp_stdata_bits_fflags_bits_uop_uses_stq),
    .io_core_fp_stdata_bits_fflags_bits_uop_is_sys_pc2epc(lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_sys_pc2epc),
    .io_core_fp_stdata_bits_fflags_bits_uop_is_unique(lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_unique),
    .io_core_fp_stdata_bits_fflags_bits_uop_flush_on_commit(lsu_io_core_fp_stdata_bits_fflags_bits_uop_flush_on_commit),
    .io_core_fp_stdata_bits_fflags_bits_uop_ldst_is_rs1(lsu_io_core_fp_stdata_bits_fflags_bits_uop_ldst_is_rs1),
    .io_core_fp_stdata_bits_fflags_bits_uop_ldst(lsu_io_core_fp_stdata_bits_fflags_bits_uop_ldst),
    .io_core_fp_stdata_bits_fflags_bits_uop_lrs1(lsu_io_core_fp_stdata_bits_fflags_bits_uop_lrs1),
    .io_core_fp_stdata_bits_fflags_bits_uop_lrs2(lsu_io_core_fp_stdata_bits_fflags_bits_uop_lrs2),
    .io_core_fp_stdata_bits_fflags_bits_uop_lrs3(lsu_io_core_fp_stdata_bits_fflags_bits_uop_lrs3),
    .io_core_fp_stdata_bits_fflags_bits_uop_ldst_val(lsu_io_core_fp_stdata_bits_fflags_bits_uop_ldst_val),
    .io_core_fp_stdata_bits_fflags_bits_uop_dst_rtype(lsu_io_core_fp_stdata_bits_fflags_bits_uop_dst_rtype),
    .io_core_fp_stdata_bits_fflags_bits_uop_lrs1_rtype(lsu_io_core_fp_stdata_bits_fflags_bits_uop_lrs1_rtype),
    .io_core_fp_stdata_bits_fflags_bits_uop_lrs2_rtype(lsu_io_core_fp_stdata_bits_fflags_bits_uop_lrs2_rtype),
    .io_core_fp_stdata_bits_fflags_bits_uop_frs3_en(lsu_io_core_fp_stdata_bits_fflags_bits_uop_frs3_en),
    .io_core_fp_stdata_bits_fflags_bits_uop_fp_val(lsu_io_core_fp_stdata_bits_fflags_bits_uop_fp_val),
    .io_core_fp_stdata_bits_fflags_bits_uop_fp_single(lsu_io_core_fp_stdata_bits_fflags_bits_uop_fp_single),
    .io_core_fp_stdata_bits_fflags_bits_uop_xcpt_pf_if(lsu_io_core_fp_stdata_bits_fflags_bits_uop_xcpt_pf_if),
    .io_core_fp_stdata_bits_fflags_bits_uop_xcpt_ae_if(lsu_io_core_fp_stdata_bits_fflags_bits_uop_xcpt_ae_if),
    .io_core_fp_stdata_bits_fflags_bits_uop_xcpt_ma_if(lsu_io_core_fp_stdata_bits_fflags_bits_uop_xcpt_ma_if),
    .io_core_fp_stdata_bits_fflags_bits_uop_bp_debug_if(lsu_io_core_fp_stdata_bits_fflags_bits_uop_bp_debug_if),
    .io_core_fp_stdata_bits_fflags_bits_uop_bp_xcpt_if(lsu_io_core_fp_stdata_bits_fflags_bits_uop_bp_xcpt_if),
    .io_core_fp_stdata_bits_fflags_bits_uop_debug_fsrc(lsu_io_core_fp_stdata_bits_fflags_bits_uop_debug_fsrc),
    .io_core_fp_stdata_bits_fflags_bits_uop_debug_tsrc(lsu_io_core_fp_stdata_bits_fflags_bits_uop_debug_tsrc),
    .io_core_fp_stdata_bits_fflags_bits_flags(lsu_io_core_fp_stdata_bits_fflags_bits_flags),
    .io_core_fp_stdata_bits_flagdata(lsu_io_core_fp_stdata_bits_flagdata),
    .io_core_fp_stdata_bits_fflagdata_valid(lsu_io_core_fp_stdata_bits_fflagdata_valid),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_switch(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_switch),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_switch_off(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_switch_off),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_is_unicore(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_unicore),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_shift(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_shift),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_lrs3_rtype(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_lrs3_rtype),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_rflag(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_rflag),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_wflag(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_wflag),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_prflag(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_prflag),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_pwflag(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_pwflag),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_pflag_busy(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_pflag_busy),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_stale_pflag(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_stale_pflag),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_op1_sel(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_op1_sel),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_op2_sel(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_op2_sel),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_split_num(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_split_num),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_self_index(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_self_index),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_rob_inst_idx(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_rob_inst_idx),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_address_num(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_address_num),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_uopc(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_uopc),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_inst(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_inst),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_debug_inst(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_debug_inst),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_is_rvc(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_rvc),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_debug_pc(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_debug_pc),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_iq_type(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_iq_type),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_fu_code(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_fu_code),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_br_type(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_br_type),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_op1_sel(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_op1_sel),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_op2_sel(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_op2_sel),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_imm_sel(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_imm_sel),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_op_fcn(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_op_fcn),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_fcn_dw(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_fcn_dw),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_csr_cmd(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_csr_cmd),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_load(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_load),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_sta(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_sta),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_std(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_std),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_op3_sel(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_op3_sel),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_iw_state(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_iw_state),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_iw_p1_poisoned(
      lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_iw_p1_poisoned),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_iw_p2_poisoned(
      lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_iw_p2_poisoned),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_is_br(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_br),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_is_jalr(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_jalr),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_is_jal(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_jal),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_is_sfb(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_sfb),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_br_mask(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_br_mask),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_br_tag(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_br_tag),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_ftq_idx(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ftq_idx),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_edge_inst(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_edge_inst),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_pc_lob(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_pc_lob),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_taken(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_taken),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_imm_packed(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_imm_packed),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_csr_addr(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_csr_addr),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_rob_idx(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_rob_idx),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_ldq_idx(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ldq_idx),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_stq_idx(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_stq_idx),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_rxq_idx(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_rxq_idx),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_pdst(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_pdst),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_prs1(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_prs1),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_prs2(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_prs2),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_prs3(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_prs3),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_ppred(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ppred),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_prs1_busy(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_prs1_busy),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_prs2_busy(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_prs2_busy),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_prs3_busy(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_prs3_busy),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_ppred_busy(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ppred_busy),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_stale_pdst(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_stale_pdst),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_exception(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_exception),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_exc_cause(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_exc_cause),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_bypassable(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_bypassable),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_mem_cmd(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_mem_cmd),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_mem_size(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_mem_size),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_mem_signed(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_mem_signed),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_is_fence(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_fence),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_is_fencei(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_fencei),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_is_amo(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_amo),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_uses_ldq(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_uses_ldq),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_uses_stq(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_uses_stq),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_is_sys_pc2epc(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_sys_pc2epc
      ),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_is_unique(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_unique),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_flush_on_commit(
      lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_flush_on_commit),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_ldst_is_rs1(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ldst_is_rs1),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_ldst(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ldst),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_lrs1(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_lrs1),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_lrs2(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_lrs2),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_lrs3(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_lrs3),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_ldst_val(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ldst_val),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_dst_rtype(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_dst_rtype),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_lrs1_rtype(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_lrs1_rtype),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_lrs2_rtype(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_lrs2_rtype),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_frs3_en(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_frs3_en),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_fp_val(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_fp_val),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_fp_single(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_fp_single),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_xcpt_pf_if(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_xcpt_pf_if),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_xcpt_ae_if(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_xcpt_ae_if),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_xcpt_ma_if(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_xcpt_ma_if),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_bp_debug_if(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_bp_debug_if),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_bp_xcpt_if(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_bp_xcpt_if),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_debug_fsrc(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_debug_fsrc),
    .io_core_fp_stdata_bits_fflagdata_bits_uop_debug_tsrc(lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_debug_tsrc),
    .io_core_fp_stdata_bits_fflagdata_bits_fflag(lsu_io_core_fp_stdata_bits_fflagdata_bits_fflag),
    .io_core_commit_valids_0(lsu_io_core_commit_valids_0),
    .io_core_commit_valids_1(lsu_io_core_commit_valids_1),
    .io_core_commit_arch_valids_0(lsu_io_core_commit_arch_valids_0),
    .io_core_commit_arch_valids_1(lsu_io_core_commit_arch_valids_1),
    .io_core_commit_uops_0_switch(lsu_io_core_commit_uops_0_switch),
    .io_core_commit_uops_0_switch_off(lsu_io_core_commit_uops_0_switch_off),
    .io_core_commit_uops_0_is_unicore(lsu_io_core_commit_uops_0_is_unicore),
    .io_core_commit_uops_0_shift(lsu_io_core_commit_uops_0_shift),
    .io_core_commit_uops_0_lrs3_rtype(lsu_io_core_commit_uops_0_lrs3_rtype),
    .io_core_commit_uops_0_rflag(lsu_io_core_commit_uops_0_rflag),
    .io_core_commit_uops_0_wflag(lsu_io_core_commit_uops_0_wflag),
    .io_core_commit_uops_0_prflag(lsu_io_core_commit_uops_0_prflag),
    .io_core_commit_uops_0_pwflag(lsu_io_core_commit_uops_0_pwflag),
    .io_core_commit_uops_0_pflag_busy(lsu_io_core_commit_uops_0_pflag_busy),
    .io_core_commit_uops_0_stale_pflag(lsu_io_core_commit_uops_0_stale_pflag),
    .io_core_commit_uops_0_op1_sel(lsu_io_core_commit_uops_0_op1_sel),
    .io_core_commit_uops_0_op2_sel(lsu_io_core_commit_uops_0_op2_sel),
    .io_core_commit_uops_0_split_num(lsu_io_core_commit_uops_0_split_num),
    .io_core_commit_uops_0_self_index(lsu_io_core_commit_uops_0_self_index),
    .io_core_commit_uops_0_rob_inst_idx(lsu_io_core_commit_uops_0_rob_inst_idx),
    .io_core_commit_uops_0_address_num(lsu_io_core_commit_uops_0_address_num),
    .io_core_commit_uops_0_uopc(lsu_io_core_commit_uops_0_uopc),
    .io_core_commit_uops_0_inst(lsu_io_core_commit_uops_0_inst),
    .io_core_commit_uops_0_debug_inst(lsu_io_core_commit_uops_0_debug_inst),
    .io_core_commit_uops_0_is_rvc(lsu_io_core_commit_uops_0_is_rvc),
    .io_core_commit_uops_0_debug_pc(lsu_io_core_commit_uops_0_debug_pc),
    .io_core_commit_uops_0_iq_type(lsu_io_core_commit_uops_0_iq_type),
    .io_core_commit_uops_0_fu_code(lsu_io_core_commit_uops_0_fu_code),
    .io_core_commit_uops_0_ctrl_br_type(lsu_io_core_commit_uops_0_ctrl_br_type),
    .io_core_commit_uops_0_ctrl_op1_sel(lsu_io_core_commit_uops_0_ctrl_op1_sel),
    .io_core_commit_uops_0_ctrl_op2_sel(lsu_io_core_commit_uops_0_ctrl_op2_sel),
    .io_core_commit_uops_0_ctrl_imm_sel(lsu_io_core_commit_uops_0_ctrl_imm_sel),
    .io_core_commit_uops_0_ctrl_op_fcn(lsu_io_core_commit_uops_0_ctrl_op_fcn),
    .io_core_commit_uops_0_ctrl_fcn_dw(lsu_io_core_commit_uops_0_ctrl_fcn_dw),
    .io_core_commit_uops_0_ctrl_csr_cmd(lsu_io_core_commit_uops_0_ctrl_csr_cmd),
    .io_core_commit_uops_0_ctrl_is_load(lsu_io_core_commit_uops_0_ctrl_is_load),
    .io_core_commit_uops_0_ctrl_is_sta(lsu_io_core_commit_uops_0_ctrl_is_sta),
    .io_core_commit_uops_0_ctrl_is_std(lsu_io_core_commit_uops_0_ctrl_is_std),
    .io_core_commit_uops_0_ctrl_op3_sel(lsu_io_core_commit_uops_0_ctrl_op3_sel),
    .io_core_commit_uops_0_iw_state(lsu_io_core_commit_uops_0_iw_state),
    .io_core_commit_uops_0_iw_p1_poisoned(lsu_io_core_commit_uops_0_iw_p1_poisoned),
    .io_core_commit_uops_0_iw_p2_poisoned(lsu_io_core_commit_uops_0_iw_p2_poisoned),
    .io_core_commit_uops_0_is_br(lsu_io_core_commit_uops_0_is_br),
    .io_core_commit_uops_0_is_jalr(lsu_io_core_commit_uops_0_is_jalr),
    .io_core_commit_uops_0_is_jal(lsu_io_core_commit_uops_0_is_jal),
    .io_core_commit_uops_0_is_sfb(lsu_io_core_commit_uops_0_is_sfb),
    .io_core_commit_uops_0_br_mask(lsu_io_core_commit_uops_0_br_mask),
    .io_core_commit_uops_0_br_tag(lsu_io_core_commit_uops_0_br_tag),
    .io_core_commit_uops_0_ftq_idx(lsu_io_core_commit_uops_0_ftq_idx),
    .io_core_commit_uops_0_edge_inst(lsu_io_core_commit_uops_0_edge_inst),
    .io_core_commit_uops_0_pc_lob(lsu_io_core_commit_uops_0_pc_lob),
    .io_core_commit_uops_0_taken(lsu_io_core_commit_uops_0_taken),
    .io_core_commit_uops_0_imm_packed(lsu_io_core_commit_uops_0_imm_packed),
    .io_core_commit_uops_0_csr_addr(lsu_io_core_commit_uops_0_csr_addr),
    .io_core_commit_uops_0_rob_idx(lsu_io_core_commit_uops_0_rob_idx),
    .io_core_commit_uops_0_ldq_idx(lsu_io_core_commit_uops_0_ldq_idx),
    .io_core_commit_uops_0_stq_idx(lsu_io_core_commit_uops_0_stq_idx),
    .io_core_commit_uops_0_rxq_idx(lsu_io_core_commit_uops_0_rxq_idx),
    .io_core_commit_uops_0_pdst(lsu_io_core_commit_uops_0_pdst),
    .io_core_commit_uops_0_prs1(lsu_io_core_commit_uops_0_prs1),
    .io_core_commit_uops_0_prs2(lsu_io_core_commit_uops_0_prs2),
    .io_core_commit_uops_0_prs3(lsu_io_core_commit_uops_0_prs3),
    .io_core_commit_uops_0_ppred(lsu_io_core_commit_uops_0_ppred),
    .io_core_commit_uops_0_prs1_busy(lsu_io_core_commit_uops_0_prs1_busy),
    .io_core_commit_uops_0_prs2_busy(lsu_io_core_commit_uops_0_prs2_busy),
    .io_core_commit_uops_0_prs3_busy(lsu_io_core_commit_uops_0_prs3_busy),
    .io_core_commit_uops_0_ppred_busy(lsu_io_core_commit_uops_0_ppred_busy),
    .io_core_commit_uops_0_stale_pdst(lsu_io_core_commit_uops_0_stale_pdst),
    .io_core_commit_uops_0_exception(lsu_io_core_commit_uops_0_exception),
    .io_core_commit_uops_0_exc_cause(lsu_io_core_commit_uops_0_exc_cause),
    .io_core_commit_uops_0_bypassable(lsu_io_core_commit_uops_0_bypassable),
    .io_core_commit_uops_0_mem_cmd(lsu_io_core_commit_uops_0_mem_cmd),
    .io_core_commit_uops_0_mem_size(lsu_io_core_commit_uops_0_mem_size),
    .io_core_commit_uops_0_mem_signed(lsu_io_core_commit_uops_0_mem_signed),
    .io_core_commit_uops_0_is_fence(lsu_io_core_commit_uops_0_is_fence),
    .io_core_commit_uops_0_is_fencei(lsu_io_core_commit_uops_0_is_fencei),
    .io_core_commit_uops_0_is_amo(lsu_io_core_commit_uops_0_is_amo),
    .io_core_commit_uops_0_uses_ldq(lsu_io_core_commit_uops_0_uses_ldq),
    .io_core_commit_uops_0_uses_stq(lsu_io_core_commit_uops_0_uses_stq),
    .io_core_commit_uops_0_is_sys_pc2epc(lsu_io_core_commit_uops_0_is_sys_pc2epc),
    .io_core_commit_uops_0_is_unique(lsu_io_core_commit_uops_0_is_unique),
    .io_core_commit_uops_0_flush_on_commit(lsu_io_core_commit_uops_0_flush_on_commit),
    .io_core_commit_uops_0_ldst_is_rs1(lsu_io_core_commit_uops_0_ldst_is_rs1),
    .io_core_commit_uops_0_ldst(lsu_io_core_commit_uops_0_ldst),
    .io_core_commit_uops_0_lrs1(lsu_io_core_commit_uops_0_lrs1),
    .io_core_commit_uops_0_lrs2(lsu_io_core_commit_uops_0_lrs2),
    .io_core_commit_uops_0_lrs3(lsu_io_core_commit_uops_0_lrs3),
    .io_core_commit_uops_0_ldst_val(lsu_io_core_commit_uops_0_ldst_val),
    .io_core_commit_uops_0_dst_rtype(lsu_io_core_commit_uops_0_dst_rtype),
    .io_core_commit_uops_0_lrs1_rtype(lsu_io_core_commit_uops_0_lrs1_rtype),
    .io_core_commit_uops_0_lrs2_rtype(lsu_io_core_commit_uops_0_lrs2_rtype),
    .io_core_commit_uops_0_frs3_en(lsu_io_core_commit_uops_0_frs3_en),
    .io_core_commit_uops_0_fp_val(lsu_io_core_commit_uops_0_fp_val),
    .io_core_commit_uops_0_fp_single(lsu_io_core_commit_uops_0_fp_single),
    .io_core_commit_uops_0_xcpt_pf_if(lsu_io_core_commit_uops_0_xcpt_pf_if),
    .io_core_commit_uops_0_xcpt_ae_if(lsu_io_core_commit_uops_0_xcpt_ae_if),
    .io_core_commit_uops_0_xcpt_ma_if(lsu_io_core_commit_uops_0_xcpt_ma_if),
    .io_core_commit_uops_0_bp_debug_if(lsu_io_core_commit_uops_0_bp_debug_if),
    .io_core_commit_uops_0_bp_xcpt_if(lsu_io_core_commit_uops_0_bp_xcpt_if),
    .io_core_commit_uops_0_debug_fsrc(lsu_io_core_commit_uops_0_debug_fsrc),
    .io_core_commit_uops_0_debug_tsrc(lsu_io_core_commit_uops_0_debug_tsrc),
    .io_core_commit_uops_1_switch(lsu_io_core_commit_uops_1_switch),
    .io_core_commit_uops_1_switch_off(lsu_io_core_commit_uops_1_switch_off),
    .io_core_commit_uops_1_is_unicore(lsu_io_core_commit_uops_1_is_unicore),
    .io_core_commit_uops_1_shift(lsu_io_core_commit_uops_1_shift),
    .io_core_commit_uops_1_lrs3_rtype(lsu_io_core_commit_uops_1_lrs3_rtype),
    .io_core_commit_uops_1_rflag(lsu_io_core_commit_uops_1_rflag),
    .io_core_commit_uops_1_wflag(lsu_io_core_commit_uops_1_wflag),
    .io_core_commit_uops_1_prflag(lsu_io_core_commit_uops_1_prflag),
    .io_core_commit_uops_1_pwflag(lsu_io_core_commit_uops_1_pwflag),
    .io_core_commit_uops_1_pflag_busy(lsu_io_core_commit_uops_1_pflag_busy),
    .io_core_commit_uops_1_stale_pflag(lsu_io_core_commit_uops_1_stale_pflag),
    .io_core_commit_uops_1_op1_sel(lsu_io_core_commit_uops_1_op1_sel),
    .io_core_commit_uops_1_op2_sel(lsu_io_core_commit_uops_1_op2_sel),
    .io_core_commit_uops_1_split_num(lsu_io_core_commit_uops_1_split_num),
    .io_core_commit_uops_1_self_index(lsu_io_core_commit_uops_1_self_index),
    .io_core_commit_uops_1_rob_inst_idx(lsu_io_core_commit_uops_1_rob_inst_idx),
    .io_core_commit_uops_1_address_num(lsu_io_core_commit_uops_1_address_num),
    .io_core_commit_uops_1_uopc(lsu_io_core_commit_uops_1_uopc),
    .io_core_commit_uops_1_inst(lsu_io_core_commit_uops_1_inst),
    .io_core_commit_uops_1_debug_inst(lsu_io_core_commit_uops_1_debug_inst),
    .io_core_commit_uops_1_is_rvc(lsu_io_core_commit_uops_1_is_rvc),
    .io_core_commit_uops_1_debug_pc(lsu_io_core_commit_uops_1_debug_pc),
    .io_core_commit_uops_1_iq_type(lsu_io_core_commit_uops_1_iq_type),
    .io_core_commit_uops_1_fu_code(lsu_io_core_commit_uops_1_fu_code),
    .io_core_commit_uops_1_ctrl_br_type(lsu_io_core_commit_uops_1_ctrl_br_type),
    .io_core_commit_uops_1_ctrl_op1_sel(lsu_io_core_commit_uops_1_ctrl_op1_sel),
    .io_core_commit_uops_1_ctrl_op2_sel(lsu_io_core_commit_uops_1_ctrl_op2_sel),
    .io_core_commit_uops_1_ctrl_imm_sel(lsu_io_core_commit_uops_1_ctrl_imm_sel),
    .io_core_commit_uops_1_ctrl_op_fcn(lsu_io_core_commit_uops_1_ctrl_op_fcn),
    .io_core_commit_uops_1_ctrl_fcn_dw(lsu_io_core_commit_uops_1_ctrl_fcn_dw),
    .io_core_commit_uops_1_ctrl_csr_cmd(lsu_io_core_commit_uops_1_ctrl_csr_cmd),
    .io_core_commit_uops_1_ctrl_is_load(lsu_io_core_commit_uops_1_ctrl_is_load),
    .io_core_commit_uops_1_ctrl_is_sta(lsu_io_core_commit_uops_1_ctrl_is_sta),
    .io_core_commit_uops_1_ctrl_is_std(lsu_io_core_commit_uops_1_ctrl_is_std),
    .io_core_commit_uops_1_ctrl_op3_sel(lsu_io_core_commit_uops_1_ctrl_op3_sel),
    .io_core_commit_uops_1_iw_state(lsu_io_core_commit_uops_1_iw_state),
    .io_core_commit_uops_1_iw_p1_poisoned(lsu_io_core_commit_uops_1_iw_p1_poisoned),
    .io_core_commit_uops_1_iw_p2_poisoned(lsu_io_core_commit_uops_1_iw_p2_poisoned),
    .io_core_commit_uops_1_is_br(lsu_io_core_commit_uops_1_is_br),
    .io_core_commit_uops_1_is_jalr(lsu_io_core_commit_uops_1_is_jalr),
    .io_core_commit_uops_1_is_jal(lsu_io_core_commit_uops_1_is_jal),
    .io_core_commit_uops_1_is_sfb(lsu_io_core_commit_uops_1_is_sfb),
    .io_core_commit_uops_1_br_mask(lsu_io_core_commit_uops_1_br_mask),
    .io_core_commit_uops_1_br_tag(lsu_io_core_commit_uops_1_br_tag),
    .io_core_commit_uops_1_ftq_idx(lsu_io_core_commit_uops_1_ftq_idx),
    .io_core_commit_uops_1_edge_inst(lsu_io_core_commit_uops_1_edge_inst),
    .io_core_commit_uops_1_pc_lob(lsu_io_core_commit_uops_1_pc_lob),
    .io_core_commit_uops_1_taken(lsu_io_core_commit_uops_1_taken),
    .io_core_commit_uops_1_imm_packed(lsu_io_core_commit_uops_1_imm_packed),
    .io_core_commit_uops_1_csr_addr(lsu_io_core_commit_uops_1_csr_addr),
    .io_core_commit_uops_1_rob_idx(lsu_io_core_commit_uops_1_rob_idx),
    .io_core_commit_uops_1_ldq_idx(lsu_io_core_commit_uops_1_ldq_idx),
    .io_core_commit_uops_1_stq_idx(lsu_io_core_commit_uops_1_stq_idx),
    .io_core_commit_uops_1_rxq_idx(lsu_io_core_commit_uops_1_rxq_idx),
    .io_core_commit_uops_1_pdst(lsu_io_core_commit_uops_1_pdst),
    .io_core_commit_uops_1_prs1(lsu_io_core_commit_uops_1_prs1),
    .io_core_commit_uops_1_prs2(lsu_io_core_commit_uops_1_prs2),
    .io_core_commit_uops_1_prs3(lsu_io_core_commit_uops_1_prs3),
    .io_core_commit_uops_1_ppred(lsu_io_core_commit_uops_1_ppred),
    .io_core_commit_uops_1_prs1_busy(lsu_io_core_commit_uops_1_prs1_busy),
    .io_core_commit_uops_1_prs2_busy(lsu_io_core_commit_uops_1_prs2_busy),
    .io_core_commit_uops_1_prs3_busy(lsu_io_core_commit_uops_1_prs3_busy),
    .io_core_commit_uops_1_ppred_busy(lsu_io_core_commit_uops_1_ppred_busy),
    .io_core_commit_uops_1_stale_pdst(lsu_io_core_commit_uops_1_stale_pdst),
    .io_core_commit_uops_1_exception(lsu_io_core_commit_uops_1_exception),
    .io_core_commit_uops_1_exc_cause(lsu_io_core_commit_uops_1_exc_cause),
    .io_core_commit_uops_1_bypassable(lsu_io_core_commit_uops_1_bypassable),
    .io_core_commit_uops_1_mem_cmd(lsu_io_core_commit_uops_1_mem_cmd),
    .io_core_commit_uops_1_mem_size(lsu_io_core_commit_uops_1_mem_size),
    .io_core_commit_uops_1_mem_signed(lsu_io_core_commit_uops_1_mem_signed),
    .io_core_commit_uops_1_is_fence(lsu_io_core_commit_uops_1_is_fence),
    .io_core_commit_uops_1_is_fencei(lsu_io_core_commit_uops_1_is_fencei),
    .io_core_commit_uops_1_is_amo(lsu_io_core_commit_uops_1_is_amo),
    .io_core_commit_uops_1_uses_ldq(lsu_io_core_commit_uops_1_uses_ldq),
    .io_core_commit_uops_1_uses_stq(lsu_io_core_commit_uops_1_uses_stq),
    .io_core_commit_uops_1_is_sys_pc2epc(lsu_io_core_commit_uops_1_is_sys_pc2epc),
    .io_core_commit_uops_1_is_unique(lsu_io_core_commit_uops_1_is_unique),
    .io_core_commit_uops_1_flush_on_commit(lsu_io_core_commit_uops_1_flush_on_commit),
    .io_core_commit_uops_1_ldst_is_rs1(lsu_io_core_commit_uops_1_ldst_is_rs1),
    .io_core_commit_uops_1_ldst(lsu_io_core_commit_uops_1_ldst),
    .io_core_commit_uops_1_lrs1(lsu_io_core_commit_uops_1_lrs1),
    .io_core_commit_uops_1_lrs2(lsu_io_core_commit_uops_1_lrs2),
    .io_core_commit_uops_1_lrs3(lsu_io_core_commit_uops_1_lrs3),
    .io_core_commit_uops_1_ldst_val(lsu_io_core_commit_uops_1_ldst_val),
    .io_core_commit_uops_1_dst_rtype(lsu_io_core_commit_uops_1_dst_rtype),
    .io_core_commit_uops_1_lrs1_rtype(lsu_io_core_commit_uops_1_lrs1_rtype),
    .io_core_commit_uops_1_lrs2_rtype(lsu_io_core_commit_uops_1_lrs2_rtype),
    .io_core_commit_uops_1_frs3_en(lsu_io_core_commit_uops_1_frs3_en),
    .io_core_commit_uops_1_fp_val(lsu_io_core_commit_uops_1_fp_val),
    .io_core_commit_uops_1_fp_single(lsu_io_core_commit_uops_1_fp_single),
    .io_core_commit_uops_1_xcpt_pf_if(lsu_io_core_commit_uops_1_xcpt_pf_if),
    .io_core_commit_uops_1_xcpt_ae_if(lsu_io_core_commit_uops_1_xcpt_ae_if),
    .io_core_commit_uops_1_xcpt_ma_if(lsu_io_core_commit_uops_1_xcpt_ma_if),
    .io_core_commit_uops_1_bp_debug_if(lsu_io_core_commit_uops_1_bp_debug_if),
    .io_core_commit_uops_1_bp_xcpt_if(lsu_io_core_commit_uops_1_bp_xcpt_if),
    .io_core_commit_uops_1_debug_fsrc(lsu_io_core_commit_uops_1_debug_fsrc),
    .io_core_commit_uops_1_debug_tsrc(lsu_io_core_commit_uops_1_debug_tsrc),
    .io_core_commit_fflags_valid(lsu_io_core_commit_fflags_valid),
    .io_core_commit_fflags_bits(lsu_io_core_commit_fflags_bits),
    .io_core_commit_fflag_exception_valid(lsu_io_core_commit_fflag_exception_valid),
    .io_core_commit_fflag_exception_bits(lsu_io_core_commit_fflag_exception_bits),
    .io_core_commit_debug_insts_0(lsu_io_core_commit_debug_insts_0),
    .io_core_commit_debug_insts_1(lsu_io_core_commit_debug_insts_1),
    .io_core_commit_rbk_valids_0(lsu_io_core_commit_rbk_valids_0),
    .io_core_commit_rbk_valids_1(lsu_io_core_commit_rbk_valids_1),
    .io_core_commit_rollback(lsu_io_core_commit_rollback),
    .io_core_commit_debug_wdata_0(lsu_io_core_commit_debug_wdata_0),
    .io_core_commit_debug_wdata_1(lsu_io_core_commit_debug_wdata_1),
    .io_core_commit_debug_wflagdata_0(lsu_io_core_commit_debug_wflagdata_0),
    .io_core_commit_debug_wflagdata_1(lsu_io_core_commit_debug_wflagdata_1),
    .io_core_commit_load_at_rob_head(lsu_io_core_commit_load_at_rob_head),
    .io_core_clr_bsy_0_valid(lsu_io_core_clr_bsy_0_valid),
    .io_core_clr_bsy_0_bits(lsu_io_core_clr_bsy_0_bits),
    .io_core_clr_bsy_1_valid(lsu_io_core_clr_bsy_1_valid),
    .io_core_clr_bsy_1_bits(lsu_io_core_clr_bsy_1_bits),
    .io_core_clr_unsafe_0_valid(lsu_io_core_clr_unsafe_0_valid),
    .io_core_clr_unsafe_0_bits(lsu_io_core_clr_unsafe_0_bits),
    .io_core_clr_bsy_first_idx_0(lsu_io_core_clr_bsy_first_idx_0),
    .io_core_clr_bsy_first_idx_1(lsu_io_core_clr_bsy_first_idx_1),
    .io_core_clr_bsy_self_idx_0(lsu_io_core_clr_bsy_self_idx_0),
    .io_core_clr_bsy_self_idx_1(lsu_io_core_clr_bsy_self_idx_1),
    .io_core_fence_dmem(lsu_io_core_fence_dmem),
    .io_core_spec_ld_wakeup_0_valid(lsu_io_core_spec_ld_wakeup_0_valid),
    .io_core_spec_ld_wakeup_0_bits(lsu_io_core_spec_ld_wakeup_0_bits),
    .io_core_ld_miss(lsu_io_core_ld_miss),
    .io_core_brupdate_b1_resolve_mask(lsu_io_core_brupdate_b1_resolve_mask),
    .io_core_brupdate_b1_mispredict_mask(lsu_io_core_brupdate_b1_mispredict_mask),
    .io_core_brupdate_b2_uop_switch(lsu_io_core_brupdate_b2_uop_switch),
    .io_core_brupdate_b2_uop_switch_off(lsu_io_core_brupdate_b2_uop_switch_off),
    .io_core_brupdate_b2_uop_is_unicore(lsu_io_core_brupdate_b2_uop_is_unicore),
    .io_core_brupdate_b2_uop_shift(lsu_io_core_brupdate_b2_uop_shift),
    .io_core_brupdate_b2_uop_lrs3_rtype(lsu_io_core_brupdate_b2_uop_lrs3_rtype),
    .io_core_brupdate_b2_uop_rflag(lsu_io_core_brupdate_b2_uop_rflag),
    .io_core_brupdate_b2_uop_wflag(lsu_io_core_brupdate_b2_uop_wflag),
    .io_core_brupdate_b2_uop_prflag(lsu_io_core_brupdate_b2_uop_prflag),
    .io_core_brupdate_b2_uop_pwflag(lsu_io_core_brupdate_b2_uop_pwflag),
    .io_core_brupdate_b2_uop_pflag_busy(lsu_io_core_brupdate_b2_uop_pflag_busy),
    .io_core_brupdate_b2_uop_stale_pflag(lsu_io_core_brupdate_b2_uop_stale_pflag),
    .io_core_brupdate_b2_uop_op1_sel(lsu_io_core_brupdate_b2_uop_op1_sel),
    .io_core_brupdate_b2_uop_op2_sel(lsu_io_core_brupdate_b2_uop_op2_sel),
    .io_core_brupdate_b2_uop_split_num(lsu_io_core_brupdate_b2_uop_split_num),
    .io_core_brupdate_b2_uop_self_index(lsu_io_core_brupdate_b2_uop_self_index),
    .io_core_brupdate_b2_uop_rob_inst_idx(lsu_io_core_brupdate_b2_uop_rob_inst_idx),
    .io_core_brupdate_b2_uop_address_num(lsu_io_core_brupdate_b2_uop_address_num),
    .io_core_brupdate_b2_uop_uopc(lsu_io_core_brupdate_b2_uop_uopc),
    .io_core_brupdate_b2_uop_inst(lsu_io_core_brupdate_b2_uop_inst),
    .io_core_brupdate_b2_uop_debug_inst(lsu_io_core_brupdate_b2_uop_debug_inst),
    .io_core_brupdate_b2_uop_is_rvc(lsu_io_core_brupdate_b2_uop_is_rvc),
    .io_core_brupdate_b2_uop_debug_pc(lsu_io_core_brupdate_b2_uop_debug_pc),
    .io_core_brupdate_b2_uop_iq_type(lsu_io_core_brupdate_b2_uop_iq_type),
    .io_core_brupdate_b2_uop_fu_code(lsu_io_core_brupdate_b2_uop_fu_code),
    .io_core_brupdate_b2_uop_ctrl_br_type(lsu_io_core_brupdate_b2_uop_ctrl_br_type),
    .io_core_brupdate_b2_uop_ctrl_op1_sel(lsu_io_core_brupdate_b2_uop_ctrl_op1_sel),
    .io_core_brupdate_b2_uop_ctrl_op2_sel(lsu_io_core_brupdate_b2_uop_ctrl_op2_sel),
    .io_core_brupdate_b2_uop_ctrl_imm_sel(lsu_io_core_brupdate_b2_uop_ctrl_imm_sel),
    .io_core_brupdate_b2_uop_ctrl_op_fcn(lsu_io_core_brupdate_b2_uop_ctrl_op_fcn),
    .io_core_brupdate_b2_uop_ctrl_fcn_dw(lsu_io_core_brupdate_b2_uop_ctrl_fcn_dw),
    .io_core_brupdate_b2_uop_ctrl_csr_cmd(lsu_io_core_brupdate_b2_uop_ctrl_csr_cmd),
    .io_core_brupdate_b2_uop_ctrl_is_load(lsu_io_core_brupdate_b2_uop_ctrl_is_load),
    .io_core_brupdate_b2_uop_ctrl_is_sta(lsu_io_core_brupdate_b2_uop_ctrl_is_sta),
    .io_core_brupdate_b2_uop_ctrl_is_std(lsu_io_core_brupdate_b2_uop_ctrl_is_std),
    .io_core_brupdate_b2_uop_ctrl_op3_sel(lsu_io_core_brupdate_b2_uop_ctrl_op3_sel),
    .io_core_brupdate_b2_uop_iw_state(lsu_io_core_brupdate_b2_uop_iw_state),
    .io_core_brupdate_b2_uop_iw_p1_poisoned(lsu_io_core_brupdate_b2_uop_iw_p1_poisoned),
    .io_core_brupdate_b2_uop_iw_p2_poisoned(lsu_io_core_brupdate_b2_uop_iw_p2_poisoned),
    .io_core_brupdate_b2_uop_is_br(lsu_io_core_brupdate_b2_uop_is_br),
    .io_core_brupdate_b2_uop_is_jalr(lsu_io_core_brupdate_b2_uop_is_jalr),
    .io_core_brupdate_b2_uop_is_jal(lsu_io_core_brupdate_b2_uop_is_jal),
    .io_core_brupdate_b2_uop_is_sfb(lsu_io_core_brupdate_b2_uop_is_sfb),
    .io_core_brupdate_b2_uop_br_mask(lsu_io_core_brupdate_b2_uop_br_mask),
    .io_core_brupdate_b2_uop_br_tag(lsu_io_core_brupdate_b2_uop_br_tag),
    .io_core_brupdate_b2_uop_ftq_idx(lsu_io_core_brupdate_b2_uop_ftq_idx),
    .io_core_brupdate_b2_uop_edge_inst(lsu_io_core_brupdate_b2_uop_edge_inst),
    .io_core_brupdate_b2_uop_pc_lob(lsu_io_core_brupdate_b2_uop_pc_lob),
    .io_core_brupdate_b2_uop_taken(lsu_io_core_brupdate_b2_uop_taken),
    .io_core_brupdate_b2_uop_imm_packed(lsu_io_core_brupdate_b2_uop_imm_packed),
    .io_core_brupdate_b2_uop_csr_addr(lsu_io_core_brupdate_b2_uop_csr_addr),
    .io_core_brupdate_b2_uop_rob_idx(lsu_io_core_brupdate_b2_uop_rob_idx),
    .io_core_brupdate_b2_uop_ldq_idx(lsu_io_core_brupdate_b2_uop_ldq_idx),
    .io_core_brupdate_b2_uop_stq_idx(lsu_io_core_brupdate_b2_uop_stq_idx),
    .io_core_brupdate_b2_uop_rxq_idx(lsu_io_core_brupdate_b2_uop_rxq_idx),
    .io_core_brupdate_b2_uop_pdst(lsu_io_core_brupdate_b2_uop_pdst),
    .io_core_brupdate_b2_uop_prs1(lsu_io_core_brupdate_b2_uop_prs1),
    .io_core_brupdate_b2_uop_prs2(lsu_io_core_brupdate_b2_uop_prs2),
    .io_core_brupdate_b2_uop_prs3(lsu_io_core_brupdate_b2_uop_prs3),
    .io_core_brupdate_b2_uop_ppred(lsu_io_core_brupdate_b2_uop_ppred),
    .io_core_brupdate_b2_uop_prs1_busy(lsu_io_core_brupdate_b2_uop_prs1_busy),
    .io_core_brupdate_b2_uop_prs2_busy(lsu_io_core_brupdate_b2_uop_prs2_busy),
    .io_core_brupdate_b2_uop_prs3_busy(lsu_io_core_brupdate_b2_uop_prs3_busy),
    .io_core_brupdate_b2_uop_ppred_busy(lsu_io_core_brupdate_b2_uop_ppred_busy),
    .io_core_brupdate_b2_uop_stale_pdst(lsu_io_core_brupdate_b2_uop_stale_pdst),
    .io_core_brupdate_b2_uop_exception(lsu_io_core_brupdate_b2_uop_exception),
    .io_core_brupdate_b2_uop_exc_cause(lsu_io_core_brupdate_b2_uop_exc_cause),
    .io_core_brupdate_b2_uop_bypassable(lsu_io_core_brupdate_b2_uop_bypassable),
    .io_core_brupdate_b2_uop_mem_cmd(lsu_io_core_brupdate_b2_uop_mem_cmd),
    .io_core_brupdate_b2_uop_mem_size(lsu_io_core_brupdate_b2_uop_mem_size),
    .io_core_brupdate_b2_uop_mem_signed(lsu_io_core_brupdate_b2_uop_mem_signed),
    .io_core_brupdate_b2_uop_is_fence(lsu_io_core_brupdate_b2_uop_is_fence),
    .io_core_brupdate_b2_uop_is_fencei(lsu_io_core_brupdate_b2_uop_is_fencei),
    .io_core_brupdate_b2_uop_is_amo(lsu_io_core_brupdate_b2_uop_is_amo),
    .io_core_brupdate_b2_uop_uses_ldq(lsu_io_core_brupdate_b2_uop_uses_ldq),
    .io_core_brupdate_b2_uop_uses_stq(lsu_io_core_brupdate_b2_uop_uses_stq),
    .io_core_brupdate_b2_uop_is_sys_pc2epc(lsu_io_core_brupdate_b2_uop_is_sys_pc2epc),
    .io_core_brupdate_b2_uop_is_unique(lsu_io_core_brupdate_b2_uop_is_unique),
    .io_core_brupdate_b2_uop_flush_on_commit(lsu_io_core_brupdate_b2_uop_flush_on_commit),
    .io_core_brupdate_b2_uop_ldst_is_rs1(lsu_io_core_brupdate_b2_uop_ldst_is_rs1),
    .io_core_brupdate_b2_uop_ldst(lsu_io_core_brupdate_b2_uop_ldst),
    .io_core_brupdate_b2_uop_lrs1(lsu_io_core_brupdate_b2_uop_lrs1),
    .io_core_brupdate_b2_uop_lrs2(lsu_io_core_brupdate_b2_uop_lrs2),
    .io_core_brupdate_b2_uop_lrs3(lsu_io_core_brupdate_b2_uop_lrs3),
    .io_core_brupdate_b2_uop_ldst_val(lsu_io_core_brupdate_b2_uop_ldst_val),
    .io_core_brupdate_b2_uop_dst_rtype(lsu_io_core_brupdate_b2_uop_dst_rtype),
    .io_core_brupdate_b2_uop_lrs1_rtype(lsu_io_core_brupdate_b2_uop_lrs1_rtype),
    .io_core_brupdate_b2_uop_lrs2_rtype(lsu_io_core_brupdate_b2_uop_lrs2_rtype),
    .io_core_brupdate_b2_uop_frs3_en(lsu_io_core_brupdate_b2_uop_frs3_en),
    .io_core_brupdate_b2_uop_fp_val(lsu_io_core_brupdate_b2_uop_fp_val),
    .io_core_brupdate_b2_uop_fp_single(lsu_io_core_brupdate_b2_uop_fp_single),
    .io_core_brupdate_b2_uop_xcpt_pf_if(lsu_io_core_brupdate_b2_uop_xcpt_pf_if),
    .io_core_brupdate_b2_uop_xcpt_ae_if(lsu_io_core_brupdate_b2_uop_xcpt_ae_if),
    .io_core_brupdate_b2_uop_xcpt_ma_if(lsu_io_core_brupdate_b2_uop_xcpt_ma_if),
    .io_core_brupdate_b2_uop_bp_debug_if(lsu_io_core_brupdate_b2_uop_bp_debug_if),
    .io_core_brupdate_b2_uop_bp_xcpt_if(lsu_io_core_brupdate_b2_uop_bp_xcpt_if),
    .io_core_brupdate_b2_uop_debug_fsrc(lsu_io_core_brupdate_b2_uop_debug_fsrc),
    .io_core_brupdate_b2_uop_debug_tsrc(lsu_io_core_brupdate_b2_uop_debug_tsrc),
    .io_core_brupdate_b2_valid(lsu_io_core_brupdate_b2_valid),
    .io_core_brupdate_b2_mispredict(lsu_io_core_brupdate_b2_mispredict),
    .io_core_brupdate_b2_taken(lsu_io_core_brupdate_b2_taken),
    .io_core_brupdate_b2_cfi_type(lsu_io_core_brupdate_b2_cfi_type),
    .io_core_brupdate_b2_pc_sel(lsu_io_core_brupdate_b2_pc_sel),
    .io_core_brupdate_b2_jalr_target(lsu_io_core_brupdate_b2_jalr_target),
    .io_core_brupdate_b2_target_offset(lsu_io_core_brupdate_b2_target_offset),
    .io_core_rob_pnr_idx(lsu_io_core_rob_pnr_idx),
    .io_core_rob_head_idx(lsu_io_core_rob_head_idx),
    .io_core_exception(lsu_io_core_exception),
    .io_core_fencei_rdy(lsu_io_core_fencei_rdy),
    .io_core_lxcpt_valid(lsu_io_core_lxcpt_valid),
    .io_core_lxcpt_bits_uop_switch(lsu_io_core_lxcpt_bits_uop_switch),
    .io_core_lxcpt_bits_uop_switch_off(lsu_io_core_lxcpt_bits_uop_switch_off),
    .io_core_lxcpt_bits_uop_is_unicore(lsu_io_core_lxcpt_bits_uop_is_unicore),
    .io_core_lxcpt_bits_uop_shift(lsu_io_core_lxcpt_bits_uop_shift),
    .io_core_lxcpt_bits_uop_lrs3_rtype(lsu_io_core_lxcpt_bits_uop_lrs3_rtype),
    .io_core_lxcpt_bits_uop_rflag(lsu_io_core_lxcpt_bits_uop_rflag),
    .io_core_lxcpt_bits_uop_wflag(lsu_io_core_lxcpt_bits_uop_wflag),
    .io_core_lxcpt_bits_uop_prflag(lsu_io_core_lxcpt_bits_uop_prflag),
    .io_core_lxcpt_bits_uop_pwflag(lsu_io_core_lxcpt_bits_uop_pwflag),
    .io_core_lxcpt_bits_uop_pflag_busy(lsu_io_core_lxcpt_bits_uop_pflag_busy),
    .io_core_lxcpt_bits_uop_stale_pflag(lsu_io_core_lxcpt_bits_uop_stale_pflag),
    .io_core_lxcpt_bits_uop_op1_sel(lsu_io_core_lxcpt_bits_uop_op1_sel),
    .io_core_lxcpt_bits_uop_op2_sel(lsu_io_core_lxcpt_bits_uop_op2_sel),
    .io_core_lxcpt_bits_uop_split_num(lsu_io_core_lxcpt_bits_uop_split_num),
    .io_core_lxcpt_bits_uop_self_index(lsu_io_core_lxcpt_bits_uop_self_index),
    .io_core_lxcpt_bits_uop_rob_inst_idx(lsu_io_core_lxcpt_bits_uop_rob_inst_idx),
    .io_core_lxcpt_bits_uop_address_num(lsu_io_core_lxcpt_bits_uop_address_num),
    .io_core_lxcpt_bits_uop_uopc(lsu_io_core_lxcpt_bits_uop_uopc),
    .io_core_lxcpt_bits_uop_inst(lsu_io_core_lxcpt_bits_uop_inst),
    .io_core_lxcpt_bits_uop_debug_inst(lsu_io_core_lxcpt_bits_uop_debug_inst),
    .io_core_lxcpt_bits_uop_is_rvc(lsu_io_core_lxcpt_bits_uop_is_rvc),
    .io_core_lxcpt_bits_uop_debug_pc(lsu_io_core_lxcpt_bits_uop_debug_pc),
    .io_core_lxcpt_bits_uop_iq_type(lsu_io_core_lxcpt_bits_uop_iq_type),
    .io_core_lxcpt_bits_uop_fu_code(lsu_io_core_lxcpt_bits_uop_fu_code),
    .io_core_lxcpt_bits_uop_ctrl_br_type(lsu_io_core_lxcpt_bits_uop_ctrl_br_type),
    .io_core_lxcpt_bits_uop_ctrl_op1_sel(lsu_io_core_lxcpt_bits_uop_ctrl_op1_sel),
    .io_core_lxcpt_bits_uop_ctrl_op2_sel(lsu_io_core_lxcpt_bits_uop_ctrl_op2_sel),
    .io_core_lxcpt_bits_uop_ctrl_imm_sel(lsu_io_core_lxcpt_bits_uop_ctrl_imm_sel),
    .io_core_lxcpt_bits_uop_ctrl_op_fcn(lsu_io_core_lxcpt_bits_uop_ctrl_op_fcn),
    .io_core_lxcpt_bits_uop_ctrl_fcn_dw(lsu_io_core_lxcpt_bits_uop_ctrl_fcn_dw),
    .io_core_lxcpt_bits_uop_ctrl_csr_cmd(lsu_io_core_lxcpt_bits_uop_ctrl_csr_cmd),
    .io_core_lxcpt_bits_uop_ctrl_is_load(lsu_io_core_lxcpt_bits_uop_ctrl_is_load),
    .io_core_lxcpt_bits_uop_ctrl_is_sta(lsu_io_core_lxcpt_bits_uop_ctrl_is_sta),
    .io_core_lxcpt_bits_uop_ctrl_is_std(lsu_io_core_lxcpt_bits_uop_ctrl_is_std),
    .io_core_lxcpt_bits_uop_ctrl_op3_sel(lsu_io_core_lxcpt_bits_uop_ctrl_op3_sel),
    .io_core_lxcpt_bits_uop_iw_state(lsu_io_core_lxcpt_bits_uop_iw_state),
    .io_core_lxcpt_bits_uop_iw_p1_poisoned(lsu_io_core_lxcpt_bits_uop_iw_p1_poisoned),
    .io_core_lxcpt_bits_uop_iw_p2_poisoned(lsu_io_core_lxcpt_bits_uop_iw_p2_poisoned),
    .io_core_lxcpt_bits_uop_is_br(lsu_io_core_lxcpt_bits_uop_is_br),
    .io_core_lxcpt_bits_uop_is_jalr(lsu_io_core_lxcpt_bits_uop_is_jalr),
    .io_core_lxcpt_bits_uop_is_jal(lsu_io_core_lxcpt_bits_uop_is_jal),
    .io_core_lxcpt_bits_uop_is_sfb(lsu_io_core_lxcpt_bits_uop_is_sfb),
    .io_core_lxcpt_bits_uop_br_mask(lsu_io_core_lxcpt_bits_uop_br_mask),
    .io_core_lxcpt_bits_uop_br_tag(lsu_io_core_lxcpt_bits_uop_br_tag),
    .io_core_lxcpt_bits_uop_ftq_idx(lsu_io_core_lxcpt_bits_uop_ftq_idx),
    .io_core_lxcpt_bits_uop_edge_inst(lsu_io_core_lxcpt_bits_uop_edge_inst),
    .io_core_lxcpt_bits_uop_pc_lob(lsu_io_core_lxcpt_bits_uop_pc_lob),
    .io_core_lxcpt_bits_uop_taken(lsu_io_core_lxcpt_bits_uop_taken),
    .io_core_lxcpt_bits_uop_imm_packed(lsu_io_core_lxcpt_bits_uop_imm_packed),
    .io_core_lxcpt_bits_uop_csr_addr(lsu_io_core_lxcpt_bits_uop_csr_addr),
    .io_core_lxcpt_bits_uop_rob_idx(lsu_io_core_lxcpt_bits_uop_rob_idx),
    .io_core_lxcpt_bits_uop_ldq_idx(lsu_io_core_lxcpt_bits_uop_ldq_idx),
    .io_core_lxcpt_bits_uop_stq_idx(lsu_io_core_lxcpt_bits_uop_stq_idx),
    .io_core_lxcpt_bits_uop_rxq_idx(lsu_io_core_lxcpt_bits_uop_rxq_idx),
    .io_core_lxcpt_bits_uop_pdst(lsu_io_core_lxcpt_bits_uop_pdst),
    .io_core_lxcpt_bits_uop_prs1(lsu_io_core_lxcpt_bits_uop_prs1),
    .io_core_lxcpt_bits_uop_prs2(lsu_io_core_lxcpt_bits_uop_prs2),
    .io_core_lxcpt_bits_uop_prs3(lsu_io_core_lxcpt_bits_uop_prs3),
    .io_core_lxcpt_bits_uop_ppred(lsu_io_core_lxcpt_bits_uop_ppred),
    .io_core_lxcpt_bits_uop_prs1_busy(lsu_io_core_lxcpt_bits_uop_prs1_busy),
    .io_core_lxcpt_bits_uop_prs2_busy(lsu_io_core_lxcpt_bits_uop_prs2_busy),
    .io_core_lxcpt_bits_uop_prs3_busy(lsu_io_core_lxcpt_bits_uop_prs3_busy),
    .io_core_lxcpt_bits_uop_ppred_busy(lsu_io_core_lxcpt_bits_uop_ppred_busy),
    .io_core_lxcpt_bits_uop_stale_pdst(lsu_io_core_lxcpt_bits_uop_stale_pdst),
    .io_core_lxcpt_bits_uop_exception(lsu_io_core_lxcpt_bits_uop_exception),
    .io_core_lxcpt_bits_uop_exc_cause(lsu_io_core_lxcpt_bits_uop_exc_cause),
    .io_core_lxcpt_bits_uop_bypassable(lsu_io_core_lxcpt_bits_uop_bypassable),
    .io_core_lxcpt_bits_uop_mem_cmd(lsu_io_core_lxcpt_bits_uop_mem_cmd),
    .io_core_lxcpt_bits_uop_mem_size(lsu_io_core_lxcpt_bits_uop_mem_size),
    .io_core_lxcpt_bits_uop_mem_signed(lsu_io_core_lxcpt_bits_uop_mem_signed),
    .io_core_lxcpt_bits_uop_is_fence(lsu_io_core_lxcpt_bits_uop_is_fence),
    .io_core_lxcpt_bits_uop_is_fencei(lsu_io_core_lxcpt_bits_uop_is_fencei),
    .io_core_lxcpt_bits_uop_is_amo(lsu_io_core_lxcpt_bits_uop_is_amo),
    .io_core_lxcpt_bits_uop_uses_ldq(lsu_io_core_lxcpt_bits_uop_uses_ldq),
    .io_core_lxcpt_bits_uop_uses_stq(lsu_io_core_lxcpt_bits_uop_uses_stq),
    .io_core_lxcpt_bits_uop_is_sys_pc2epc(lsu_io_core_lxcpt_bits_uop_is_sys_pc2epc),
    .io_core_lxcpt_bits_uop_is_unique(lsu_io_core_lxcpt_bits_uop_is_unique),
    .io_core_lxcpt_bits_uop_flush_on_commit(lsu_io_core_lxcpt_bits_uop_flush_on_commit),
    .io_core_lxcpt_bits_uop_ldst_is_rs1(lsu_io_core_lxcpt_bits_uop_ldst_is_rs1),
    .io_core_lxcpt_bits_uop_ldst(lsu_io_core_lxcpt_bits_uop_ldst),
    .io_core_lxcpt_bits_uop_lrs1(lsu_io_core_lxcpt_bits_uop_lrs1),
    .io_core_lxcpt_bits_uop_lrs2(lsu_io_core_lxcpt_bits_uop_lrs2),
    .io_core_lxcpt_bits_uop_lrs3(lsu_io_core_lxcpt_bits_uop_lrs3),
    .io_core_lxcpt_bits_uop_ldst_val(lsu_io_core_lxcpt_bits_uop_ldst_val),
    .io_core_lxcpt_bits_uop_dst_rtype(lsu_io_core_lxcpt_bits_uop_dst_rtype),
    .io_core_lxcpt_bits_uop_lrs1_rtype(lsu_io_core_lxcpt_bits_uop_lrs1_rtype),
    .io_core_lxcpt_bits_uop_lrs2_rtype(lsu_io_core_lxcpt_bits_uop_lrs2_rtype),
    .io_core_lxcpt_bits_uop_frs3_en(lsu_io_core_lxcpt_bits_uop_frs3_en),
    .io_core_lxcpt_bits_uop_fp_val(lsu_io_core_lxcpt_bits_uop_fp_val),
    .io_core_lxcpt_bits_uop_fp_single(lsu_io_core_lxcpt_bits_uop_fp_single),
    .io_core_lxcpt_bits_uop_xcpt_pf_if(lsu_io_core_lxcpt_bits_uop_xcpt_pf_if),
    .io_core_lxcpt_bits_uop_xcpt_ae_if(lsu_io_core_lxcpt_bits_uop_xcpt_ae_if),
    .io_core_lxcpt_bits_uop_xcpt_ma_if(lsu_io_core_lxcpt_bits_uop_xcpt_ma_if),
    .io_core_lxcpt_bits_uop_bp_debug_if(lsu_io_core_lxcpt_bits_uop_bp_debug_if),
    .io_core_lxcpt_bits_uop_bp_xcpt_if(lsu_io_core_lxcpt_bits_uop_bp_xcpt_if),
    .io_core_lxcpt_bits_uop_debug_fsrc(lsu_io_core_lxcpt_bits_uop_debug_fsrc),
    .io_core_lxcpt_bits_uop_debug_tsrc(lsu_io_core_lxcpt_bits_uop_debug_tsrc),
    .io_core_lxcpt_bits_cause(lsu_io_core_lxcpt_bits_cause),
    .io_core_lxcpt_bits_badvaddr(lsu_io_core_lxcpt_bits_badvaddr),
    .io_core_tsc_reg(lsu_io_core_tsc_reg),
    .io_core_perf_acquire(lsu_io_core_perf_acquire),
    .io_core_perf_release(lsu_io_core_perf_release),
    .io_core_perf_tlbMiss(lsu_io_core_perf_tlbMiss),
    .io_dmem_req_ready(lsu_io_dmem_req_ready),
    .io_dmem_req_valid(lsu_io_dmem_req_valid),
    .io_dmem_req_bits_0_valid(lsu_io_dmem_req_bits_0_valid),
    .io_dmem_req_bits_0_bits_uop_switch(lsu_io_dmem_req_bits_0_bits_uop_switch),
    .io_dmem_req_bits_0_bits_uop_switch_off(lsu_io_dmem_req_bits_0_bits_uop_switch_off),
    .io_dmem_req_bits_0_bits_uop_is_unicore(lsu_io_dmem_req_bits_0_bits_uop_is_unicore),
    .io_dmem_req_bits_0_bits_uop_shift(lsu_io_dmem_req_bits_0_bits_uop_shift),
    .io_dmem_req_bits_0_bits_uop_lrs3_rtype(lsu_io_dmem_req_bits_0_bits_uop_lrs3_rtype),
    .io_dmem_req_bits_0_bits_uop_rflag(lsu_io_dmem_req_bits_0_bits_uop_rflag),
    .io_dmem_req_bits_0_bits_uop_wflag(lsu_io_dmem_req_bits_0_bits_uop_wflag),
    .io_dmem_req_bits_0_bits_uop_prflag(lsu_io_dmem_req_bits_0_bits_uop_prflag),
    .io_dmem_req_bits_0_bits_uop_pwflag(lsu_io_dmem_req_bits_0_bits_uop_pwflag),
    .io_dmem_req_bits_0_bits_uop_pflag_busy(lsu_io_dmem_req_bits_0_bits_uop_pflag_busy),
    .io_dmem_req_bits_0_bits_uop_stale_pflag(lsu_io_dmem_req_bits_0_bits_uop_stale_pflag),
    .io_dmem_req_bits_0_bits_uop_op1_sel(lsu_io_dmem_req_bits_0_bits_uop_op1_sel),
    .io_dmem_req_bits_0_bits_uop_op2_sel(lsu_io_dmem_req_bits_0_bits_uop_op2_sel),
    .io_dmem_req_bits_0_bits_uop_split_num(lsu_io_dmem_req_bits_0_bits_uop_split_num),
    .io_dmem_req_bits_0_bits_uop_self_index(lsu_io_dmem_req_bits_0_bits_uop_self_index),
    .io_dmem_req_bits_0_bits_uop_rob_inst_idx(lsu_io_dmem_req_bits_0_bits_uop_rob_inst_idx),
    .io_dmem_req_bits_0_bits_uop_address_num(lsu_io_dmem_req_bits_0_bits_uop_address_num),
    .io_dmem_req_bits_0_bits_uop_uopc(lsu_io_dmem_req_bits_0_bits_uop_uopc),
    .io_dmem_req_bits_0_bits_uop_inst(lsu_io_dmem_req_bits_0_bits_uop_inst),
    .io_dmem_req_bits_0_bits_uop_debug_inst(lsu_io_dmem_req_bits_0_bits_uop_debug_inst),
    .io_dmem_req_bits_0_bits_uop_is_rvc(lsu_io_dmem_req_bits_0_bits_uop_is_rvc),
    .io_dmem_req_bits_0_bits_uop_debug_pc(lsu_io_dmem_req_bits_0_bits_uop_debug_pc),
    .io_dmem_req_bits_0_bits_uop_iq_type(lsu_io_dmem_req_bits_0_bits_uop_iq_type),
    .io_dmem_req_bits_0_bits_uop_fu_code(lsu_io_dmem_req_bits_0_bits_uop_fu_code),
    .io_dmem_req_bits_0_bits_uop_ctrl_br_type(lsu_io_dmem_req_bits_0_bits_uop_ctrl_br_type),
    .io_dmem_req_bits_0_bits_uop_ctrl_op1_sel(lsu_io_dmem_req_bits_0_bits_uop_ctrl_op1_sel),
    .io_dmem_req_bits_0_bits_uop_ctrl_op2_sel(lsu_io_dmem_req_bits_0_bits_uop_ctrl_op2_sel),
    .io_dmem_req_bits_0_bits_uop_ctrl_imm_sel(lsu_io_dmem_req_bits_0_bits_uop_ctrl_imm_sel),
    .io_dmem_req_bits_0_bits_uop_ctrl_op_fcn(lsu_io_dmem_req_bits_0_bits_uop_ctrl_op_fcn),
    .io_dmem_req_bits_0_bits_uop_ctrl_fcn_dw(lsu_io_dmem_req_bits_0_bits_uop_ctrl_fcn_dw),
    .io_dmem_req_bits_0_bits_uop_ctrl_csr_cmd(lsu_io_dmem_req_bits_0_bits_uop_ctrl_csr_cmd),
    .io_dmem_req_bits_0_bits_uop_ctrl_is_load(lsu_io_dmem_req_bits_0_bits_uop_ctrl_is_load),
    .io_dmem_req_bits_0_bits_uop_ctrl_is_sta(lsu_io_dmem_req_bits_0_bits_uop_ctrl_is_sta),
    .io_dmem_req_bits_0_bits_uop_ctrl_is_std(lsu_io_dmem_req_bits_0_bits_uop_ctrl_is_std),
    .io_dmem_req_bits_0_bits_uop_ctrl_op3_sel(lsu_io_dmem_req_bits_0_bits_uop_ctrl_op3_sel),
    .io_dmem_req_bits_0_bits_uop_iw_state(lsu_io_dmem_req_bits_0_bits_uop_iw_state),
    .io_dmem_req_bits_0_bits_uop_iw_p1_poisoned(lsu_io_dmem_req_bits_0_bits_uop_iw_p1_poisoned),
    .io_dmem_req_bits_0_bits_uop_iw_p2_poisoned(lsu_io_dmem_req_bits_0_bits_uop_iw_p2_poisoned),
    .io_dmem_req_bits_0_bits_uop_is_br(lsu_io_dmem_req_bits_0_bits_uop_is_br),
    .io_dmem_req_bits_0_bits_uop_is_jalr(lsu_io_dmem_req_bits_0_bits_uop_is_jalr),
    .io_dmem_req_bits_0_bits_uop_is_jal(lsu_io_dmem_req_bits_0_bits_uop_is_jal),
    .io_dmem_req_bits_0_bits_uop_is_sfb(lsu_io_dmem_req_bits_0_bits_uop_is_sfb),
    .io_dmem_req_bits_0_bits_uop_br_mask(lsu_io_dmem_req_bits_0_bits_uop_br_mask),
    .io_dmem_req_bits_0_bits_uop_br_tag(lsu_io_dmem_req_bits_0_bits_uop_br_tag),
    .io_dmem_req_bits_0_bits_uop_ftq_idx(lsu_io_dmem_req_bits_0_bits_uop_ftq_idx),
    .io_dmem_req_bits_0_bits_uop_edge_inst(lsu_io_dmem_req_bits_0_bits_uop_edge_inst),
    .io_dmem_req_bits_0_bits_uop_pc_lob(lsu_io_dmem_req_bits_0_bits_uop_pc_lob),
    .io_dmem_req_bits_0_bits_uop_taken(lsu_io_dmem_req_bits_0_bits_uop_taken),
    .io_dmem_req_bits_0_bits_uop_imm_packed(lsu_io_dmem_req_bits_0_bits_uop_imm_packed),
    .io_dmem_req_bits_0_bits_uop_csr_addr(lsu_io_dmem_req_bits_0_bits_uop_csr_addr),
    .io_dmem_req_bits_0_bits_uop_rob_idx(lsu_io_dmem_req_bits_0_bits_uop_rob_idx),
    .io_dmem_req_bits_0_bits_uop_ldq_idx(lsu_io_dmem_req_bits_0_bits_uop_ldq_idx),
    .io_dmem_req_bits_0_bits_uop_stq_idx(lsu_io_dmem_req_bits_0_bits_uop_stq_idx),
    .io_dmem_req_bits_0_bits_uop_rxq_idx(lsu_io_dmem_req_bits_0_bits_uop_rxq_idx),
    .io_dmem_req_bits_0_bits_uop_pdst(lsu_io_dmem_req_bits_0_bits_uop_pdst),
    .io_dmem_req_bits_0_bits_uop_prs1(lsu_io_dmem_req_bits_0_bits_uop_prs1),
    .io_dmem_req_bits_0_bits_uop_prs2(lsu_io_dmem_req_bits_0_bits_uop_prs2),
    .io_dmem_req_bits_0_bits_uop_prs3(lsu_io_dmem_req_bits_0_bits_uop_prs3),
    .io_dmem_req_bits_0_bits_uop_ppred(lsu_io_dmem_req_bits_0_bits_uop_ppred),
    .io_dmem_req_bits_0_bits_uop_prs1_busy(lsu_io_dmem_req_bits_0_bits_uop_prs1_busy),
    .io_dmem_req_bits_0_bits_uop_prs2_busy(lsu_io_dmem_req_bits_0_bits_uop_prs2_busy),
    .io_dmem_req_bits_0_bits_uop_prs3_busy(lsu_io_dmem_req_bits_0_bits_uop_prs3_busy),
    .io_dmem_req_bits_0_bits_uop_ppred_busy(lsu_io_dmem_req_bits_0_bits_uop_ppred_busy),
    .io_dmem_req_bits_0_bits_uop_stale_pdst(lsu_io_dmem_req_bits_0_bits_uop_stale_pdst),
    .io_dmem_req_bits_0_bits_uop_exception(lsu_io_dmem_req_bits_0_bits_uop_exception),
    .io_dmem_req_bits_0_bits_uop_exc_cause(lsu_io_dmem_req_bits_0_bits_uop_exc_cause),
    .io_dmem_req_bits_0_bits_uop_bypassable(lsu_io_dmem_req_bits_0_bits_uop_bypassable),
    .io_dmem_req_bits_0_bits_uop_mem_cmd(lsu_io_dmem_req_bits_0_bits_uop_mem_cmd),
    .io_dmem_req_bits_0_bits_uop_mem_size(lsu_io_dmem_req_bits_0_bits_uop_mem_size),
    .io_dmem_req_bits_0_bits_uop_mem_signed(lsu_io_dmem_req_bits_0_bits_uop_mem_signed),
    .io_dmem_req_bits_0_bits_uop_is_fence(lsu_io_dmem_req_bits_0_bits_uop_is_fence),
    .io_dmem_req_bits_0_bits_uop_is_fencei(lsu_io_dmem_req_bits_0_bits_uop_is_fencei),
    .io_dmem_req_bits_0_bits_uop_is_amo(lsu_io_dmem_req_bits_0_bits_uop_is_amo),
    .io_dmem_req_bits_0_bits_uop_uses_ldq(lsu_io_dmem_req_bits_0_bits_uop_uses_ldq),
    .io_dmem_req_bits_0_bits_uop_uses_stq(lsu_io_dmem_req_bits_0_bits_uop_uses_stq),
    .io_dmem_req_bits_0_bits_uop_is_sys_pc2epc(lsu_io_dmem_req_bits_0_bits_uop_is_sys_pc2epc),
    .io_dmem_req_bits_0_bits_uop_is_unique(lsu_io_dmem_req_bits_0_bits_uop_is_unique),
    .io_dmem_req_bits_0_bits_uop_flush_on_commit(lsu_io_dmem_req_bits_0_bits_uop_flush_on_commit),
    .io_dmem_req_bits_0_bits_uop_ldst_is_rs1(lsu_io_dmem_req_bits_0_bits_uop_ldst_is_rs1),
    .io_dmem_req_bits_0_bits_uop_ldst(lsu_io_dmem_req_bits_0_bits_uop_ldst),
    .io_dmem_req_bits_0_bits_uop_lrs1(lsu_io_dmem_req_bits_0_bits_uop_lrs1),
    .io_dmem_req_bits_0_bits_uop_lrs2(lsu_io_dmem_req_bits_0_bits_uop_lrs2),
    .io_dmem_req_bits_0_bits_uop_lrs3(lsu_io_dmem_req_bits_0_bits_uop_lrs3),
    .io_dmem_req_bits_0_bits_uop_ldst_val(lsu_io_dmem_req_bits_0_bits_uop_ldst_val),
    .io_dmem_req_bits_0_bits_uop_dst_rtype(lsu_io_dmem_req_bits_0_bits_uop_dst_rtype),
    .io_dmem_req_bits_0_bits_uop_lrs1_rtype(lsu_io_dmem_req_bits_0_bits_uop_lrs1_rtype),
    .io_dmem_req_bits_0_bits_uop_lrs2_rtype(lsu_io_dmem_req_bits_0_bits_uop_lrs2_rtype),
    .io_dmem_req_bits_0_bits_uop_frs3_en(lsu_io_dmem_req_bits_0_bits_uop_frs3_en),
    .io_dmem_req_bits_0_bits_uop_fp_val(lsu_io_dmem_req_bits_0_bits_uop_fp_val),
    .io_dmem_req_bits_0_bits_uop_fp_single(lsu_io_dmem_req_bits_0_bits_uop_fp_single),
    .io_dmem_req_bits_0_bits_uop_xcpt_pf_if(lsu_io_dmem_req_bits_0_bits_uop_xcpt_pf_if),
    .io_dmem_req_bits_0_bits_uop_xcpt_ae_if(lsu_io_dmem_req_bits_0_bits_uop_xcpt_ae_if),
    .io_dmem_req_bits_0_bits_uop_xcpt_ma_if(lsu_io_dmem_req_bits_0_bits_uop_xcpt_ma_if),
    .io_dmem_req_bits_0_bits_uop_bp_debug_if(lsu_io_dmem_req_bits_0_bits_uop_bp_debug_if),
    .io_dmem_req_bits_0_bits_uop_bp_xcpt_if(lsu_io_dmem_req_bits_0_bits_uop_bp_xcpt_if),
    .io_dmem_req_bits_0_bits_uop_debug_fsrc(lsu_io_dmem_req_bits_0_bits_uop_debug_fsrc),
    .io_dmem_req_bits_0_bits_uop_debug_tsrc(lsu_io_dmem_req_bits_0_bits_uop_debug_tsrc),
    .io_dmem_req_bits_0_bits_addr(lsu_io_dmem_req_bits_0_bits_addr),
    .io_dmem_req_bits_0_bits_data(lsu_io_dmem_req_bits_0_bits_data),
    .io_dmem_req_bits_0_bits_is_hella(lsu_io_dmem_req_bits_0_bits_is_hella),
    .io_dmem_s1_kill_0(lsu_io_dmem_s1_kill_0),
    .io_dmem_resp_0_valid(lsu_io_dmem_resp_0_valid),
    .io_dmem_resp_0_bits_uop_switch(lsu_io_dmem_resp_0_bits_uop_switch),
    .io_dmem_resp_0_bits_uop_switch_off(lsu_io_dmem_resp_0_bits_uop_switch_off),
    .io_dmem_resp_0_bits_uop_is_unicore(lsu_io_dmem_resp_0_bits_uop_is_unicore),
    .io_dmem_resp_0_bits_uop_shift(lsu_io_dmem_resp_0_bits_uop_shift),
    .io_dmem_resp_0_bits_uop_lrs3_rtype(lsu_io_dmem_resp_0_bits_uop_lrs3_rtype),
    .io_dmem_resp_0_bits_uop_rflag(lsu_io_dmem_resp_0_bits_uop_rflag),
    .io_dmem_resp_0_bits_uop_wflag(lsu_io_dmem_resp_0_bits_uop_wflag),
    .io_dmem_resp_0_bits_uop_prflag(lsu_io_dmem_resp_0_bits_uop_prflag),
    .io_dmem_resp_0_bits_uop_pwflag(lsu_io_dmem_resp_0_bits_uop_pwflag),
    .io_dmem_resp_0_bits_uop_pflag_busy(lsu_io_dmem_resp_0_bits_uop_pflag_busy),
    .io_dmem_resp_0_bits_uop_stale_pflag(lsu_io_dmem_resp_0_bits_uop_stale_pflag),
    .io_dmem_resp_0_bits_uop_op1_sel(lsu_io_dmem_resp_0_bits_uop_op1_sel),
    .io_dmem_resp_0_bits_uop_op2_sel(lsu_io_dmem_resp_0_bits_uop_op2_sel),
    .io_dmem_resp_0_bits_uop_split_num(lsu_io_dmem_resp_0_bits_uop_split_num),
    .io_dmem_resp_0_bits_uop_self_index(lsu_io_dmem_resp_0_bits_uop_self_index),
    .io_dmem_resp_0_bits_uop_rob_inst_idx(lsu_io_dmem_resp_0_bits_uop_rob_inst_idx),
    .io_dmem_resp_0_bits_uop_address_num(lsu_io_dmem_resp_0_bits_uop_address_num),
    .io_dmem_resp_0_bits_uop_uopc(lsu_io_dmem_resp_0_bits_uop_uopc),
    .io_dmem_resp_0_bits_uop_inst(lsu_io_dmem_resp_0_bits_uop_inst),
    .io_dmem_resp_0_bits_uop_debug_inst(lsu_io_dmem_resp_0_bits_uop_debug_inst),
    .io_dmem_resp_0_bits_uop_is_rvc(lsu_io_dmem_resp_0_bits_uop_is_rvc),
    .io_dmem_resp_0_bits_uop_debug_pc(lsu_io_dmem_resp_0_bits_uop_debug_pc),
    .io_dmem_resp_0_bits_uop_iq_type(lsu_io_dmem_resp_0_bits_uop_iq_type),
    .io_dmem_resp_0_bits_uop_fu_code(lsu_io_dmem_resp_0_bits_uop_fu_code),
    .io_dmem_resp_0_bits_uop_ctrl_br_type(lsu_io_dmem_resp_0_bits_uop_ctrl_br_type),
    .io_dmem_resp_0_bits_uop_ctrl_op1_sel(lsu_io_dmem_resp_0_bits_uop_ctrl_op1_sel),
    .io_dmem_resp_0_bits_uop_ctrl_op2_sel(lsu_io_dmem_resp_0_bits_uop_ctrl_op2_sel),
    .io_dmem_resp_0_bits_uop_ctrl_imm_sel(lsu_io_dmem_resp_0_bits_uop_ctrl_imm_sel),
    .io_dmem_resp_0_bits_uop_ctrl_op_fcn(lsu_io_dmem_resp_0_bits_uop_ctrl_op_fcn),
    .io_dmem_resp_0_bits_uop_ctrl_fcn_dw(lsu_io_dmem_resp_0_bits_uop_ctrl_fcn_dw),
    .io_dmem_resp_0_bits_uop_ctrl_csr_cmd(lsu_io_dmem_resp_0_bits_uop_ctrl_csr_cmd),
    .io_dmem_resp_0_bits_uop_ctrl_is_load(lsu_io_dmem_resp_0_bits_uop_ctrl_is_load),
    .io_dmem_resp_0_bits_uop_ctrl_is_sta(lsu_io_dmem_resp_0_bits_uop_ctrl_is_sta),
    .io_dmem_resp_0_bits_uop_ctrl_is_std(lsu_io_dmem_resp_0_bits_uop_ctrl_is_std),
    .io_dmem_resp_0_bits_uop_ctrl_op3_sel(lsu_io_dmem_resp_0_bits_uop_ctrl_op3_sel),
    .io_dmem_resp_0_bits_uop_iw_state(lsu_io_dmem_resp_0_bits_uop_iw_state),
    .io_dmem_resp_0_bits_uop_iw_p1_poisoned(lsu_io_dmem_resp_0_bits_uop_iw_p1_poisoned),
    .io_dmem_resp_0_bits_uop_iw_p2_poisoned(lsu_io_dmem_resp_0_bits_uop_iw_p2_poisoned),
    .io_dmem_resp_0_bits_uop_is_br(lsu_io_dmem_resp_0_bits_uop_is_br),
    .io_dmem_resp_0_bits_uop_is_jalr(lsu_io_dmem_resp_0_bits_uop_is_jalr),
    .io_dmem_resp_0_bits_uop_is_jal(lsu_io_dmem_resp_0_bits_uop_is_jal),
    .io_dmem_resp_0_bits_uop_is_sfb(lsu_io_dmem_resp_0_bits_uop_is_sfb),
    .io_dmem_resp_0_bits_uop_br_mask(lsu_io_dmem_resp_0_bits_uop_br_mask),
    .io_dmem_resp_0_bits_uop_br_tag(lsu_io_dmem_resp_0_bits_uop_br_tag),
    .io_dmem_resp_0_bits_uop_ftq_idx(lsu_io_dmem_resp_0_bits_uop_ftq_idx),
    .io_dmem_resp_0_bits_uop_edge_inst(lsu_io_dmem_resp_0_bits_uop_edge_inst),
    .io_dmem_resp_0_bits_uop_pc_lob(lsu_io_dmem_resp_0_bits_uop_pc_lob),
    .io_dmem_resp_0_bits_uop_taken(lsu_io_dmem_resp_0_bits_uop_taken),
    .io_dmem_resp_0_bits_uop_imm_packed(lsu_io_dmem_resp_0_bits_uop_imm_packed),
    .io_dmem_resp_0_bits_uop_csr_addr(lsu_io_dmem_resp_0_bits_uop_csr_addr),
    .io_dmem_resp_0_bits_uop_rob_idx(lsu_io_dmem_resp_0_bits_uop_rob_idx),
    .io_dmem_resp_0_bits_uop_ldq_idx(lsu_io_dmem_resp_0_bits_uop_ldq_idx),
    .io_dmem_resp_0_bits_uop_stq_idx(lsu_io_dmem_resp_0_bits_uop_stq_idx),
    .io_dmem_resp_0_bits_uop_rxq_idx(lsu_io_dmem_resp_0_bits_uop_rxq_idx),
    .io_dmem_resp_0_bits_uop_pdst(lsu_io_dmem_resp_0_bits_uop_pdst),
    .io_dmem_resp_0_bits_uop_prs1(lsu_io_dmem_resp_0_bits_uop_prs1),
    .io_dmem_resp_0_bits_uop_prs2(lsu_io_dmem_resp_0_bits_uop_prs2),
    .io_dmem_resp_0_bits_uop_prs3(lsu_io_dmem_resp_0_bits_uop_prs3),
    .io_dmem_resp_0_bits_uop_ppred(lsu_io_dmem_resp_0_bits_uop_ppred),
    .io_dmem_resp_0_bits_uop_prs1_busy(lsu_io_dmem_resp_0_bits_uop_prs1_busy),
    .io_dmem_resp_0_bits_uop_prs2_busy(lsu_io_dmem_resp_0_bits_uop_prs2_busy),
    .io_dmem_resp_0_bits_uop_prs3_busy(lsu_io_dmem_resp_0_bits_uop_prs3_busy),
    .io_dmem_resp_0_bits_uop_ppred_busy(lsu_io_dmem_resp_0_bits_uop_ppred_busy),
    .io_dmem_resp_0_bits_uop_stale_pdst(lsu_io_dmem_resp_0_bits_uop_stale_pdst),
    .io_dmem_resp_0_bits_uop_exception(lsu_io_dmem_resp_0_bits_uop_exception),
    .io_dmem_resp_0_bits_uop_exc_cause(lsu_io_dmem_resp_0_bits_uop_exc_cause),
    .io_dmem_resp_0_bits_uop_bypassable(lsu_io_dmem_resp_0_bits_uop_bypassable),
    .io_dmem_resp_0_bits_uop_mem_cmd(lsu_io_dmem_resp_0_bits_uop_mem_cmd),
    .io_dmem_resp_0_bits_uop_mem_size(lsu_io_dmem_resp_0_bits_uop_mem_size),
    .io_dmem_resp_0_bits_uop_mem_signed(lsu_io_dmem_resp_0_bits_uop_mem_signed),
    .io_dmem_resp_0_bits_uop_is_fence(lsu_io_dmem_resp_0_bits_uop_is_fence),
    .io_dmem_resp_0_bits_uop_is_fencei(lsu_io_dmem_resp_0_bits_uop_is_fencei),
    .io_dmem_resp_0_bits_uop_is_amo(lsu_io_dmem_resp_0_bits_uop_is_amo),
    .io_dmem_resp_0_bits_uop_uses_ldq(lsu_io_dmem_resp_0_bits_uop_uses_ldq),
    .io_dmem_resp_0_bits_uop_uses_stq(lsu_io_dmem_resp_0_bits_uop_uses_stq),
    .io_dmem_resp_0_bits_uop_is_sys_pc2epc(lsu_io_dmem_resp_0_bits_uop_is_sys_pc2epc),
    .io_dmem_resp_0_bits_uop_is_unique(lsu_io_dmem_resp_0_bits_uop_is_unique),
    .io_dmem_resp_0_bits_uop_flush_on_commit(lsu_io_dmem_resp_0_bits_uop_flush_on_commit),
    .io_dmem_resp_0_bits_uop_ldst_is_rs1(lsu_io_dmem_resp_0_bits_uop_ldst_is_rs1),
    .io_dmem_resp_0_bits_uop_ldst(lsu_io_dmem_resp_0_bits_uop_ldst),
    .io_dmem_resp_0_bits_uop_lrs1(lsu_io_dmem_resp_0_bits_uop_lrs1),
    .io_dmem_resp_0_bits_uop_lrs2(lsu_io_dmem_resp_0_bits_uop_lrs2),
    .io_dmem_resp_0_bits_uop_lrs3(lsu_io_dmem_resp_0_bits_uop_lrs3),
    .io_dmem_resp_0_bits_uop_ldst_val(lsu_io_dmem_resp_0_bits_uop_ldst_val),
    .io_dmem_resp_0_bits_uop_dst_rtype(lsu_io_dmem_resp_0_bits_uop_dst_rtype),
    .io_dmem_resp_0_bits_uop_lrs1_rtype(lsu_io_dmem_resp_0_bits_uop_lrs1_rtype),
    .io_dmem_resp_0_bits_uop_lrs2_rtype(lsu_io_dmem_resp_0_bits_uop_lrs2_rtype),
    .io_dmem_resp_0_bits_uop_frs3_en(lsu_io_dmem_resp_0_bits_uop_frs3_en),
    .io_dmem_resp_0_bits_uop_fp_val(lsu_io_dmem_resp_0_bits_uop_fp_val),
    .io_dmem_resp_0_bits_uop_fp_single(lsu_io_dmem_resp_0_bits_uop_fp_single),
    .io_dmem_resp_0_bits_uop_xcpt_pf_if(lsu_io_dmem_resp_0_bits_uop_xcpt_pf_if),
    .io_dmem_resp_0_bits_uop_xcpt_ae_if(lsu_io_dmem_resp_0_bits_uop_xcpt_ae_if),
    .io_dmem_resp_0_bits_uop_xcpt_ma_if(lsu_io_dmem_resp_0_bits_uop_xcpt_ma_if),
    .io_dmem_resp_0_bits_uop_bp_debug_if(lsu_io_dmem_resp_0_bits_uop_bp_debug_if),
    .io_dmem_resp_0_bits_uop_bp_xcpt_if(lsu_io_dmem_resp_0_bits_uop_bp_xcpt_if),
    .io_dmem_resp_0_bits_uop_debug_fsrc(lsu_io_dmem_resp_0_bits_uop_debug_fsrc),
    .io_dmem_resp_0_bits_uop_debug_tsrc(lsu_io_dmem_resp_0_bits_uop_debug_tsrc),
    .io_dmem_resp_0_bits_data(lsu_io_dmem_resp_0_bits_data),
    .io_dmem_resp_0_bits_is_hella(lsu_io_dmem_resp_0_bits_is_hella),
    .io_dmem_nack_0_valid(lsu_io_dmem_nack_0_valid),
    .io_dmem_nack_0_bits_uop_switch(lsu_io_dmem_nack_0_bits_uop_switch),
    .io_dmem_nack_0_bits_uop_switch_off(lsu_io_dmem_nack_0_bits_uop_switch_off),
    .io_dmem_nack_0_bits_uop_is_unicore(lsu_io_dmem_nack_0_bits_uop_is_unicore),
    .io_dmem_nack_0_bits_uop_shift(lsu_io_dmem_nack_0_bits_uop_shift),
    .io_dmem_nack_0_bits_uop_lrs3_rtype(lsu_io_dmem_nack_0_bits_uop_lrs3_rtype),
    .io_dmem_nack_0_bits_uop_rflag(lsu_io_dmem_nack_0_bits_uop_rflag),
    .io_dmem_nack_0_bits_uop_wflag(lsu_io_dmem_nack_0_bits_uop_wflag),
    .io_dmem_nack_0_bits_uop_prflag(lsu_io_dmem_nack_0_bits_uop_prflag),
    .io_dmem_nack_0_bits_uop_pwflag(lsu_io_dmem_nack_0_bits_uop_pwflag),
    .io_dmem_nack_0_bits_uop_pflag_busy(lsu_io_dmem_nack_0_bits_uop_pflag_busy),
    .io_dmem_nack_0_bits_uop_stale_pflag(lsu_io_dmem_nack_0_bits_uop_stale_pflag),
    .io_dmem_nack_0_bits_uop_op1_sel(lsu_io_dmem_nack_0_bits_uop_op1_sel),
    .io_dmem_nack_0_bits_uop_op2_sel(lsu_io_dmem_nack_0_bits_uop_op2_sel),
    .io_dmem_nack_0_bits_uop_split_num(lsu_io_dmem_nack_0_bits_uop_split_num),
    .io_dmem_nack_0_bits_uop_self_index(lsu_io_dmem_nack_0_bits_uop_self_index),
    .io_dmem_nack_0_bits_uop_rob_inst_idx(lsu_io_dmem_nack_0_bits_uop_rob_inst_idx),
    .io_dmem_nack_0_bits_uop_address_num(lsu_io_dmem_nack_0_bits_uop_address_num),
    .io_dmem_nack_0_bits_uop_uopc(lsu_io_dmem_nack_0_bits_uop_uopc),
    .io_dmem_nack_0_bits_uop_inst(lsu_io_dmem_nack_0_bits_uop_inst),
    .io_dmem_nack_0_bits_uop_debug_inst(lsu_io_dmem_nack_0_bits_uop_debug_inst),
    .io_dmem_nack_0_bits_uop_is_rvc(lsu_io_dmem_nack_0_bits_uop_is_rvc),
    .io_dmem_nack_0_bits_uop_debug_pc(lsu_io_dmem_nack_0_bits_uop_debug_pc),
    .io_dmem_nack_0_bits_uop_iq_type(lsu_io_dmem_nack_0_bits_uop_iq_type),
    .io_dmem_nack_0_bits_uop_fu_code(lsu_io_dmem_nack_0_bits_uop_fu_code),
    .io_dmem_nack_0_bits_uop_ctrl_br_type(lsu_io_dmem_nack_0_bits_uop_ctrl_br_type),
    .io_dmem_nack_0_bits_uop_ctrl_op1_sel(lsu_io_dmem_nack_0_bits_uop_ctrl_op1_sel),
    .io_dmem_nack_0_bits_uop_ctrl_op2_sel(lsu_io_dmem_nack_0_bits_uop_ctrl_op2_sel),
    .io_dmem_nack_0_bits_uop_ctrl_imm_sel(lsu_io_dmem_nack_0_bits_uop_ctrl_imm_sel),
    .io_dmem_nack_0_bits_uop_ctrl_op_fcn(lsu_io_dmem_nack_0_bits_uop_ctrl_op_fcn),
    .io_dmem_nack_0_bits_uop_ctrl_fcn_dw(lsu_io_dmem_nack_0_bits_uop_ctrl_fcn_dw),
    .io_dmem_nack_0_bits_uop_ctrl_csr_cmd(lsu_io_dmem_nack_0_bits_uop_ctrl_csr_cmd),
    .io_dmem_nack_0_bits_uop_ctrl_is_load(lsu_io_dmem_nack_0_bits_uop_ctrl_is_load),
    .io_dmem_nack_0_bits_uop_ctrl_is_sta(lsu_io_dmem_nack_0_bits_uop_ctrl_is_sta),
    .io_dmem_nack_0_bits_uop_ctrl_is_std(lsu_io_dmem_nack_0_bits_uop_ctrl_is_std),
    .io_dmem_nack_0_bits_uop_ctrl_op3_sel(lsu_io_dmem_nack_0_bits_uop_ctrl_op3_sel),
    .io_dmem_nack_0_bits_uop_iw_state(lsu_io_dmem_nack_0_bits_uop_iw_state),
    .io_dmem_nack_0_bits_uop_iw_p1_poisoned(lsu_io_dmem_nack_0_bits_uop_iw_p1_poisoned),
    .io_dmem_nack_0_bits_uop_iw_p2_poisoned(lsu_io_dmem_nack_0_bits_uop_iw_p2_poisoned),
    .io_dmem_nack_0_bits_uop_is_br(lsu_io_dmem_nack_0_bits_uop_is_br),
    .io_dmem_nack_0_bits_uop_is_jalr(lsu_io_dmem_nack_0_bits_uop_is_jalr),
    .io_dmem_nack_0_bits_uop_is_jal(lsu_io_dmem_nack_0_bits_uop_is_jal),
    .io_dmem_nack_0_bits_uop_is_sfb(lsu_io_dmem_nack_0_bits_uop_is_sfb),
    .io_dmem_nack_0_bits_uop_br_mask(lsu_io_dmem_nack_0_bits_uop_br_mask),
    .io_dmem_nack_0_bits_uop_br_tag(lsu_io_dmem_nack_0_bits_uop_br_tag),
    .io_dmem_nack_0_bits_uop_ftq_idx(lsu_io_dmem_nack_0_bits_uop_ftq_idx),
    .io_dmem_nack_0_bits_uop_edge_inst(lsu_io_dmem_nack_0_bits_uop_edge_inst),
    .io_dmem_nack_0_bits_uop_pc_lob(lsu_io_dmem_nack_0_bits_uop_pc_lob),
    .io_dmem_nack_0_bits_uop_taken(lsu_io_dmem_nack_0_bits_uop_taken),
    .io_dmem_nack_0_bits_uop_imm_packed(lsu_io_dmem_nack_0_bits_uop_imm_packed),
    .io_dmem_nack_0_bits_uop_csr_addr(lsu_io_dmem_nack_0_bits_uop_csr_addr),
    .io_dmem_nack_0_bits_uop_rob_idx(lsu_io_dmem_nack_0_bits_uop_rob_idx),
    .io_dmem_nack_0_bits_uop_ldq_idx(lsu_io_dmem_nack_0_bits_uop_ldq_idx),
    .io_dmem_nack_0_bits_uop_stq_idx(lsu_io_dmem_nack_0_bits_uop_stq_idx),
    .io_dmem_nack_0_bits_uop_rxq_idx(lsu_io_dmem_nack_0_bits_uop_rxq_idx),
    .io_dmem_nack_0_bits_uop_pdst(lsu_io_dmem_nack_0_bits_uop_pdst),
    .io_dmem_nack_0_bits_uop_prs1(lsu_io_dmem_nack_0_bits_uop_prs1),
    .io_dmem_nack_0_bits_uop_prs2(lsu_io_dmem_nack_0_bits_uop_prs2),
    .io_dmem_nack_0_bits_uop_prs3(lsu_io_dmem_nack_0_bits_uop_prs3),
    .io_dmem_nack_0_bits_uop_ppred(lsu_io_dmem_nack_0_bits_uop_ppred),
    .io_dmem_nack_0_bits_uop_prs1_busy(lsu_io_dmem_nack_0_bits_uop_prs1_busy),
    .io_dmem_nack_0_bits_uop_prs2_busy(lsu_io_dmem_nack_0_bits_uop_prs2_busy),
    .io_dmem_nack_0_bits_uop_prs3_busy(lsu_io_dmem_nack_0_bits_uop_prs3_busy),
    .io_dmem_nack_0_bits_uop_ppred_busy(lsu_io_dmem_nack_0_bits_uop_ppred_busy),
    .io_dmem_nack_0_bits_uop_stale_pdst(lsu_io_dmem_nack_0_bits_uop_stale_pdst),
    .io_dmem_nack_0_bits_uop_exception(lsu_io_dmem_nack_0_bits_uop_exception),
    .io_dmem_nack_0_bits_uop_exc_cause(lsu_io_dmem_nack_0_bits_uop_exc_cause),
    .io_dmem_nack_0_bits_uop_bypassable(lsu_io_dmem_nack_0_bits_uop_bypassable),
    .io_dmem_nack_0_bits_uop_mem_cmd(lsu_io_dmem_nack_0_bits_uop_mem_cmd),
    .io_dmem_nack_0_bits_uop_mem_size(lsu_io_dmem_nack_0_bits_uop_mem_size),
    .io_dmem_nack_0_bits_uop_mem_signed(lsu_io_dmem_nack_0_bits_uop_mem_signed),
    .io_dmem_nack_0_bits_uop_is_fence(lsu_io_dmem_nack_0_bits_uop_is_fence),
    .io_dmem_nack_0_bits_uop_is_fencei(lsu_io_dmem_nack_0_bits_uop_is_fencei),
    .io_dmem_nack_0_bits_uop_is_amo(lsu_io_dmem_nack_0_bits_uop_is_amo),
    .io_dmem_nack_0_bits_uop_uses_ldq(lsu_io_dmem_nack_0_bits_uop_uses_ldq),
    .io_dmem_nack_0_bits_uop_uses_stq(lsu_io_dmem_nack_0_bits_uop_uses_stq),
    .io_dmem_nack_0_bits_uop_is_sys_pc2epc(lsu_io_dmem_nack_0_bits_uop_is_sys_pc2epc),
    .io_dmem_nack_0_bits_uop_is_unique(lsu_io_dmem_nack_0_bits_uop_is_unique),
    .io_dmem_nack_0_bits_uop_flush_on_commit(lsu_io_dmem_nack_0_bits_uop_flush_on_commit),
    .io_dmem_nack_0_bits_uop_ldst_is_rs1(lsu_io_dmem_nack_0_bits_uop_ldst_is_rs1),
    .io_dmem_nack_0_bits_uop_ldst(lsu_io_dmem_nack_0_bits_uop_ldst),
    .io_dmem_nack_0_bits_uop_lrs1(lsu_io_dmem_nack_0_bits_uop_lrs1),
    .io_dmem_nack_0_bits_uop_lrs2(lsu_io_dmem_nack_0_bits_uop_lrs2),
    .io_dmem_nack_0_bits_uop_lrs3(lsu_io_dmem_nack_0_bits_uop_lrs3),
    .io_dmem_nack_0_bits_uop_ldst_val(lsu_io_dmem_nack_0_bits_uop_ldst_val),
    .io_dmem_nack_0_bits_uop_dst_rtype(lsu_io_dmem_nack_0_bits_uop_dst_rtype),
    .io_dmem_nack_0_bits_uop_lrs1_rtype(lsu_io_dmem_nack_0_bits_uop_lrs1_rtype),
    .io_dmem_nack_0_bits_uop_lrs2_rtype(lsu_io_dmem_nack_0_bits_uop_lrs2_rtype),
    .io_dmem_nack_0_bits_uop_frs3_en(lsu_io_dmem_nack_0_bits_uop_frs3_en),
    .io_dmem_nack_0_bits_uop_fp_val(lsu_io_dmem_nack_0_bits_uop_fp_val),
    .io_dmem_nack_0_bits_uop_fp_single(lsu_io_dmem_nack_0_bits_uop_fp_single),
    .io_dmem_nack_0_bits_uop_xcpt_pf_if(lsu_io_dmem_nack_0_bits_uop_xcpt_pf_if),
    .io_dmem_nack_0_bits_uop_xcpt_ae_if(lsu_io_dmem_nack_0_bits_uop_xcpt_ae_if),
    .io_dmem_nack_0_bits_uop_xcpt_ma_if(lsu_io_dmem_nack_0_bits_uop_xcpt_ma_if),
    .io_dmem_nack_0_bits_uop_bp_debug_if(lsu_io_dmem_nack_0_bits_uop_bp_debug_if),
    .io_dmem_nack_0_bits_uop_bp_xcpt_if(lsu_io_dmem_nack_0_bits_uop_bp_xcpt_if),
    .io_dmem_nack_0_bits_uop_debug_fsrc(lsu_io_dmem_nack_0_bits_uop_debug_fsrc),
    .io_dmem_nack_0_bits_uop_debug_tsrc(lsu_io_dmem_nack_0_bits_uop_debug_tsrc),
    .io_dmem_nack_0_bits_addr(lsu_io_dmem_nack_0_bits_addr),
    .io_dmem_nack_0_bits_data(lsu_io_dmem_nack_0_bits_data),
    .io_dmem_nack_0_bits_is_hella(lsu_io_dmem_nack_0_bits_is_hella),
    .io_dmem_brupdate_b1_resolve_mask(lsu_io_dmem_brupdate_b1_resolve_mask),
    .io_dmem_brupdate_b1_mispredict_mask(lsu_io_dmem_brupdate_b1_mispredict_mask),
    .io_dmem_brupdate_b2_uop_switch(lsu_io_dmem_brupdate_b2_uop_switch),
    .io_dmem_brupdate_b2_uop_switch_off(lsu_io_dmem_brupdate_b2_uop_switch_off),
    .io_dmem_brupdate_b2_uop_is_unicore(lsu_io_dmem_brupdate_b2_uop_is_unicore),
    .io_dmem_brupdate_b2_uop_shift(lsu_io_dmem_brupdate_b2_uop_shift),
    .io_dmem_brupdate_b2_uop_lrs3_rtype(lsu_io_dmem_brupdate_b2_uop_lrs3_rtype),
    .io_dmem_brupdate_b2_uop_rflag(lsu_io_dmem_brupdate_b2_uop_rflag),
    .io_dmem_brupdate_b2_uop_wflag(lsu_io_dmem_brupdate_b2_uop_wflag),
    .io_dmem_brupdate_b2_uop_prflag(lsu_io_dmem_brupdate_b2_uop_prflag),
    .io_dmem_brupdate_b2_uop_pwflag(lsu_io_dmem_brupdate_b2_uop_pwflag),
    .io_dmem_brupdate_b2_uop_pflag_busy(lsu_io_dmem_brupdate_b2_uop_pflag_busy),
    .io_dmem_brupdate_b2_uop_stale_pflag(lsu_io_dmem_brupdate_b2_uop_stale_pflag),
    .io_dmem_brupdate_b2_uop_op1_sel(lsu_io_dmem_brupdate_b2_uop_op1_sel),
    .io_dmem_brupdate_b2_uop_op2_sel(lsu_io_dmem_brupdate_b2_uop_op2_sel),
    .io_dmem_brupdate_b2_uop_split_num(lsu_io_dmem_brupdate_b2_uop_split_num),
    .io_dmem_brupdate_b2_uop_self_index(lsu_io_dmem_brupdate_b2_uop_self_index),
    .io_dmem_brupdate_b2_uop_rob_inst_idx(lsu_io_dmem_brupdate_b2_uop_rob_inst_idx),
    .io_dmem_brupdate_b2_uop_address_num(lsu_io_dmem_brupdate_b2_uop_address_num),
    .io_dmem_brupdate_b2_uop_uopc(lsu_io_dmem_brupdate_b2_uop_uopc),
    .io_dmem_brupdate_b2_uop_inst(lsu_io_dmem_brupdate_b2_uop_inst),
    .io_dmem_brupdate_b2_uop_debug_inst(lsu_io_dmem_brupdate_b2_uop_debug_inst),
    .io_dmem_brupdate_b2_uop_is_rvc(lsu_io_dmem_brupdate_b2_uop_is_rvc),
    .io_dmem_brupdate_b2_uop_debug_pc(lsu_io_dmem_brupdate_b2_uop_debug_pc),
    .io_dmem_brupdate_b2_uop_iq_type(lsu_io_dmem_brupdate_b2_uop_iq_type),
    .io_dmem_brupdate_b2_uop_fu_code(lsu_io_dmem_brupdate_b2_uop_fu_code),
    .io_dmem_brupdate_b2_uop_ctrl_br_type(lsu_io_dmem_brupdate_b2_uop_ctrl_br_type),
    .io_dmem_brupdate_b2_uop_ctrl_op1_sel(lsu_io_dmem_brupdate_b2_uop_ctrl_op1_sel),
    .io_dmem_brupdate_b2_uop_ctrl_op2_sel(lsu_io_dmem_brupdate_b2_uop_ctrl_op2_sel),
    .io_dmem_brupdate_b2_uop_ctrl_imm_sel(lsu_io_dmem_brupdate_b2_uop_ctrl_imm_sel),
    .io_dmem_brupdate_b2_uop_ctrl_op_fcn(lsu_io_dmem_brupdate_b2_uop_ctrl_op_fcn),
    .io_dmem_brupdate_b2_uop_ctrl_fcn_dw(lsu_io_dmem_brupdate_b2_uop_ctrl_fcn_dw),
    .io_dmem_brupdate_b2_uop_ctrl_csr_cmd(lsu_io_dmem_brupdate_b2_uop_ctrl_csr_cmd),
    .io_dmem_brupdate_b2_uop_ctrl_is_load(lsu_io_dmem_brupdate_b2_uop_ctrl_is_load),
    .io_dmem_brupdate_b2_uop_ctrl_is_sta(lsu_io_dmem_brupdate_b2_uop_ctrl_is_sta),
    .io_dmem_brupdate_b2_uop_ctrl_is_std(lsu_io_dmem_brupdate_b2_uop_ctrl_is_std),
    .io_dmem_brupdate_b2_uop_ctrl_op3_sel(lsu_io_dmem_brupdate_b2_uop_ctrl_op3_sel),
    .io_dmem_brupdate_b2_uop_iw_state(lsu_io_dmem_brupdate_b2_uop_iw_state),
    .io_dmem_brupdate_b2_uop_iw_p1_poisoned(lsu_io_dmem_brupdate_b2_uop_iw_p1_poisoned),
    .io_dmem_brupdate_b2_uop_iw_p2_poisoned(lsu_io_dmem_brupdate_b2_uop_iw_p2_poisoned),
    .io_dmem_brupdate_b2_uop_is_br(lsu_io_dmem_brupdate_b2_uop_is_br),
    .io_dmem_brupdate_b2_uop_is_jalr(lsu_io_dmem_brupdate_b2_uop_is_jalr),
    .io_dmem_brupdate_b2_uop_is_jal(lsu_io_dmem_brupdate_b2_uop_is_jal),
    .io_dmem_brupdate_b2_uop_is_sfb(lsu_io_dmem_brupdate_b2_uop_is_sfb),
    .io_dmem_brupdate_b2_uop_br_mask(lsu_io_dmem_brupdate_b2_uop_br_mask),
    .io_dmem_brupdate_b2_uop_br_tag(lsu_io_dmem_brupdate_b2_uop_br_tag),
    .io_dmem_brupdate_b2_uop_ftq_idx(lsu_io_dmem_brupdate_b2_uop_ftq_idx),
    .io_dmem_brupdate_b2_uop_edge_inst(lsu_io_dmem_brupdate_b2_uop_edge_inst),
    .io_dmem_brupdate_b2_uop_pc_lob(lsu_io_dmem_brupdate_b2_uop_pc_lob),
    .io_dmem_brupdate_b2_uop_taken(lsu_io_dmem_brupdate_b2_uop_taken),
    .io_dmem_brupdate_b2_uop_imm_packed(lsu_io_dmem_brupdate_b2_uop_imm_packed),
    .io_dmem_brupdate_b2_uop_csr_addr(lsu_io_dmem_brupdate_b2_uop_csr_addr),
    .io_dmem_brupdate_b2_uop_rob_idx(lsu_io_dmem_brupdate_b2_uop_rob_idx),
    .io_dmem_brupdate_b2_uop_ldq_idx(lsu_io_dmem_brupdate_b2_uop_ldq_idx),
    .io_dmem_brupdate_b2_uop_stq_idx(lsu_io_dmem_brupdate_b2_uop_stq_idx),
    .io_dmem_brupdate_b2_uop_rxq_idx(lsu_io_dmem_brupdate_b2_uop_rxq_idx),
    .io_dmem_brupdate_b2_uop_pdst(lsu_io_dmem_brupdate_b2_uop_pdst),
    .io_dmem_brupdate_b2_uop_prs1(lsu_io_dmem_brupdate_b2_uop_prs1),
    .io_dmem_brupdate_b2_uop_prs2(lsu_io_dmem_brupdate_b2_uop_prs2),
    .io_dmem_brupdate_b2_uop_prs3(lsu_io_dmem_brupdate_b2_uop_prs3),
    .io_dmem_brupdate_b2_uop_ppred(lsu_io_dmem_brupdate_b2_uop_ppred),
    .io_dmem_brupdate_b2_uop_prs1_busy(lsu_io_dmem_brupdate_b2_uop_prs1_busy),
    .io_dmem_brupdate_b2_uop_prs2_busy(lsu_io_dmem_brupdate_b2_uop_prs2_busy),
    .io_dmem_brupdate_b2_uop_prs3_busy(lsu_io_dmem_brupdate_b2_uop_prs3_busy),
    .io_dmem_brupdate_b2_uop_ppred_busy(lsu_io_dmem_brupdate_b2_uop_ppred_busy),
    .io_dmem_brupdate_b2_uop_stale_pdst(lsu_io_dmem_brupdate_b2_uop_stale_pdst),
    .io_dmem_brupdate_b2_uop_exception(lsu_io_dmem_brupdate_b2_uop_exception),
    .io_dmem_brupdate_b2_uop_exc_cause(lsu_io_dmem_brupdate_b2_uop_exc_cause),
    .io_dmem_brupdate_b2_uop_bypassable(lsu_io_dmem_brupdate_b2_uop_bypassable),
    .io_dmem_brupdate_b2_uop_mem_cmd(lsu_io_dmem_brupdate_b2_uop_mem_cmd),
    .io_dmem_brupdate_b2_uop_mem_size(lsu_io_dmem_brupdate_b2_uop_mem_size),
    .io_dmem_brupdate_b2_uop_mem_signed(lsu_io_dmem_brupdate_b2_uop_mem_signed),
    .io_dmem_brupdate_b2_uop_is_fence(lsu_io_dmem_brupdate_b2_uop_is_fence),
    .io_dmem_brupdate_b2_uop_is_fencei(lsu_io_dmem_brupdate_b2_uop_is_fencei),
    .io_dmem_brupdate_b2_uop_is_amo(lsu_io_dmem_brupdate_b2_uop_is_amo),
    .io_dmem_brupdate_b2_uop_uses_ldq(lsu_io_dmem_brupdate_b2_uop_uses_ldq),
    .io_dmem_brupdate_b2_uop_uses_stq(lsu_io_dmem_brupdate_b2_uop_uses_stq),
    .io_dmem_brupdate_b2_uop_is_sys_pc2epc(lsu_io_dmem_brupdate_b2_uop_is_sys_pc2epc),
    .io_dmem_brupdate_b2_uop_is_unique(lsu_io_dmem_brupdate_b2_uop_is_unique),
    .io_dmem_brupdate_b2_uop_flush_on_commit(lsu_io_dmem_brupdate_b2_uop_flush_on_commit),
    .io_dmem_brupdate_b2_uop_ldst_is_rs1(lsu_io_dmem_brupdate_b2_uop_ldst_is_rs1),
    .io_dmem_brupdate_b2_uop_ldst(lsu_io_dmem_brupdate_b2_uop_ldst),
    .io_dmem_brupdate_b2_uop_lrs1(lsu_io_dmem_brupdate_b2_uop_lrs1),
    .io_dmem_brupdate_b2_uop_lrs2(lsu_io_dmem_brupdate_b2_uop_lrs2),
    .io_dmem_brupdate_b2_uop_lrs3(lsu_io_dmem_brupdate_b2_uop_lrs3),
    .io_dmem_brupdate_b2_uop_ldst_val(lsu_io_dmem_brupdate_b2_uop_ldst_val),
    .io_dmem_brupdate_b2_uop_dst_rtype(lsu_io_dmem_brupdate_b2_uop_dst_rtype),
    .io_dmem_brupdate_b2_uop_lrs1_rtype(lsu_io_dmem_brupdate_b2_uop_lrs1_rtype),
    .io_dmem_brupdate_b2_uop_lrs2_rtype(lsu_io_dmem_brupdate_b2_uop_lrs2_rtype),
    .io_dmem_brupdate_b2_uop_frs3_en(lsu_io_dmem_brupdate_b2_uop_frs3_en),
    .io_dmem_brupdate_b2_uop_fp_val(lsu_io_dmem_brupdate_b2_uop_fp_val),
    .io_dmem_brupdate_b2_uop_fp_single(lsu_io_dmem_brupdate_b2_uop_fp_single),
    .io_dmem_brupdate_b2_uop_xcpt_pf_if(lsu_io_dmem_brupdate_b2_uop_xcpt_pf_if),
    .io_dmem_brupdate_b2_uop_xcpt_ae_if(lsu_io_dmem_brupdate_b2_uop_xcpt_ae_if),
    .io_dmem_brupdate_b2_uop_xcpt_ma_if(lsu_io_dmem_brupdate_b2_uop_xcpt_ma_if),
    .io_dmem_brupdate_b2_uop_bp_debug_if(lsu_io_dmem_brupdate_b2_uop_bp_debug_if),
    .io_dmem_brupdate_b2_uop_bp_xcpt_if(lsu_io_dmem_brupdate_b2_uop_bp_xcpt_if),
    .io_dmem_brupdate_b2_uop_debug_fsrc(lsu_io_dmem_brupdate_b2_uop_debug_fsrc),
    .io_dmem_brupdate_b2_uop_debug_tsrc(lsu_io_dmem_brupdate_b2_uop_debug_tsrc),
    .io_dmem_brupdate_b2_valid(lsu_io_dmem_brupdate_b2_valid),
    .io_dmem_brupdate_b2_mispredict(lsu_io_dmem_brupdate_b2_mispredict),
    .io_dmem_brupdate_b2_taken(lsu_io_dmem_brupdate_b2_taken),
    .io_dmem_brupdate_b2_cfi_type(lsu_io_dmem_brupdate_b2_cfi_type),
    .io_dmem_brupdate_b2_pc_sel(lsu_io_dmem_brupdate_b2_pc_sel),
    .io_dmem_brupdate_b2_jalr_target(lsu_io_dmem_brupdate_b2_jalr_target),
    .io_dmem_brupdate_b2_target_offset(lsu_io_dmem_brupdate_b2_target_offset),
    .io_dmem_exception(lsu_io_dmem_exception),
    .io_dmem_rob_pnr_idx(lsu_io_dmem_rob_pnr_idx),
    .io_dmem_rob_head_idx(lsu_io_dmem_rob_head_idx),
    .io_dmem_release_ready(lsu_io_dmem_release_ready),
    .io_dmem_release_valid(lsu_io_dmem_release_valid),
    .io_dmem_release_bits_opcode(lsu_io_dmem_release_bits_opcode),
    .io_dmem_release_bits_param(lsu_io_dmem_release_bits_param),
    .io_dmem_release_bits_size(lsu_io_dmem_release_bits_size),
    .io_dmem_release_bits_source(lsu_io_dmem_release_bits_source),
    .io_dmem_release_bits_address(lsu_io_dmem_release_bits_address),
    .io_dmem_release_bits_data(lsu_io_dmem_release_bits_data),
    .io_dmem_release_bits_corrupt(lsu_io_dmem_release_bits_corrupt),
    .io_dmem_force_order(lsu_io_dmem_force_order),
    .io_dmem_ordered(lsu_io_dmem_ordered),
    .io_dmem_perf_acquire(lsu_io_dmem_perf_acquire),
    .io_dmem_perf_release(lsu_io_dmem_perf_release),
    .io_hellacache_req_ready(lsu_io_hellacache_req_ready),
    .io_hellacache_req_valid(lsu_io_hellacache_req_valid),
    .io_hellacache_req_bits_addr(lsu_io_hellacache_req_bits_addr),
    .io_hellacache_req_bits_tag(lsu_io_hellacache_req_bits_tag),
    .io_hellacache_req_bits_cmd(lsu_io_hellacache_req_bits_cmd),
    .io_hellacache_req_bits_size(lsu_io_hellacache_req_bits_size),
    .io_hellacache_req_bits_signed(lsu_io_hellacache_req_bits_signed),
    .io_hellacache_req_bits_dprv(lsu_io_hellacache_req_bits_dprv),
    .io_hellacache_req_bits_phys(lsu_io_hellacache_req_bits_phys),
    .io_hellacache_req_bits_no_alloc(lsu_io_hellacache_req_bits_no_alloc),
    .io_hellacache_req_bits_no_xcpt(lsu_io_hellacache_req_bits_no_xcpt),
    .io_hellacache_req_bits_data(lsu_io_hellacache_req_bits_data),
    .io_hellacache_req_bits_mask(lsu_io_hellacache_req_bits_mask),
    .io_hellacache_s1_kill(lsu_io_hellacache_s1_kill),
    .io_hellacache_s1_data_data(lsu_io_hellacache_s1_data_data),
    .io_hellacache_s1_data_mask(lsu_io_hellacache_s1_data_mask),
    .io_hellacache_s2_nack(lsu_io_hellacache_s2_nack),
    .io_hellacache_s2_nack_cause_raw(lsu_io_hellacache_s2_nack_cause_raw),
    .io_hellacache_s2_kill(lsu_io_hellacache_s2_kill),
    .io_hellacache_s2_uncached(lsu_io_hellacache_s2_uncached),
    .io_hellacache_s2_paddr(lsu_io_hellacache_s2_paddr),
    .io_hellacache_resp_valid(lsu_io_hellacache_resp_valid),
    .io_hellacache_resp_bits_addr(lsu_io_hellacache_resp_bits_addr),
    .io_hellacache_resp_bits_tag(lsu_io_hellacache_resp_bits_tag),
    .io_hellacache_resp_bits_cmd(lsu_io_hellacache_resp_bits_cmd),
    .io_hellacache_resp_bits_size(lsu_io_hellacache_resp_bits_size),
    .io_hellacache_resp_bits_signed(lsu_io_hellacache_resp_bits_signed),
    .io_hellacache_resp_bits_dprv(lsu_io_hellacache_resp_bits_dprv),
    .io_hellacache_resp_bits_data(lsu_io_hellacache_resp_bits_data),
    .io_hellacache_resp_bits_mask(lsu_io_hellacache_resp_bits_mask),
    .io_hellacache_resp_bits_replay(lsu_io_hellacache_resp_bits_replay),
    .io_hellacache_resp_bits_has_data(lsu_io_hellacache_resp_bits_has_data),
    .io_hellacache_resp_bits_data_word_bypass(lsu_io_hellacache_resp_bits_data_word_bypass),
    .io_hellacache_resp_bits_data_raw(lsu_io_hellacache_resp_bits_data_raw),
    .io_hellacache_resp_bits_store_data(lsu_io_hellacache_resp_bits_store_data),
    .io_hellacache_replay_next(lsu_io_hellacache_replay_next),
    .io_hellacache_s2_xcpt_ma_ld(lsu_io_hellacache_s2_xcpt_ma_ld),
    .io_hellacache_s2_xcpt_ma_st(lsu_io_hellacache_s2_xcpt_ma_st),
    .io_hellacache_s2_xcpt_pf_ld(lsu_io_hellacache_s2_xcpt_pf_ld),
    .io_hellacache_s2_xcpt_pf_st(lsu_io_hellacache_s2_xcpt_pf_st),
    .io_hellacache_s2_xcpt_ae_ld(lsu_io_hellacache_s2_xcpt_ae_ld),
    .io_hellacache_s2_xcpt_ae_st(lsu_io_hellacache_s2_xcpt_ae_st),
    .io_hellacache_ordered(lsu_io_hellacache_ordered),
    .io_hellacache_perf_acquire(lsu_io_hellacache_perf_acquire),
    .io_hellacache_perf_release(lsu_io_hellacache_perf_release),
    .io_hellacache_perf_grant(lsu_io_hellacache_perf_grant),
    .io_hellacache_perf_tlbMiss(lsu_io_hellacache_perf_tlbMiss),
    .io_hellacache_perf_blocked(lsu_io_hellacache_perf_blocked),
    .io_hellacache_perf_canAcceptStoreThenLoad(lsu_io_hellacache_perf_canAcceptStoreThenLoad),
    .io_hellacache_perf_canAcceptStoreThenRMW(lsu_io_hellacache_perf_canAcceptStoreThenRMW),
    .io_hellacache_perf_canAcceptLoadThenLoad(lsu_io_hellacache_perf_canAcceptLoadThenLoad),
    .io_hellacache_perf_storeBufferEmptyAfterLoad(lsu_io_hellacache_perf_storeBufferEmptyAfterLoad),
    .io_hellacache_perf_storeBufferEmptyAfterStore(lsu_io_hellacache_perf_storeBufferEmptyAfterStore),
    .io_hellacache_keep_clock_enabled(lsu_io_hellacache_keep_clock_enabled),
    .io_hellacache_clock_enabled(lsu_io_hellacache_clock_enabled)
  );
  PTW ptw ( // @[tile.scala 230:20]
    .clock(ptw_clock),
    .reset(ptw_reset),
    .io_requestor_0_req_ready(ptw_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(ptw_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_valid(ptw_io_requestor_0_req_bits_valid),
    .io_requestor_0_req_bits_bits_addr(ptw_io_requestor_0_req_bits_bits_addr),
    .io_requestor_0_resp_valid(ptw_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_ae(ptw_io_requestor_0_resp_bits_ae),
    .io_requestor_0_resp_bits_pte_ppn(ptw_io_requestor_0_resp_bits_pte_ppn),
    .io_requestor_0_resp_bits_pte_reserved_for_software(ptw_io_requestor_0_resp_bits_pte_reserved_for_software),
    .io_requestor_0_resp_bits_pte_d(ptw_io_requestor_0_resp_bits_pte_d),
    .io_requestor_0_resp_bits_pte_a(ptw_io_requestor_0_resp_bits_pte_a),
    .io_requestor_0_resp_bits_pte_g(ptw_io_requestor_0_resp_bits_pte_g),
    .io_requestor_0_resp_bits_pte_u(ptw_io_requestor_0_resp_bits_pte_u),
    .io_requestor_0_resp_bits_pte_x(ptw_io_requestor_0_resp_bits_pte_x),
    .io_requestor_0_resp_bits_pte_w(ptw_io_requestor_0_resp_bits_pte_w),
    .io_requestor_0_resp_bits_pte_r(ptw_io_requestor_0_resp_bits_pte_r),
    .io_requestor_0_resp_bits_pte_v(ptw_io_requestor_0_resp_bits_pte_v),
    .io_requestor_0_resp_bits_level(ptw_io_requestor_0_resp_bits_level),
    .io_requestor_0_resp_bits_fragmented_superpage(ptw_io_requestor_0_resp_bits_fragmented_superpage),
    .io_requestor_0_resp_bits_homogeneous(ptw_io_requestor_0_resp_bits_homogeneous),
    .io_requestor_0_ptbr_mode(ptw_io_requestor_0_ptbr_mode),
    .io_requestor_0_ptbr_asid(ptw_io_requestor_0_ptbr_asid),
    .io_requestor_0_ptbr_ppn(ptw_io_requestor_0_ptbr_ppn),
    .io_requestor_0_status_debug(ptw_io_requestor_0_status_debug),
    .io_requestor_0_status_cease(ptw_io_requestor_0_status_cease),
    .io_requestor_0_status_wfi(ptw_io_requestor_0_status_wfi),
    .io_requestor_0_status_isa(ptw_io_requestor_0_status_isa),
    .io_requestor_0_status_dprv(ptw_io_requestor_0_status_dprv),
    .io_requestor_0_status_prv(ptw_io_requestor_0_status_prv),
    .io_requestor_0_status_sd(ptw_io_requestor_0_status_sd),
    .io_requestor_0_status_zero2(ptw_io_requestor_0_status_zero2),
    .io_requestor_0_status_sxl(ptw_io_requestor_0_status_sxl),
    .io_requestor_0_status_uxl(ptw_io_requestor_0_status_uxl),
    .io_requestor_0_status_sd_rv32(ptw_io_requestor_0_status_sd_rv32),
    .io_requestor_0_status_zero1(ptw_io_requestor_0_status_zero1),
    .io_requestor_0_status_tsr(ptw_io_requestor_0_status_tsr),
    .io_requestor_0_status_tw(ptw_io_requestor_0_status_tw),
    .io_requestor_0_status_tvm(ptw_io_requestor_0_status_tvm),
    .io_requestor_0_status_mxr(ptw_io_requestor_0_status_mxr),
    .io_requestor_0_status_sum(ptw_io_requestor_0_status_sum),
    .io_requestor_0_status_mprv(ptw_io_requestor_0_status_mprv),
    .io_requestor_0_status_xs(ptw_io_requestor_0_status_xs),
    .io_requestor_0_status_fs(ptw_io_requestor_0_status_fs),
    .io_requestor_0_status_mpp(ptw_io_requestor_0_status_mpp),
    .io_requestor_0_status_vs(ptw_io_requestor_0_status_vs),
    .io_requestor_0_status_spp(ptw_io_requestor_0_status_spp),
    .io_requestor_0_status_mpie(ptw_io_requestor_0_status_mpie),
    .io_requestor_0_status_hpie(ptw_io_requestor_0_status_hpie),
    .io_requestor_0_status_spie(ptw_io_requestor_0_status_spie),
    .io_requestor_0_status_upie(ptw_io_requestor_0_status_upie),
    .io_requestor_0_status_mie(ptw_io_requestor_0_status_mie),
    .io_requestor_0_status_hie(ptw_io_requestor_0_status_hie),
    .io_requestor_0_status_sie(ptw_io_requestor_0_status_sie),
    .io_requestor_0_status_uie(ptw_io_requestor_0_status_uie),
    .io_requestor_0_pmp_0_cfg_l(ptw_io_requestor_0_pmp_0_cfg_l),
    .io_requestor_0_pmp_0_cfg_res(ptw_io_requestor_0_pmp_0_cfg_res),
    .io_requestor_0_pmp_0_cfg_a(ptw_io_requestor_0_pmp_0_cfg_a),
    .io_requestor_0_pmp_0_cfg_x(ptw_io_requestor_0_pmp_0_cfg_x),
    .io_requestor_0_pmp_0_cfg_w(ptw_io_requestor_0_pmp_0_cfg_w),
    .io_requestor_0_pmp_0_cfg_r(ptw_io_requestor_0_pmp_0_cfg_r),
    .io_requestor_0_pmp_0_addr(ptw_io_requestor_0_pmp_0_addr),
    .io_requestor_0_pmp_0_mask(ptw_io_requestor_0_pmp_0_mask),
    .io_requestor_0_pmp_1_cfg_l(ptw_io_requestor_0_pmp_1_cfg_l),
    .io_requestor_0_pmp_1_cfg_res(ptw_io_requestor_0_pmp_1_cfg_res),
    .io_requestor_0_pmp_1_cfg_a(ptw_io_requestor_0_pmp_1_cfg_a),
    .io_requestor_0_pmp_1_cfg_x(ptw_io_requestor_0_pmp_1_cfg_x),
    .io_requestor_0_pmp_1_cfg_w(ptw_io_requestor_0_pmp_1_cfg_w),
    .io_requestor_0_pmp_1_cfg_r(ptw_io_requestor_0_pmp_1_cfg_r),
    .io_requestor_0_pmp_1_addr(ptw_io_requestor_0_pmp_1_addr),
    .io_requestor_0_pmp_1_mask(ptw_io_requestor_0_pmp_1_mask),
    .io_requestor_0_pmp_2_cfg_l(ptw_io_requestor_0_pmp_2_cfg_l),
    .io_requestor_0_pmp_2_cfg_res(ptw_io_requestor_0_pmp_2_cfg_res),
    .io_requestor_0_pmp_2_cfg_a(ptw_io_requestor_0_pmp_2_cfg_a),
    .io_requestor_0_pmp_2_cfg_x(ptw_io_requestor_0_pmp_2_cfg_x),
    .io_requestor_0_pmp_2_cfg_w(ptw_io_requestor_0_pmp_2_cfg_w),
    .io_requestor_0_pmp_2_cfg_r(ptw_io_requestor_0_pmp_2_cfg_r),
    .io_requestor_0_pmp_2_addr(ptw_io_requestor_0_pmp_2_addr),
    .io_requestor_0_pmp_2_mask(ptw_io_requestor_0_pmp_2_mask),
    .io_requestor_0_pmp_3_cfg_l(ptw_io_requestor_0_pmp_3_cfg_l),
    .io_requestor_0_pmp_3_cfg_res(ptw_io_requestor_0_pmp_3_cfg_res),
    .io_requestor_0_pmp_3_cfg_a(ptw_io_requestor_0_pmp_3_cfg_a),
    .io_requestor_0_pmp_3_cfg_x(ptw_io_requestor_0_pmp_3_cfg_x),
    .io_requestor_0_pmp_3_cfg_w(ptw_io_requestor_0_pmp_3_cfg_w),
    .io_requestor_0_pmp_3_cfg_r(ptw_io_requestor_0_pmp_3_cfg_r),
    .io_requestor_0_pmp_3_addr(ptw_io_requestor_0_pmp_3_addr),
    .io_requestor_0_pmp_3_mask(ptw_io_requestor_0_pmp_3_mask),
    .io_requestor_0_pmp_4_cfg_l(ptw_io_requestor_0_pmp_4_cfg_l),
    .io_requestor_0_pmp_4_cfg_res(ptw_io_requestor_0_pmp_4_cfg_res),
    .io_requestor_0_pmp_4_cfg_a(ptw_io_requestor_0_pmp_4_cfg_a),
    .io_requestor_0_pmp_4_cfg_x(ptw_io_requestor_0_pmp_4_cfg_x),
    .io_requestor_0_pmp_4_cfg_w(ptw_io_requestor_0_pmp_4_cfg_w),
    .io_requestor_0_pmp_4_cfg_r(ptw_io_requestor_0_pmp_4_cfg_r),
    .io_requestor_0_pmp_4_addr(ptw_io_requestor_0_pmp_4_addr),
    .io_requestor_0_pmp_4_mask(ptw_io_requestor_0_pmp_4_mask),
    .io_requestor_0_pmp_5_cfg_l(ptw_io_requestor_0_pmp_5_cfg_l),
    .io_requestor_0_pmp_5_cfg_res(ptw_io_requestor_0_pmp_5_cfg_res),
    .io_requestor_0_pmp_5_cfg_a(ptw_io_requestor_0_pmp_5_cfg_a),
    .io_requestor_0_pmp_5_cfg_x(ptw_io_requestor_0_pmp_5_cfg_x),
    .io_requestor_0_pmp_5_cfg_w(ptw_io_requestor_0_pmp_5_cfg_w),
    .io_requestor_0_pmp_5_cfg_r(ptw_io_requestor_0_pmp_5_cfg_r),
    .io_requestor_0_pmp_5_addr(ptw_io_requestor_0_pmp_5_addr),
    .io_requestor_0_pmp_5_mask(ptw_io_requestor_0_pmp_5_mask),
    .io_requestor_0_pmp_6_cfg_l(ptw_io_requestor_0_pmp_6_cfg_l),
    .io_requestor_0_pmp_6_cfg_res(ptw_io_requestor_0_pmp_6_cfg_res),
    .io_requestor_0_pmp_6_cfg_a(ptw_io_requestor_0_pmp_6_cfg_a),
    .io_requestor_0_pmp_6_cfg_x(ptw_io_requestor_0_pmp_6_cfg_x),
    .io_requestor_0_pmp_6_cfg_w(ptw_io_requestor_0_pmp_6_cfg_w),
    .io_requestor_0_pmp_6_cfg_r(ptw_io_requestor_0_pmp_6_cfg_r),
    .io_requestor_0_pmp_6_addr(ptw_io_requestor_0_pmp_6_addr),
    .io_requestor_0_pmp_6_mask(ptw_io_requestor_0_pmp_6_mask),
    .io_requestor_0_pmp_7_cfg_l(ptw_io_requestor_0_pmp_7_cfg_l),
    .io_requestor_0_pmp_7_cfg_res(ptw_io_requestor_0_pmp_7_cfg_res),
    .io_requestor_0_pmp_7_cfg_a(ptw_io_requestor_0_pmp_7_cfg_a),
    .io_requestor_0_pmp_7_cfg_x(ptw_io_requestor_0_pmp_7_cfg_x),
    .io_requestor_0_pmp_7_cfg_w(ptw_io_requestor_0_pmp_7_cfg_w),
    .io_requestor_0_pmp_7_cfg_r(ptw_io_requestor_0_pmp_7_cfg_r),
    .io_requestor_0_pmp_7_addr(ptw_io_requestor_0_pmp_7_addr),
    .io_requestor_0_pmp_7_mask(ptw_io_requestor_0_pmp_7_mask),
    .io_requestor_0_customCSRs_csrs_0_wen(ptw_io_requestor_0_customCSRs_csrs_0_wen),
    .io_requestor_0_customCSRs_csrs_0_wdata(ptw_io_requestor_0_customCSRs_csrs_0_wdata),
    .io_requestor_0_customCSRs_csrs_0_value(ptw_io_requestor_0_customCSRs_csrs_0_value),
    .io_requestor_1_req_ready(ptw_io_requestor_1_req_ready),
    .io_requestor_1_req_valid(ptw_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_valid(ptw_io_requestor_1_req_bits_valid),
    .io_requestor_1_req_bits_bits_addr(ptw_io_requestor_1_req_bits_bits_addr),
    .io_requestor_1_resp_valid(ptw_io_requestor_1_resp_valid),
    .io_requestor_1_resp_bits_ae(ptw_io_requestor_1_resp_bits_ae),
    .io_requestor_1_resp_bits_pte_ppn(ptw_io_requestor_1_resp_bits_pte_ppn),
    .io_requestor_1_resp_bits_pte_reserved_for_software(ptw_io_requestor_1_resp_bits_pte_reserved_for_software),
    .io_requestor_1_resp_bits_pte_d(ptw_io_requestor_1_resp_bits_pte_d),
    .io_requestor_1_resp_bits_pte_a(ptw_io_requestor_1_resp_bits_pte_a),
    .io_requestor_1_resp_bits_pte_g(ptw_io_requestor_1_resp_bits_pte_g),
    .io_requestor_1_resp_bits_pte_u(ptw_io_requestor_1_resp_bits_pte_u),
    .io_requestor_1_resp_bits_pte_x(ptw_io_requestor_1_resp_bits_pte_x),
    .io_requestor_1_resp_bits_pte_w(ptw_io_requestor_1_resp_bits_pte_w),
    .io_requestor_1_resp_bits_pte_r(ptw_io_requestor_1_resp_bits_pte_r),
    .io_requestor_1_resp_bits_pte_v(ptw_io_requestor_1_resp_bits_pte_v),
    .io_requestor_1_resp_bits_level(ptw_io_requestor_1_resp_bits_level),
    .io_requestor_1_resp_bits_fragmented_superpage(ptw_io_requestor_1_resp_bits_fragmented_superpage),
    .io_requestor_1_resp_bits_homogeneous(ptw_io_requestor_1_resp_bits_homogeneous),
    .io_requestor_1_ptbr_mode(ptw_io_requestor_1_ptbr_mode),
    .io_requestor_1_ptbr_asid(ptw_io_requestor_1_ptbr_asid),
    .io_requestor_1_ptbr_ppn(ptw_io_requestor_1_ptbr_ppn),
    .io_requestor_1_status_debug(ptw_io_requestor_1_status_debug),
    .io_requestor_1_status_cease(ptw_io_requestor_1_status_cease),
    .io_requestor_1_status_wfi(ptw_io_requestor_1_status_wfi),
    .io_requestor_1_status_isa(ptw_io_requestor_1_status_isa),
    .io_requestor_1_status_dprv(ptw_io_requestor_1_status_dprv),
    .io_requestor_1_status_prv(ptw_io_requestor_1_status_prv),
    .io_requestor_1_status_sd(ptw_io_requestor_1_status_sd),
    .io_requestor_1_status_zero2(ptw_io_requestor_1_status_zero2),
    .io_requestor_1_status_sxl(ptw_io_requestor_1_status_sxl),
    .io_requestor_1_status_uxl(ptw_io_requestor_1_status_uxl),
    .io_requestor_1_status_sd_rv32(ptw_io_requestor_1_status_sd_rv32),
    .io_requestor_1_status_zero1(ptw_io_requestor_1_status_zero1),
    .io_requestor_1_status_tsr(ptw_io_requestor_1_status_tsr),
    .io_requestor_1_status_tw(ptw_io_requestor_1_status_tw),
    .io_requestor_1_status_tvm(ptw_io_requestor_1_status_tvm),
    .io_requestor_1_status_mxr(ptw_io_requestor_1_status_mxr),
    .io_requestor_1_status_sum(ptw_io_requestor_1_status_sum),
    .io_requestor_1_status_mprv(ptw_io_requestor_1_status_mprv),
    .io_requestor_1_status_xs(ptw_io_requestor_1_status_xs),
    .io_requestor_1_status_fs(ptw_io_requestor_1_status_fs),
    .io_requestor_1_status_mpp(ptw_io_requestor_1_status_mpp),
    .io_requestor_1_status_vs(ptw_io_requestor_1_status_vs),
    .io_requestor_1_status_spp(ptw_io_requestor_1_status_spp),
    .io_requestor_1_status_mpie(ptw_io_requestor_1_status_mpie),
    .io_requestor_1_status_hpie(ptw_io_requestor_1_status_hpie),
    .io_requestor_1_status_spie(ptw_io_requestor_1_status_spie),
    .io_requestor_1_status_upie(ptw_io_requestor_1_status_upie),
    .io_requestor_1_status_mie(ptw_io_requestor_1_status_mie),
    .io_requestor_1_status_hie(ptw_io_requestor_1_status_hie),
    .io_requestor_1_status_sie(ptw_io_requestor_1_status_sie),
    .io_requestor_1_status_uie(ptw_io_requestor_1_status_uie),
    .io_requestor_1_pmp_0_cfg_l(ptw_io_requestor_1_pmp_0_cfg_l),
    .io_requestor_1_pmp_0_cfg_res(ptw_io_requestor_1_pmp_0_cfg_res),
    .io_requestor_1_pmp_0_cfg_a(ptw_io_requestor_1_pmp_0_cfg_a),
    .io_requestor_1_pmp_0_cfg_x(ptw_io_requestor_1_pmp_0_cfg_x),
    .io_requestor_1_pmp_0_cfg_w(ptw_io_requestor_1_pmp_0_cfg_w),
    .io_requestor_1_pmp_0_cfg_r(ptw_io_requestor_1_pmp_0_cfg_r),
    .io_requestor_1_pmp_0_addr(ptw_io_requestor_1_pmp_0_addr),
    .io_requestor_1_pmp_0_mask(ptw_io_requestor_1_pmp_0_mask),
    .io_requestor_1_pmp_1_cfg_l(ptw_io_requestor_1_pmp_1_cfg_l),
    .io_requestor_1_pmp_1_cfg_res(ptw_io_requestor_1_pmp_1_cfg_res),
    .io_requestor_1_pmp_1_cfg_a(ptw_io_requestor_1_pmp_1_cfg_a),
    .io_requestor_1_pmp_1_cfg_x(ptw_io_requestor_1_pmp_1_cfg_x),
    .io_requestor_1_pmp_1_cfg_w(ptw_io_requestor_1_pmp_1_cfg_w),
    .io_requestor_1_pmp_1_cfg_r(ptw_io_requestor_1_pmp_1_cfg_r),
    .io_requestor_1_pmp_1_addr(ptw_io_requestor_1_pmp_1_addr),
    .io_requestor_1_pmp_1_mask(ptw_io_requestor_1_pmp_1_mask),
    .io_requestor_1_pmp_2_cfg_l(ptw_io_requestor_1_pmp_2_cfg_l),
    .io_requestor_1_pmp_2_cfg_res(ptw_io_requestor_1_pmp_2_cfg_res),
    .io_requestor_1_pmp_2_cfg_a(ptw_io_requestor_1_pmp_2_cfg_a),
    .io_requestor_1_pmp_2_cfg_x(ptw_io_requestor_1_pmp_2_cfg_x),
    .io_requestor_1_pmp_2_cfg_w(ptw_io_requestor_1_pmp_2_cfg_w),
    .io_requestor_1_pmp_2_cfg_r(ptw_io_requestor_1_pmp_2_cfg_r),
    .io_requestor_1_pmp_2_addr(ptw_io_requestor_1_pmp_2_addr),
    .io_requestor_1_pmp_2_mask(ptw_io_requestor_1_pmp_2_mask),
    .io_requestor_1_pmp_3_cfg_l(ptw_io_requestor_1_pmp_3_cfg_l),
    .io_requestor_1_pmp_3_cfg_res(ptw_io_requestor_1_pmp_3_cfg_res),
    .io_requestor_1_pmp_3_cfg_a(ptw_io_requestor_1_pmp_3_cfg_a),
    .io_requestor_1_pmp_3_cfg_x(ptw_io_requestor_1_pmp_3_cfg_x),
    .io_requestor_1_pmp_3_cfg_w(ptw_io_requestor_1_pmp_3_cfg_w),
    .io_requestor_1_pmp_3_cfg_r(ptw_io_requestor_1_pmp_3_cfg_r),
    .io_requestor_1_pmp_3_addr(ptw_io_requestor_1_pmp_3_addr),
    .io_requestor_1_pmp_3_mask(ptw_io_requestor_1_pmp_3_mask),
    .io_requestor_1_pmp_4_cfg_l(ptw_io_requestor_1_pmp_4_cfg_l),
    .io_requestor_1_pmp_4_cfg_res(ptw_io_requestor_1_pmp_4_cfg_res),
    .io_requestor_1_pmp_4_cfg_a(ptw_io_requestor_1_pmp_4_cfg_a),
    .io_requestor_1_pmp_4_cfg_x(ptw_io_requestor_1_pmp_4_cfg_x),
    .io_requestor_1_pmp_4_cfg_w(ptw_io_requestor_1_pmp_4_cfg_w),
    .io_requestor_1_pmp_4_cfg_r(ptw_io_requestor_1_pmp_4_cfg_r),
    .io_requestor_1_pmp_4_addr(ptw_io_requestor_1_pmp_4_addr),
    .io_requestor_1_pmp_4_mask(ptw_io_requestor_1_pmp_4_mask),
    .io_requestor_1_pmp_5_cfg_l(ptw_io_requestor_1_pmp_5_cfg_l),
    .io_requestor_1_pmp_5_cfg_res(ptw_io_requestor_1_pmp_5_cfg_res),
    .io_requestor_1_pmp_5_cfg_a(ptw_io_requestor_1_pmp_5_cfg_a),
    .io_requestor_1_pmp_5_cfg_x(ptw_io_requestor_1_pmp_5_cfg_x),
    .io_requestor_1_pmp_5_cfg_w(ptw_io_requestor_1_pmp_5_cfg_w),
    .io_requestor_1_pmp_5_cfg_r(ptw_io_requestor_1_pmp_5_cfg_r),
    .io_requestor_1_pmp_5_addr(ptw_io_requestor_1_pmp_5_addr),
    .io_requestor_1_pmp_5_mask(ptw_io_requestor_1_pmp_5_mask),
    .io_requestor_1_pmp_6_cfg_l(ptw_io_requestor_1_pmp_6_cfg_l),
    .io_requestor_1_pmp_6_cfg_res(ptw_io_requestor_1_pmp_6_cfg_res),
    .io_requestor_1_pmp_6_cfg_a(ptw_io_requestor_1_pmp_6_cfg_a),
    .io_requestor_1_pmp_6_cfg_x(ptw_io_requestor_1_pmp_6_cfg_x),
    .io_requestor_1_pmp_6_cfg_w(ptw_io_requestor_1_pmp_6_cfg_w),
    .io_requestor_1_pmp_6_cfg_r(ptw_io_requestor_1_pmp_6_cfg_r),
    .io_requestor_1_pmp_6_addr(ptw_io_requestor_1_pmp_6_addr),
    .io_requestor_1_pmp_6_mask(ptw_io_requestor_1_pmp_6_mask),
    .io_requestor_1_pmp_7_cfg_l(ptw_io_requestor_1_pmp_7_cfg_l),
    .io_requestor_1_pmp_7_cfg_res(ptw_io_requestor_1_pmp_7_cfg_res),
    .io_requestor_1_pmp_7_cfg_a(ptw_io_requestor_1_pmp_7_cfg_a),
    .io_requestor_1_pmp_7_cfg_x(ptw_io_requestor_1_pmp_7_cfg_x),
    .io_requestor_1_pmp_7_cfg_w(ptw_io_requestor_1_pmp_7_cfg_w),
    .io_requestor_1_pmp_7_cfg_r(ptw_io_requestor_1_pmp_7_cfg_r),
    .io_requestor_1_pmp_7_addr(ptw_io_requestor_1_pmp_7_addr),
    .io_requestor_1_pmp_7_mask(ptw_io_requestor_1_pmp_7_mask),
    .io_requestor_1_customCSRs_csrs_0_wen(ptw_io_requestor_1_customCSRs_csrs_0_wen),
    .io_requestor_1_customCSRs_csrs_0_wdata(ptw_io_requestor_1_customCSRs_csrs_0_wdata),
    .io_requestor_1_customCSRs_csrs_0_value(ptw_io_requestor_1_customCSRs_csrs_0_value),
    .io_requestor_2_req_ready(ptw_io_requestor_2_req_ready),
    .io_requestor_2_req_valid(ptw_io_requestor_2_req_valid),
    .io_requestor_2_req_bits_valid(ptw_io_requestor_2_req_bits_valid),
    .io_requestor_2_req_bits_bits_addr(ptw_io_requestor_2_req_bits_bits_addr),
    .io_requestor_2_resp_valid(ptw_io_requestor_2_resp_valid),
    .io_requestor_2_resp_bits_ae(ptw_io_requestor_2_resp_bits_ae),
    .io_requestor_2_resp_bits_pte_ppn(ptw_io_requestor_2_resp_bits_pte_ppn),
    .io_requestor_2_resp_bits_pte_reserved_for_software(ptw_io_requestor_2_resp_bits_pte_reserved_for_software),
    .io_requestor_2_resp_bits_pte_d(ptw_io_requestor_2_resp_bits_pte_d),
    .io_requestor_2_resp_bits_pte_a(ptw_io_requestor_2_resp_bits_pte_a),
    .io_requestor_2_resp_bits_pte_g(ptw_io_requestor_2_resp_bits_pte_g),
    .io_requestor_2_resp_bits_pte_u(ptw_io_requestor_2_resp_bits_pte_u),
    .io_requestor_2_resp_bits_pte_x(ptw_io_requestor_2_resp_bits_pte_x),
    .io_requestor_2_resp_bits_pte_w(ptw_io_requestor_2_resp_bits_pte_w),
    .io_requestor_2_resp_bits_pte_r(ptw_io_requestor_2_resp_bits_pte_r),
    .io_requestor_2_resp_bits_pte_v(ptw_io_requestor_2_resp_bits_pte_v),
    .io_requestor_2_resp_bits_level(ptw_io_requestor_2_resp_bits_level),
    .io_requestor_2_resp_bits_fragmented_superpage(ptw_io_requestor_2_resp_bits_fragmented_superpage),
    .io_requestor_2_resp_bits_homogeneous(ptw_io_requestor_2_resp_bits_homogeneous),
    .io_requestor_2_ptbr_mode(ptw_io_requestor_2_ptbr_mode),
    .io_requestor_2_ptbr_asid(ptw_io_requestor_2_ptbr_asid),
    .io_requestor_2_ptbr_ppn(ptw_io_requestor_2_ptbr_ppn),
    .io_requestor_2_status_debug(ptw_io_requestor_2_status_debug),
    .io_requestor_2_status_cease(ptw_io_requestor_2_status_cease),
    .io_requestor_2_status_wfi(ptw_io_requestor_2_status_wfi),
    .io_requestor_2_status_isa(ptw_io_requestor_2_status_isa),
    .io_requestor_2_status_dprv(ptw_io_requestor_2_status_dprv),
    .io_requestor_2_status_prv(ptw_io_requestor_2_status_prv),
    .io_requestor_2_status_sd(ptw_io_requestor_2_status_sd),
    .io_requestor_2_status_zero2(ptw_io_requestor_2_status_zero2),
    .io_requestor_2_status_sxl(ptw_io_requestor_2_status_sxl),
    .io_requestor_2_status_uxl(ptw_io_requestor_2_status_uxl),
    .io_requestor_2_status_sd_rv32(ptw_io_requestor_2_status_sd_rv32),
    .io_requestor_2_status_zero1(ptw_io_requestor_2_status_zero1),
    .io_requestor_2_status_tsr(ptw_io_requestor_2_status_tsr),
    .io_requestor_2_status_tw(ptw_io_requestor_2_status_tw),
    .io_requestor_2_status_tvm(ptw_io_requestor_2_status_tvm),
    .io_requestor_2_status_mxr(ptw_io_requestor_2_status_mxr),
    .io_requestor_2_status_sum(ptw_io_requestor_2_status_sum),
    .io_requestor_2_status_mprv(ptw_io_requestor_2_status_mprv),
    .io_requestor_2_status_xs(ptw_io_requestor_2_status_xs),
    .io_requestor_2_status_fs(ptw_io_requestor_2_status_fs),
    .io_requestor_2_status_mpp(ptw_io_requestor_2_status_mpp),
    .io_requestor_2_status_vs(ptw_io_requestor_2_status_vs),
    .io_requestor_2_status_spp(ptw_io_requestor_2_status_spp),
    .io_requestor_2_status_mpie(ptw_io_requestor_2_status_mpie),
    .io_requestor_2_status_hpie(ptw_io_requestor_2_status_hpie),
    .io_requestor_2_status_spie(ptw_io_requestor_2_status_spie),
    .io_requestor_2_status_upie(ptw_io_requestor_2_status_upie),
    .io_requestor_2_status_mie(ptw_io_requestor_2_status_mie),
    .io_requestor_2_status_hie(ptw_io_requestor_2_status_hie),
    .io_requestor_2_status_sie(ptw_io_requestor_2_status_sie),
    .io_requestor_2_status_uie(ptw_io_requestor_2_status_uie),
    .io_requestor_2_pmp_0_cfg_l(ptw_io_requestor_2_pmp_0_cfg_l),
    .io_requestor_2_pmp_0_cfg_res(ptw_io_requestor_2_pmp_0_cfg_res),
    .io_requestor_2_pmp_0_cfg_a(ptw_io_requestor_2_pmp_0_cfg_a),
    .io_requestor_2_pmp_0_cfg_x(ptw_io_requestor_2_pmp_0_cfg_x),
    .io_requestor_2_pmp_0_cfg_w(ptw_io_requestor_2_pmp_0_cfg_w),
    .io_requestor_2_pmp_0_cfg_r(ptw_io_requestor_2_pmp_0_cfg_r),
    .io_requestor_2_pmp_0_addr(ptw_io_requestor_2_pmp_0_addr),
    .io_requestor_2_pmp_0_mask(ptw_io_requestor_2_pmp_0_mask),
    .io_requestor_2_pmp_1_cfg_l(ptw_io_requestor_2_pmp_1_cfg_l),
    .io_requestor_2_pmp_1_cfg_res(ptw_io_requestor_2_pmp_1_cfg_res),
    .io_requestor_2_pmp_1_cfg_a(ptw_io_requestor_2_pmp_1_cfg_a),
    .io_requestor_2_pmp_1_cfg_x(ptw_io_requestor_2_pmp_1_cfg_x),
    .io_requestor_2_pmp_1_cfg_w(ptw_io_requestor_2_pmp_1_cfg_w),
    .io_requestor_2_pmp_1_cfg_r(ptw_io_requestor_2_pmp_1_cfg_r),
    .io_requestor_2_pmp_1_addr(ptw_io_requestor_2_pmp_1_addr),
    .io_requestor_2_pmp_1_mask(ptw_io_requestor_2_pmp_1_mask),
    .io_requestor_2_pmp_2_cfg_l(ptw_io_requestor_2_pmp_2_cfg_l),
    .io_requestor_2_pmp_2_cfg_res(ptw_io_requestor_2_pmp_2_cfg_res),
    .io_requestor_2_pmp_2_cfg_a(ptw_io_requestor_2_pmp_2_cfg_a),
    .io_requestor_2_pmp_2_cfg_x(ptw_io_requestor_2_pmp_2_cfg_x),
    .io_requestor_2_pmp_2_cfg_w(ptw_io_requestor_2_pmp_2_cfg_w),
    .io_requestor_2_pmp_2_cfg_r(ptw_io_requestor_2_pmp_2_cfg_r),
    .io_requestor_2_pmp_2_addr(ptw_io_requestor_2_pmp_2_addr),
    .io_requestor_2_pmp_2_mask(ptw_io_requestor_2_pmp_2_mask),
    .io_requestor_2_pmp_3_cfg_l(ptw_io_requestor_2_pmp_3_cfg_l),
    .io_requestor_2_pmp_3_cfg_res(ptw_io_requestor_2_pmp_3_cfg_res),
    .io_requestor_2_pmp_3_cfg_a(ptw_io_requestor_2_pmp_3_cfg_a),
    .io_requestor_2_pmp_3_cfg_x(ptw_io_requestor_2_pmp_3_cfg_x),
    .io_requestor_2_pmp_3_cfg_w(ptw_io_requestor_2_pmp_3_cfg_w),
    .io_requestor_2_pmp_3_cfg_r(ptw_io_requestor_2_pmp_3_cfg_r),
    .io_requestor_2_pmp_3_addr(ptw_io_requestor_2_pmp_3_addr),
    .io_requestor_2_pmp_3_mask(ptw_io_requestor_2_pmp_3_mask),
    .io_requestor_2_pmp_4_cfg_l(ptw_io_requestor_2_pmp_4_cfg_l),
    .io_requestor_2_pmp_4_cfg_res(ptw_io_requestor_2_pmp_4_cfg_res),
    .io_requestor_2_pmp_4_cfg_a(ptw_io_requestor_2_pmp_4_cfg_a),
    .io_requestor_2_pmp_4_cfg_x(ptw_io_requestor_2_pmp_4_cfg_x),
    .io_requestor_2_pmp_4_cfg_w(ptw_io_requestor_2_pmp_4_cfg_w),
    .io_requestor_2_pmp_4_cfg_r(ptw_io_requestor_2_pmp_4_cfg_r),
    .io_requestor_2_pmp_4_addr(ptw_io_requestor_2_pmp_4_addr),
    .io_requestor_2_pmp_4_mask(ptw_io_requestor_2_pmp_4_mask),
    .io_requestor_2_pmp_5_cfg_l(ptw_io_requestor_2_pmp_5_cfg_l),
    .io_requestor_2_pmp_5_cfg_res(ptw_io_requestor_2_pmp_5_cfg_res),
    .io_requestor_2_pmp_5_cfg_a(ptw_io_requestor_2_pmp_5_cfg_a),
    .io_requestor_2_pmp_5_cfg_x(ptw_io_requestor_2_pmp_5_cfg_x),
    .io_requestor_2_pmp_5_cfg_w(ptw_io_requestor_2_pmp_5_cfg_w),
    .io_requestor_2_pmp_5_cfg_r(ptw_io_requestor_2_pmp_5_cfg_r),
    .io_requestor_2_pmp_5_addr(ptw_io_requestor_2_pmp_5_addr),
    .io_requestor_2_pmp_5_mask(ptw_io_requestor_2_pmp_5_mask),
    .io_requestor_2_pmp_6_cfg_l(ptw_io_requestor_2_pmp_6_cfg_l),
    .io_requestor_2_pmp_6_cfg_res(ptw_io_requestor_2_pmp_6_cfg_res),
    .io_requestor_2_pmp_6_cfg_a(ptw_io_requestor_2_pmp_6_cfg_a),
    .io_requestor_2_pmp_6_cfg_x(ptw_io_requestor_2_pmp_6_cfg_x),
    .io_requestor_2_pmp_6_cfg_w(ptw_io_requestor_2_pmp_6_cfg_w),
    .io_requestor_2_pmp_6_cfg_r(ptw_io_requestor_2_pmp_6_cfg_r),
    .io_requestor_2_pmp_6_addr(ptw_io_requestor_2_pmp_6_addr),
    .io_requestor_2_pmp_6_mask(ptw_io_requestor_2_pmp_6_mask),
    .io_requestor_2_pmp_7_cfg_l(ptw_io_requestor_2_pmp_7_cfg_l),
    .io_requestor_2_pmp_7_cfg_res(ptw_io_requestor_2_pmp_7_cfg_res),
    .io_requestor_2_pmp_7_cfg_a(ptw_io_requestor_2_pmp_7_cfg_a),
    .io_requestor_2_pmp_7_cfg_x(ptw_io_requestor_2_pmp_7_cfg_x),
    .io_requestor_2_pmp_7_cfg_w(ptw_io_requestor_2_pmp_7_cfg_w),
    .io_requestor_2_pmp_7_cfg_r(ptw_io_requestor_2_pmp_7_cfg_r),
    .io_requestor_2_pmp_7_addr(ptw_io_requestor_2_pmp_7_addr),
    .io_requestor_2_pmp_7_mask(ptw_io_requestor_2_pmp_7_mask),
    .io_requestor_2_customCSRs_csrs_0_wen(ptw_io_requestor_2_customCSRs_csrs_0_wen),
    .io_requestor_2_customCSRs_csrs_0_wdata(ptw_io_requestor_2_customCSRs_csrs_0_wdata),
    .io_requestor_2_customCSRs_csrs_0_value(ptw_io_requestor_2_customCSRs_csrs_0_value),
    .io_mem_req_ready(ptw_io_mem_req_ready),
    .io_mem_req_valid(ptw_io_mem_req_valid),
    .io_mem_req_bits_addr(ptw_io_mem_req_bits_addr),
    .io_mem_req_bits_tag(ptw_io_mem_req_bits_tag),
    .io_mem_req_bits_cmd(ptw_io_mem_req_bits_cmd),
    .io_mem_req_bits_size(ptw_io_mem_req_bits_size),
    .io_mem_req_bits_signed(ptw_io_mem_req_bits_signed),
    .io_mem_req_bits_dprv(ptw_io_mem_req_bits_dprv),
    .io_mem_req_bits_phys(ptw_io_mem_req_bits_phys),
    .io_mem_req_bits_no_alloc(ptw_io_mem_req_bits_no_alloc),
    .io_mem_req_bits_no_xcpt(ptw_io_mem_req_bits_no_xcpt),
    .io_mem_req_bits_data(ptw_io_mem_req_bits_data),
    .io_mem_req_bits_mask(ptw_io_mem_req_bits_mask),
    .io_mem_s1_kill(ptw_io_mem_s1_kill),
    .io_mem_s1_data_data(ptw_io_mem_s1_data_data),
    .io_mem_s1_data_mask(ptw_io_mem_s1_data_mask),
    .io_mem_s2_nack(ptw_io_mem_s2_nack),
    .io_mem_s2_nack_cause_raw(ptw_io_mem_s2_nack_cause_raw),
    .io_mem_s2_kill(ptw_io_mem_s2_kill),
    .io_mem_s2_uncached(ptw_io_mem_s2_uncached),
    .io_mem_s2_paddr(ptw_io_mem_s2_paddr),
    .io_mem_resp_valid(ptw_io_mem_resp_valid),
    .io_mem_resp_bits_addr(ptw_io_mem_resp_bits_addr),
    .io_mem_resp_bits_tag(ptw_io_mem_resp_bits_tag),
    .io_mem_resp_bits_cmd(ptw_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_size(ptw_io_mem_resp_bits_size),
    .io_mem_resp_bits_signed(ptw_io_mem_resp_bits_signed),
    .io_mem_resp_bits_dprv(ptw_io_mem_resp_bits_dprv),
    .io_mem_resp_bits_data(ptw_io_mem_resp_bits_data),
    .io_mem_resp_bits_mask(ptw_io_mem_resp_bits_mask),
    .io_mem_resp_bits_replay(ptw_io_mem_resp_bits_replay),
    .io_mem_resp_bits_has_data(ptw_io_mem_resp_bits_has_data),
    .io_mem_resp_bits_data_word_bypass(ptw_io_mem_resp_bits_data_word_bypass),
    .io_mem_resp_bits_data_raw(ptw_io_mem_resp_bits_data_raw),
    .io_mem_resp_bits_store_data(ptw_io_mem_resp_bits_store_data),
    .io_mem_replay_next(ptw_io_mem_replay_next),
    .io_mem_s2_xcpt_ma_ld(ptw_io_mem_s2_xcpt_ma_ld),
    .io_mem_s2_xcpt_ma_st(ptw_io_mem_s2_xcpt_ma_st),
    .io_mem_s2_xcpt_pf_ld(ptw_io_mem_s2_xcpt_pf_ld),
    .io_mem_s2_xcpt_pf_st(ptw_io_mem_s2_xcpt_pf_st),
    .io_mem_s2_xcpt_ae_ld(ptw_io_mem_s2_xcpt_ae_ld),
    .io_mem_s2_xcpt_ae_st(ptw_io_mem_s2_xcpt_ae_st),
    .io_mem_ordered(ptw_io_mem_ordered),
    .io_mem_perf_acquire(ptw_io_mem_perf_acquire),
    .io_mem_perf_release(ptw_io_mem_perf_release),
    .io_mem_perf_grant(ptw_io_mem_perf_grant),
    .io_mem_perf_tlbMiss(ptw_io_mem_perf_tlbMiss),
    .io_mem_perf_blocked(ptw_io_mem_perf_blocked),
    .io_mem_perf_canAcceptStoreThenLoad(ptw_io_mem_perf_canAcceptStoreThenLoad),
    .io_mem_perf_canAcceptStoreThenRMW(ptw_io_mem_perf_canAcceptStoreThenRMW),
    .io_mem_perf_canAcceptLoadThenLoad(ptw_io_mem_perf_canAcceptLoadThenLoad),
    .io_mem_perf_storeBufferEmptyAfterLoad(ptw_io_mem_perf_storeBufferEmptyAfterLoad),
    .io_mem_perf_storeBufferEmptyAfterStore(ptw_io_mem_perf_storeBufferEmptyAfterStore),
    .io_mem_keep_clock_enabled(ptw_io_mem_keep_clock_enabled),
    .io_mem_clock_enabled(ptw_io_mem_clock_enabled),
    .io_dpath_ptbr_mode(ptw_io_dpath_ptbr_mode),
    .io_dpath_ptbr_asid(ptw_io_dpath_ptbr_asid),
    .io_dpath_ptbr_ppn(ptw_io_dpath_ptbr_ppn),
    .io_dpath_sfence_valid(ptw_io_dpath_sfence_valid),
    .io_dpath_sfence_bits_rs1(ptw_io_dpath_sfence_bits_rs1),
    .io_dpath_sfence_bits_rs2(ptw_io_dpath_sfence_bits_rs2),
    .io_dpath_sfence_bits_addr(ptw_io_dpath_sfence_bits_addr),
    .io_dpath_sfence_bits_asid(ptw_io_dpath_sfence_bits_asid),
    .io_dpath_status_debug(ptw_io_dpath_status_debug),
    .io_dpath_status_cease(ptw_io_dpath_status_cease),
    .io_dpath_status_wfi(ptw_io_dpath_status_wfi),
    .io_dpath_status_isa(ptw_io_dpath_status_isa),
    .io_dpath_status_dprv(ptw_io_dpath_status_dprv),
    .io_dpath_status_prv(ptw_io_dpath_status_prv),
    .io_dpath_status_sd(ptw_io_dpath_status_sd),
    .io_dpath_status_zero2(ptw_io_dpath_status_zero2),
    .io_dpath_status_sxl(ptw_io_dpath_status_sxl),
    .io_dpath_status_uxl(ptw_io_dpath_status_uxl),
    .io_dpath_status_sd_rv32(ptw_io_dpath_status_sd_rv32),
    .io_dpath_status_zero1(ptw_io_dpath_status_zero1),
    .io_dpath_status_tsr(ptw_io_dpath_status_tsr),
    .io_dpath_status_tw(ptw_io_dpath_status_tw),
    .io_dpath_status_tvm(ptw_io_dpath_status_tvm),
    .io_dpath_status_mxr(ptw_io_dpath_status_mxr),
    .io_dpath_status_sum(ptw_io_dpath_status_sum),
    .io_dpath_status_mprv(ptw_io_dpath_status_mprv),
    .io_dpath_status_xs(ptw_io_dpath_status_xs),
    .io_dpath_status_fs(ptw_io_dpath_status_fs),
    .io_dpath_status_mpp(ptw_io_dpath_status_mpp),
    .io_dpath_status_vs(ptw_io_dpath_status_vs),
    .io_dpath_status_spp(ptw_io_dpath_status_spp),
    .io_dpath_status_mpie(ptw_io_dpath_status_mpie),
    .io_dpath_status_hpie(ptw_io_dpath_status_hpie),
    .io_dpath_status_spie(ptw_io_dpath_status_spie),
    .io_dpath_status_upie(ptw_io_dpath_status_upie),
    .io_dpath_status_mie(ptw_io_dpath_status_mie),
    .io_dpath_status_hie(ptw_io_dpath_status_hie),
    .io_dpath_status_sie(ptw_io_dpath_status_sie),
    .io_dpath_status_uie(ptw_io_dpath_status_uie),
    .io_dpath_pmp_0_cfg_l(ptw_io_dpath_pmp_0_cfg_l),
    .io_dpath_pmp_0_cfg_res(ptw_io_dpath_pmp_0_cfg_res),
    .io_dpath_pmp_0_cfg_a(ptw_io_dpath_pmp_0_cfg_a),
    .io_dpath_pmp_0_cfg_x(ptw_io_dpath_pmp_0_cfg_x),
    .io_dpath_pmp_0_cfg_w(ptw_io_dpath_pmp_0_cfg_w),
    .io_dpath_pmp_0_cfg_r(ptw_io_dpath_pmp_0_cfg_r),
    .io_dpath_pmp_0_addr(ptw_io_dpath_pmp_0_addr),
    .io_dpath_pmp_0_mask(ptw_io_dpath_pmp_0_mask),
    .io_dpath_pmp_1_cfg_l(ptw_io_dpath_pmp_1_cfg_l),
    .io_dpath_pmp_1_cfg_res(ptw_io_dpath_pmp_1_cfg_res),
    .io_dpath_pmp_1_cfg_a(ptw_io_dpath_pmp_1_cfg_a),
    .io_dpath_pmp_1_cfg_x(ptw_io_dpath_pmp_1_cfg_x),
    .io_dpath_pmp_1_cfg_w(ptw_io_dpath_pmp_1_cfg_w),
    .io_dpath_pmp_1_cfg_r(ptw_io_dpath_pmp_1_cfg_r),
    .io_dpath_pmp_1_addr(ptw_io_dpath_pmp_1_addr),
    .io_dpath_pmp_1_mask(ptw_io_dpath_pmp_1_mask),
    .io_dpath_pmp_2_cfg_l(ptw_io_dpath_pmp_2_cfg_l),
    .io_dpath_pmp_2_cfg_res(ptw_io_dpath_pmp_2_cfg_res),
    .io_dpath_pmp_2_cfg_a(ptw_io_dpath_pmp_2_cfg_a),
    .io_dpath_pmp_2_cfg_x(ptw_io_dpath_pmp_2_cfg_x),
    .io_dpath_pmp_2_cfg_w(ptw_io_dpath_pmp_2_cfg_w),
    .io_dpath_pmp_2_cfg_r(ptw_io_dpath_pmp_2_cfg_r),
    .io_dpath_pmp_2_addr(ptw_io_dpath_pmp_2_addr),
    .io_dpath_pmp_2_mask(ptw_io_dpath_pmp_2_mask),
    .io_dpath_pmp_3_cfg_l(ptw_io_dpath_pmp_3_cfg_l),
    .io_dpath_pmp_3_cfg_res(ptw_io_dpath_pmp_3_cfg_res),
    .io_dpath_pmp_3_cfg_a(ptw_io_dpath_pmp_3_cfg_a),
    .io_dpath_pmp_3_cfg_x(ptw_io_dpath_pmp_3_cfg_x),
    .io_dpath_pmp_3_cfg_w(ptw_io_dpath_pmp_3_cfg_w),
    .io_dpath_pmp_3_cfg_r(ptw_io_dpath_pmp_3_cfg_r),
    .io_dpath_pmp_3_addr(ptw_io_dpath_pmp_3_addr),
    .io_dpath_pmp_3_mask(ptw_io_dpath_pmp_3_mask),
    .io_dpath_pmp_4_cfg_l(ptw_io_dpath_pmp_4_cfg_l),
    .io_dpath_pmp_4_cfg_res(ptw_io_dpath_pmp_4_cfg_res),
    .io_dpath_pmp_4_cfg_a(ptw_io_dpath_pmp_4_cfg_a),
    .io_dpath_pmp_4_cfg_x(ptw_io_dpath_pmp_4_cfg_x),
    .io_dpath_pmp_4_cfg_w(ptw_io_dpath_pmp_4_cfg_w),
    .io_dpath_pmp_4_cfg_r(ptw_io_dpath_pmp_4_cfg_r),
    .io_dpath_pmp_4_addr(ptw_io_dpath_pmp_4_addr),
    .io_dpath_pmp_4_mask(ptw_io_dpath_pmp_4_mask),
    .io_dpath_pmp_5_cfg_l(ptw_io_dpath_pmp_5_cfg_l),
    .io_dpath_pmp_5_cfg_res(ptw_io_dpath_pmp_5_cfg_res),
    .io_dpath_pmp_5_cfg_a(ptw_io_dpath_pmp_5_cfg_a),
    .io_dpath_pmp_5_cfg_x(ptw_io_dpath_pmp_5_cfg_x),
    .io_dpath_pmp_5_cfg_w(ptw_io_dpath_pmp_5_cfg_w),
    .io_dpath_pmp_5_cfg_r(ptw_io_dpath_pmp_5_cfg_r),
    .io_dpath_pmp_5_addr(ptw_io_dpath_pmp_5_addr),
    .io_dpath_pmp_5_mask(ptw_io_dpath_pmp_5_mask),
    .io_dpath_pmp_6_cfg_l(ptw_io_dpath_pmp_6_cfg_l),
    .io_dpath_pmp_6_cfg_res(ptw_io_dpath_pmp_6_cfg_res),
    .io_dpath_pmp_6_cfg_a(ptw_io_dpath_pmp_6_cfg_a),
    .io_dpath_pmp_6_cfg_x(ptw_io_dpath_pmp_6_cfg_x),
    .io_dpath_pmp_6_cfg_w(ptw_io_dpath_pmp_6_cfg_w),
    .io_dpath_pmp_6_cfg_r(ptw_io_dpath_pmp_6_cfg_r),
    .io_dpath_pmp_6_addr(ptw_io_dpath_pmp_6_addr),
    .io_dpath_pmp_6_mask(ptw_io_dpath_pmp_6_mask),
    .io_dpath_pmp_7_cfg_l(ptw_io_dpath_pmp_7_cfg_l),
    .io_dpath_pmp_7_cfg_res(ptw_io_dpath_pmp_7_cfg_res),
    .io_dpath_pmp_7_cfg_a(ptw_io_dpath_pmp_7_cfg_a),
    .io_dpath_pmp_7_cfg_x(ptw_io_dpath_pmp_7_cfg_x),
    .io_dpath_pmp_7_cfg_w(ptw_io_dpath_pmp_7_cfg_w),
    .io_dpath_pmp_7_cfg_r(ptw_io_dpath_pmp_7_cfg_r),
    .io_dpath_pmp_7_addr(ptw_io_dpath_pmp_7_addr),
    .io_dpath_pmp_7_mask(ptw_io_dpath_pmp_7_mask),
    .io_dpath_perf_l2miss(ptw_io_dpath_perf_l2miss),
    .io_dpath_perf_l2hit(ptw_io_dpath_perf_l2hit),
    .io_dpath_perf_pte_miss(ptw_io_dpath_perf_pte_miss),
    .io_dpath_perf_pte_hit(ptw_io_dpath_perf_pte_hit),
    .io_dpath_customCSRs_csrs_0_wen(ptw_io_dpath_customCSRs_csrs_0_wen),
    .io_dpath_customCSRs_csrs_0_wdata(ptw_io_dpath_customCSRs_csrs_0_wdata),
    .io_dpath_customCSRs_csrs_0_value(ptw_io_dpath_customCSRs_csrs_0_value),
    .io_dpath_clock_enabled(ptw_io_dpath_clock_enabled)
  );
  HellaCacheArbiter hellaCacheArb ( // @[tile.scala 236:29]
    .clock(hellaCacheArb_clock),
    .reset(hellaCacheArb_reset),
    .io_requestor_0_req_ready(hellaCacheArb_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(hellaCacheArb_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_addr(hellaCacheArb_io_requestor_0_req_bits_addr),
    .io_requestor_0_req_bits_tag(hellaCacheArb_io_requestor_0_req_bits_tag),
    .io_requestor_0_req_bits_cmd(hellaCacheArb_io_requestor_0_req_bits_cmd),
    .io_requestor_0_req_bits_size(hellaCacheArb_io_requestor_0_req_bits_size),
    .io_requestor_0_req_bits_signed(hellaCacheArb_io_requestor_0_req_bits_signed),
    .io_requestor_0_req_bits_dprv(hellaCacheArb_io_requestor_0_req_bits_dprv),
    .io_requestor_0_req_bits_phys(hellaCacheArb_io_requestor_0_req_bits_phys),
    .io_requestor_0_req_bits_no_alloc(hellaCacheArb_io_requestor_0_req_bits_no_alloc),
    .io_requestor_0_req_bits_no_xcpt(hellaCacheArb_io_requestor_0_req_bits_no_xcpt),
    .io_requestor_0_req_bits_data(hellaCacheArb_io_requestor_0_req_bits_data),
    .io_requestor_0_req_bits_mask(hellaCacheArb_io_requestor_0_req_bits_mask),
    .io_requestor_0_s1_kill(hellaCacheArb_io_requestor_0_s1_kill),
    .io_requestor_0_s1_data_data(hellaCacheArb_io_requestor_0_s1_data_data),
    .io_requestor_0_s1_data_mask(hellaCacheArb_io_requestor_0_s1_data_mask),
    .io_requestor_0_s2_nack(hellaCacheArb_io_requestor_0_s2_nack),
    .io_requestor_0_s2_nack_cause_raw(hellaCacheArb_io_requestor_0_s2_nack_cause_raw),
    .io_requestor_0_s2_kill(hellaCacheArb_io_requestor_0_s2_kill),
    .io_requestor_0_s2_uncached(hellaCacheArb_io_requestor_0_s2_uncached),
    .io_requestor_0_s2_paddr(hellaCacheArb_io_requestor_0_s2_paddr),
    .io_requestor_0_resp_valid(hellaCacheArb_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_addr(hellaCacheArb_io_requestor_0_resp_bits_addr),
    .io_requestor_0_resp_bits_tag(hellaCacheArb_io_requestor_0_resp_bits_tag),
    .io_requestor_0_resp_bits_cmd(hellaCacheArb_io_requestor_0_resp_bits_cmd),
    .io_requestor_0_resp_bits_size(hellaCacheArb_io_requestor_0_resp_bits_size),
    .io_requestor_0_resp_bits_signed(hellaCacheArb_io_requestor_0_resp_bits_signed),
    .io_requestor_0_resp_bits_dprv(hellaCacheArb_io_requestor_0_resp_bits_dprv),
    .io_requestor_0_resp_bits_data(hellaCacheArb_io_requestor_0_resp_bits_data),
    .io_requestor_0_resp_bits_mask(hellaCacheArb_io_requestor_0_resp_bits_mask),
    .io_requestor_0_resp_bits_replay(hellaCacheArb_io_requestor_0_resp_bits_replay),
    .io_requestor_0_resp_bits_has_data(hellaCacheArb_io_requestor_0_resp_bits_has_data),
    .io_requestor_0_resp_bits_data_word_bypass(hellaCacheArb_io_requestor_0_resp_bits_data_word_bypass),
    .io_requestor_0_resp_bits_data_raw(hellaCacheArb_io_requestor_0_resp_bits_data_raw),
    .io_requestor_0_resp_bits_store_data(hellaCacheArb_io_requestor_0_resp_bits_store_data),
    .io_requestor_0_replay_next(hellaCacheArb_io_requestor_0_replay_next),
    .io_requestor_0_s2_xcpt_ma_ld(hellaCacheArb_io_requestor_0_s2_xcpt_ma_ld),
    .io_requestor_0_s2_xcpt_ma_st(hellaCacheArb_io_requestor_0_s2_xcpt_ma_st),
    .io_requestor_0_s2_xcpt_pf_ld(hellaCacheArb_io_requestor_0_s2_xcpt_pf_ld),
    .io_requestor_0_s2_xcpt_pf_st(hellaCacheArb_io_requestor_0_s2_xcpt_pf_st),
    .io_requestor_0_s2_xcpt_ae_ld(hellaCacheArb_io_requestor_0_s2_xcpt_ae_ld),
    .io_requestor_0_s2_xcpt_ae_st(hellaCacheArb_io_requestor_0_s2_xcpt_ae_st),
    .io_requestor_0_ordered(hellaCacheArb_io_requestor_0_ordered),
    .io_requestor_0_perf_acquire(hellaCacheArb_io_requestor_0_perf_acquire),
    .io_requestor_0_perf_release(hellaCacheArb_io_requestor_0_perf_release),
    .io_requestor_0_perf_grant(hellaCacheArb_io_requestor_0_perf_grant),
    .io_requestor_0_perf_tlbMiss(hellaCacheArb_io_requestor_0_perf_tlbMiss),
    .io_requestor_0_perf_blocked(hellaCacheArb_io_requestor_0_perf_blocked),
    .io_requestor_0_perf_canAcceptStoreThenLoad(hellaCacheArb_io_requestor_0_perf_canAcceptStoreThenLoad),
    .io_requestor_0_perf_canAcceptStoreThenRMW(hellaCacheArb_io_requestor_0_perf_canAcceptStoreThenRMW),
    .io_requestor_0_perf_canAcceptLoadThenLoad(hellaCacheArb_io_requestor_0_perf_canAcceptLoadThenLoad),
    .io_requestor_0_perf_storeBufferEmptyAfterLoad(hellaCacheArb_io_requestor_0_perf_storeBufferEmptyAfterLoad),
    .io_requestor_0_perf_storeBufferEmptyAfterStore(hellaCacheArb_io_requestor_0_perf_storeBufferEmptyAfterStore),
    .io_requestor_0_keep_clock_enabled(hellaCacheArb_io_requestor_0_keep_clock_enabled),
    .io_requestor_0_clock_enabled(hellaCacheArb_io_requestor_0_clock_enabled),
    .io_mem_req_ready(hellaCacheArb_io_mem_req_ready),
    .io_mem_req_valid(hellaCacheArb_io_mem_req_valid),
    .io_mem_req_bits_addr(hellaCacheArb_io_mem_req_bits_addr),
    .io_mem_req_bits_tag(hellaCacheArb_io_mem_req_bits_tag),
    .io_mem_req_bits_cmd(hellaCacheArb_io_mem_req_bits_cmd),
    .io_mem_req_bits_size(hellaCacheArb_io_mem_req_bits_size),
    .io_mem_req_bits_signed(hellaCacheArb_io_mem_req_bits_signed),
    .io_mem_req_bits_dprv(hellaCacheArb_io_mem_req_bits_dprv),
    .io_mem_req_bits_phys(hellaCacheArb_io_mem_req_bits_phys),
    .io_mem_req_bits_no_alloc(hellaCacheArb_io_mem_req_bits_no_alloc),
    .io_mem_req_bits_no_xcpt(hellaCacheArb_io_mem_req_bits_no_xcpt),
    .io_mem_req_bits_data(hellaCacheArb_io_mem_req_bits_data),
    .io_mem_req_bits_mask(hellaCacheArb_io_mem_req_bits_mask),
    .io_mem_s1_kill(hellaCacheArb_io_mem_s1_kill),
    .io_mem_s1_data_data(hellaCacheArb_io_mem_s1_data_data),
    .io_mem_s1_data_mask(hellaCacheArb_io_mem_s1_data_mask),
    .io_mem_s2_nack(hellaCacheArb_io_mem_s2_nack),
    .io_mem_s2_nack_cause_raw(hellaCacheArb_io_mem_s2_nack_cause_raw),
    .io_mem_s2_kill(hellaCacheArb_io_mem_s2_kill),
    .io_mem_s2_uncached(hellaCacheArb_io_mem_s2_uncached),
    .io_mem_s2_paddr(hellaCacheArb_io_mem_s2_paddr),
    .io_mem_resp_valid(hellaCacheArb_io_mem_resp_valid),
    .io_mem_resp_bits_addr(hellaCacheArb_io_mem_resp_bits_addr),
    .io_mem_resp_bits_tag(hellaCacheArb_io_mem_resp_bits_tag),
    .io_mem_resp_bits_cmd(hellaCacheArb_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_size(hellaCacheArb_io_mem_resp_bits_size),
    .io_mem_resp_bits_signed(hellaCacheArb_io_mem_resp_bits_signed),
    .io_mem_resp_bits_dprv(hellaCacheArb_io_mem_resp_bits_dprv),
    .io_mem_resp_bits_data(hellaCacheArb_io_mem_resp_bits_data),
    .io_mem_resp_bits_mask(hellaCacheArb_io_mem_resp_bits_mask),
    .io_mem_resp_bits_replay(hellaCacheArb_io_mem_resp_bits_replay),
    .io_mem_resp_bits_has_data(hellaCacheArb_io_mem_resp_bits_has_data),
    .io_mem_resp_bits_data_word_bypass(hellaCacheArb_io_mem_resp_bits_data_word_bypass),
    .io_mem_resp_bits_data_raw(hellaCacheArb_io_mem_resp_bits_data_raw),
    .io_mem_resp_bits_store_data(hellaCacheArb_io_mem_resp_bits_store_data),
    .io_mem_replay_next(hellaCacheArb_io_mem_replay_next),
    .io_mem_s2_xcpt_ma_ld(hellaCacheArb_io_mem_s2_xcpt_ma_ld),
    .io_mem_s2_xcpt_ma_st(hellaCacheArb_io_mem_s2_xcpt_ma_st),
    .io_mem_s2_xcpt_pf_ld(hellaCacheArb_io_mem_s2_xcpt_pf_ld),
    .io_mem_s2_xcpt_pf_st(hellaCacheArb_io_mem_s2_xcpt_pf_st),
    .io_mem_s2_xcpt_ae_ld(hellaCacheArb_io_mem_s2_xcpt_ae_ld),
    .io_mem_s2_xcpt_ae_st(hellaCacheArb_io_mem_s2_xcpt_ae_st),
    .io_mem_ordered(hellaCacheArb_io_mem_ordered),
    .io_mem_perf_acquire(hellaCacheArb_io_mem_perf_acquire),
    .io_mem_perf_release(hellaCacheArb_io_mem_perf_release),
    .io_mem_perf_grant(hellaCacheArb_io_mem_perf_grant),
    .io_mem_perf_tlbMiss(hellaCacheArb_io_mem_perf_tlbMiss),
    .io_mem_perf_blocked(hellaCacheArb_io_mem_perf_blocked),
    .io_mem_perf_canAcceptStoreThenLoad(hellaCacheArb_io_mem_perf_canAcceptStoreThenLoad),
    .io_mem_perf_canAcceptStoreThenRMW(hellaCacheArb_io_mem_perf_canAcceptStoreThenRMW),
    .io_mem_perf_canAcceptLoadThenLoad(hellaCacheArb_io_mem_perf_canAcceptLoadThenLoad),
    .io_mem_perf_storeBufferEmptyAfterLoad(hellaCacheArb_io_mem_perf_storeBufferEmptyAfterLoad),
    .io_mem_perf_storeBufferEmptyAfterStore(hellaCacheArb_io_mem_perf_storeBufferEmptyAfterStore),
    .io_mem_keep_clock_enabled(hellaCacheArb_io_mem_keep_clock_enabled),
    .io_mem_clock_enabled(hellaCacheArb_io_mem_clock_enabled)
  );
  assign auto_trace_out_0_valid = trace_auto_out_0_valid; // @[LazyModule.scala 311:12]
  assign auto_trace_out_0_iaddr = trace_auto_out_0_iaddr; // @[LazyModule.scala 311:12]
  assign auto_trace_out_0_insn = trace_auto_out_0_insn; // @[LazyModule.scala 311:12]
  assign auto_trace_out_0_priv = trace_auto_out_0_priv; // @[LazyModule.scala 311:12]
  assign auto_trace_out_0_exception = trace_auto_out_0_exception; // @[LazyModule.scala 311:12]
  assign auto_trace_out_0_interrupt = trace_auto_out_0_interrupt; // @[LazyModule.scala 311:12]
  assign auto_trace_out_0_cause = trace_auto_out_0_cause; // @[LazyModule.scala 311:12]
  assign auto_trace_out_0_tval = trace_auto_out_0_tval; // @[LazyModule.scala 311:12]
  assign auto_trace_out_0_wdata = trace_auto_out_0_wdata; // @[LazyModule.scala 311:12]
  assign auto_trace_out_1_valid = trace_auto_out_1_valid; // @[LazyModule.scala 311:12]
  assign auto_trace_out_1_iaddr = trace_auto_out_1_iaddr; // @[LazyModule.scala 311:12]
  assign auto_trace_out_1_insn = trace_auto_out_1_insn; // @[LazyModule.scala 311:12]
  assign auto_trace_out_1_priv = trace_auto_out_1_priv; // @[LazyModule.scala 311:12]
  assign auto_trace_out_1_exception = trace_auto_out_1_exception; // @[LazyModule.scala 311:12]
  assign auto_trace_out_1_interrupt = trace_auto_out_1_interrupt; // @[LazyModule.scala 311:12]
  assign auto_trace_out_1_cause = trace_auto_out_1_cause; // @[LazyModule.scala 311:12]
  assign auto_trace_out_1_tval = trace_auto_out_1_tval; // @[LazyModule.scala 311:12]
  assign auto_trace_out_1_wdata = trace_auto_out_1_wdata; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_0_valid = broadcast_3_auto_out_0_valid; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_0_iaddr = broadcast_3_auto_out_0_iaddr; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_0_insn = broadcast_3_auto_out_0_insn; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_0_priv = broadcast_3_auto_out_0_priv; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_0_exception = broadcast_3_auto_out_0_exception; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_0_interrupt = broadcast_3_auto_out_0_interrupt; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_0_cause = broadcast_3_auto_out_0_cause; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_0_tval = broadcast_3_auto_out_0_tval; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_1_valid = broadcast_3_auto_out_1_valid; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_1_iaddr = broadcast_3_auto_out_1_iaddr; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_1_insn = broadcast_3_auto_out_1_insn; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_1_priv = broadcast_3_auto_out_1_priv; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_1_exception = broadcast_3_auto_out_1_exception; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_1_interrupt = broadcast_3_auto_out_1_interrupt; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_1_cause = broadcast_3_auto_out_1_cause; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_1_tval = broadcast_3_auto_out_1_tval; // @[LazyModule.scala 311:12]
  assign auto_wfi_out_0 = 1'h0; // @[Nodes.scala 1207:84 Interrupts.scala 129:12]
  assign auto_cease_out_0 = 1'h0; // @[LazyModule.scala 311:12]
  assign auto_halt_out_0 = 1'h0; // @[LazyModule.scala 311:12]
  assign auto_trace_core_source_out_group_0_iretire = 1'h0; // @[LazyModule.scala 311:12]
  assign auto_trace_core_source_out_group_0_iaddr = 32'h0; // @[LazyModule.scala 311:12]
  assign auto_trace_core_source_out_group_0_itype = 4'h0; // @[LazyModule.scala 311:12]
  assign auto_trace_core_source_out_group_0_ilastsize = 1'h0; // @[LazyModule.scala 311:12]
  assign auto_trace_core_source_out_priv = 4'h0; // @[LazyModule.scala 311:12]
  assign auto_trace_core_source_out_tval = 32'h0; // @[LazyModule.scala 311:12]
  assign auto_trace_core_source_out_cause = 32'h0; // @[LazyModule.scala 311:12]
  assign auto_tl_other_masters_out_a_valid = tlMasterXbar_auto_out_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_opcode = tlMasterXbar_auto_out_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_param = tlMasterXbar_auto_out_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_size = tlMasterXbar_auto_out_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_source = tlMasterXbar_auto_out_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_address = tlMasterXbar_auto_out_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_mask = tlMasterXbar_auto_out_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_data = tlMasterXbar_auto_out_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_a_bits_corrupt = tlMasterXbar_auto_out_a_bits_corrupt; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_b_ready = tlMasterXbar_auto_out_b_ready; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_c_valid = tlMasterXbar_auto_out_c_valid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_c_bits_opcode = tlMasterXbar_auto_out_c_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_c_bits_param = tlMasterXbar_auto_out_c_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_c_bits_size = tlMasterXbar_auto_out_c_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_c_bits_source = tlMasterXbar_auto_out_c_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_c_bits_address = tlMasterXbar_auto_out_c_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_c_bits_data = tlMasterXbar_auto_out_c_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_c_bits_corrupt = tlMasterXbar_auto_out_c_bits_corrupt; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_d_ready = tlMasterXbar_auto_out_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_e_valid = tlMasterXbar_auto_out_e_valid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign auto_tl_other_masters_out_e_bits_sink = tlMasterXbar_auto_out_e_bits_sink; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_clock = clock;
  assign tlMasterXbar_reset = reset;
  assign tlMasterXbar_auto_in_1_a_valid = frontend_auto_icache_master_out_a_valid; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_1_a_bits_opcode = frontend_auto_icache_master_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_1_a_bits_param = frontend_auto_icache_master_out_a_bits_param; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_1_a_bits_size = frontend_auto_icache_master_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_1_a_bits_source = frontend_auto_icache_master_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_1_a_bits_address = frontend_auto_icache_master_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_1_a_bits_mask = frontend_auto_icache_master_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_1_a_bits_data = frontend_auto_icache_master_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_1_a_bits_corrupt = frontend_auto_icache_master_out_a_bits_corrupt; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_1_d_ready = frontend_auto_icache_master_out_d_ready; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_a_valid = dcache_auto_out_a_valid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_a_bits_opcode = dcache_auto_out_a_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_a_bits_param = dcache_auto_out_a_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_a_bits_size = dcache_auto_out_a_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_a_bits_source = dcache_auto_out_a_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_a_bits_address = dcache_auto_out_a_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_a_bits_mask = dcache_auto_out_a_bits_mask; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_a_bits_data = dcache_auto_out_a_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_a_bits_corrupt = dcache_auto_out_a_bits_corrupt; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_b_ready = dcache_auto_out_b_ready; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_c_valid = dcache_auto_out_c_valid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_c_bits_opcode = dcache_auto_out_c_bits_opcode; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_c_bits_param = dcache_auto_out_c_bits_param; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_c_bits_size = dcache_auto_out_c_bits_size; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_c_bits_source = dcache_auto_out_c_bits_source; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_c_bits_address = dcache_auto_out_c_bits_address; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_c_bits_data = dcache_auto_out_c_bits_data; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_c_bits_corrupt = dcache_auto_out_c_bits_corrupt; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_d_ready = dcache_auto_out_d_ready; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_e_valid = dcache_auto_out_e_valid; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_e_bits_sink = dcache_auto_out_e_bits_sink; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_a_ready = auto_tl_other_masters_out_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_b_valid = auto_tl_other_masters_out_b_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_b_bits_opcode = auto_tl_other_masters_out_b_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_b_bits_param = auto_tl_other_masters_out_b_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_b_bits_size = auto_tl_other_masters_out_b_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_b_bits_source = auto_tl_other_masters_out_b_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_b_bits_address = auto_tl_other_masters_out_b_bits_address; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_b_bits_mask = auto_tl_other_masters_out_b_bits_mask; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_b_bits_data = auto_tl_other_masters_out_b_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_b_bits_corrupt = auto_tl_other_masters_out_b_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_c_ready = auto_tl_other_masters_out_c_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_d_valid = auto_tl_other_masters_out_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_d_bits_opcode = auto_tl_other_masters_out_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_d_bits_param = auto_tl_other_masters_out_d_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_d_bits_size = auto_tl_other_masters_out_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_d_bits_source = auto_tl_other_masters_out_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_d_bits_sink = auto_tl_other_masters_out_d_bits_sink; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_d_bits_denied = auto_tl_other_masters_out_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_d_bits_data = auto_tl_other_masters_out_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_d_bits_corrupt = auto_tl_other_masters_out_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlMasterXbar_auto_out_e_ready = auto_tl_other_masters_out_e_ready; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign tlSlaveXbar_clock = clock;
  assign tlSlaveXbar_reset = reset;
  assign intXbar_clock = clock;
  assign intXbar_reset = reset;
  assign intXbar_auto_int_in_3_0 = auto_int_local_in_3_0; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign intXbar_auto_int_in_2_0 = auto_int_local_in_2_0; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign intXbar_auto_int_in_1_0 = auto_int_local_in_1_0; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign intXbar_auto_int_in_1_1 = auto_int_local_in_1_1; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign intXbar_auto_int_in_0_0 = auto_int_local_in_0_0; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign broadcast_clock = clock;
  assign broadcast_reset = reset;
  assign broadcast_auto_in = auto_hartid_in; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign broadcast_1_clock = clock;
  assign broadcast_1_reset = reset;
  assign broadcast_1_auto_in = auto_reset_vector_in; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign broadcast_2_clock = clock;
  assign broadcast_2_reset = reset;
  assign broadcast_2_auto_in_rnmi = auto_nmi_in_rnmi; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign broadcast_2_auto_in_rnmi_interrupt_vector = auto_nmi_in_rnmi_interrupt_vector; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign broadcast_2_auto_in_rnmi_exception_vector = auto_nmi_in_rnmi_exception_vector; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign broadcast_2_auto_in_unmi = auto_nmi_in_unmi; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign broadcast_2_auto_in_unmi_interrupt_vector = auto_nmi_in_unmi_interrupt_vector; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign broadcast_2_auto_in_unmi_exception_vector = auto_nmi_in_unmi_exception_vector; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  assign nexus_clock = clock;
  assign nexus_reset = reset;
  assign broadcast_3_clock = clock;
  assign broadcast_3_reset = reset;
  assign broadcast_3_auto_in_0_valid = 1'h0; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_0_iaddr = 40'h0; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_0_insn = 32'h0; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_0_priv = 3'h0; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_0_exception = 1'h0; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_0_interrupt = 1'h0; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_0_cause = 64'h0; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_0_tval = 40'h0; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_1_valid = 1'h0; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_1_iaddr = 40'h0; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_1_insn = 32'h0; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_1_priv = 3'h0; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_1_exception = 1'h0; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_1_interrupt = 1'h0; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_1_cause = 64'h0; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_1_tval = 40'h0; // @[LazyModule.scala 298:16]
  assign nexus_1_clock = clock;
  assign nexus_1_reset = reset;
  assign broadcast_4_clock = clock;
  assign broadcast_4_reset = reset;
  assign trace_clock = clock;
  assign trace_reset = reset;
  assign trace_auto_in_0_valid = core_io_trace_0_valid; // @[Nodes.scala 1207:84 tile.scala 171:35]
  assign trace_auto_in_0_iaddr = core_io_trace_0_iaddr; // @[Nodes.scala 1207:84 tile.scala 171:35]
  assign trace_auto_in_0_insn = core_io_trace_0_insn; // @[Nodes.scala 1207:84 tile.scala 171:35]
  assign trace_auto_in_0_priv = core_io_trace_0_priv; // @[Nodes.scala 1207:84 tile.scala 171:35]
  assign trace_auto_in_0_exception = core_io_trace_0_exception; // @[Nodes.scala 1207:84 tile.scala 171:35]
  assign trace_auto_in_0_interrupt = core_io_trace_0_interrupt; // @[Nodes.scala 1207:84 tile.scala 171:35]
  assign trace_auto_in_0_cause = core_io_trace_0_cause; // @[Nodes.scala 1207:84 tile.scala 171:35]
  assign trace_auto_in_0_tval = core_io_trace_0_tval; // @[Nodes.scala 1207:84 tile.scala 171:35]
  assign trace_auto_in_0_wdata = core_io_trace_0_wdata; // @[Nodes.scala 1207:84 tile.scala 171:35]
  assign trace_auto_in_1_valid = core_io_trace_1_valid; // @[Nodes.scala 1207:84 tile.scala 171:35]
  assign trace_auto_in_1_iaddr = core_io_trace_1_iaddr; // @[Nodes.scala 1207:84 tile.scala 171:35]
  assign trace_auto_in_1_insn = core_io_trace_1_insn; // @[Nodes.scala 1207:84 tile.scala 171:35]
  assign trace_auto_in_1_priv = core_io_trace_1_priv; // @[Nodes.scala 1207:84 tile.scala 171:35]
  assign trace_auto_in_1_exception = core_io_trace_1_exception; // @[Nodes.scala 1207:84 tile.scala 171:35]
  assign trace_auto_in_1_interrupt = core_io_trace_1_interrupt; // @[Nodes.scala 1207:84 tile.scala 171:35]
  assign trace_auto_in_1_cause = core_io_trace_1_cause; // @[Nodes.scala 1207:84 tile.scala 171:35]
  assign trace_auto_in_1_tval = core_io_trace_1_tval; // @[Nodes.scala 1207:84 tile.scala 171:35]
  assign trace_auto_in_1_wdata = core_io_trace_1_wdata; // @[Nodes.scala 1207:84 tile.scala 171:35]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_auto_out_a_ready = tlMasterXbar_auto_in_0_a_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign dcache_auto_out_b_valid = tlMasterXbar_auto_in_0_b_valid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign dcache_auto_out_b_bits_opcode = tlMasterXbar_auto_in_0_b_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign dcache_auto_out_b_bits_param = tlMasterXbar_auto_in_0_b_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign dcache_auto_out_b_bits_size = tlMasterXbar_auto_in_0_b_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign dcache_auto_out_b_bits_source = tlMasterXbar_auto_in_0_b_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign dcache_auto_out_b_bits_address = tlMasterXbar_auto_in_0_b_bits_address; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign dcache_auto_out_b_bits_mask = tlMasterXbar_auto_in_0_b_bits_mask; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign dcache_auto_out_b_bits_data = tlMasterXbar_auto_in_0_b_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign dcache_auto_out_b_bits_corrupt = tlMasterXbar_auto_in_0_b_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign dcache_auto_out_c_ready = tlMasterXbar_auto_in_0_c_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign dcache_auto_out_d_valid = tlMasterXbar_auto_in_0_d_valid; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign dcache_auto_out_d_bits_opcode = tlMasterXbar_auto_in_0_d_bits_opcode; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign dcache_auto_out_d_bits_param = tlMasterXbar_auto_in_0_d_bits_param; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign dcache_auto_out_d_bits_size = tlMasterXbar_auto_in_0_d_bits_size; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign dcache_auto_out_d_bits_source = tlMasterXbar_auto_in_0_d_bits_source; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign dcache_auto_out_d_bits_sink = tlMasterXbar_auto_in_0_d_bits_sink; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign dcache_auto_out_d_bits_denied = tlMasterXbar_auto_in_0_d_bits_denied; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign dcache_auto_out_d_bits_data = tlMasterXbar_auto_in_0_d_bits_data; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign dcache_auto_out_d_bits_corrupt = tlMasterXbar_auto_in_0_d_bits_corrupt; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign dcache_auto_out_e_ready = tlMasterXbar_auto_in_0_e_ready; // @[Nodes.scala 1207:84 LazyModule.scala 298:16]
  assign dcache_io_lsu_req_valid = lsu_io_dmem_req_valid; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_valid = lsu_io_dmem_req_bits_0_valid; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_switch = lsu_io_dmem_req_bits_0_bits_uop_switch; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_switch_off = lsu_io_dmem_req_bits_0_bits_uop_switch_off; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_is_unicore = lsu_io_dmem_req_bits_0_bits_uop_is_unicore; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_shift = lsu_io_dmem_req_bits_0_bits_uop_shift; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_lrs3_rtype = lsu_io_dmem_req_bits_0_bits_uop_lrs3_rtype; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_rflag = lsu_io_dmem_req_bits_0_bits_uop_rflag; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_wflag = lsu_io_dmem_req_bits_0_bits_uop_wflag; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_prflag = lsu_io_dmem_req_bits_0_bits_uop_prflag; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_pwflag = lsu_io_dmem_req_bits_0_bits_uop_pwflag; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_pflag_busy = lsu_io_dmem_req_bits_0_bits_uop_pflag_busy; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_stale_pflag = lsu_io_dmem_req_bits_0_bits_uop_stale_pflag; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_op1_sel = lsu_io_dmem_req_bits_0_bits_uop_op1_sel; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_op2_sel = lsu_io_dmem_req_bits_0_bits_uop_op2_sel; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_split_num = lsu_io_dmem_req_bits_0_bits_uop_split_num; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_self_index = lsu_io_dmem_req_bits_0_bits_uop_self_index; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_rob_inst_idx = lsu_io_dmem_req_bits_0_bits_uop_rob_inst_idx; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_address_num = lsu_io_dmem_req_bits_0_bits_uop_address_num; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_uopc = lsu_io_dmem_req_bits_0_bits_uop_uopc; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_inst = lsu_io_dmem_req_bits_0_bits_uop_inst; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_debug_inst = lsu_io_dmem_req_bits_0_bits_uop_debug_inst; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_is_rvc = lsu_io_dmem_req_bits_0_bits_uop_is_rvc; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_debug_pc = lsu_io_dmem_req_bits_0_bits_uop_debug_pc; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_iq_type = lsu_io_dmem_req_bits_0_bits_uop_iq_type; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_fu_code = lsu_io_dmem_req_bits_0_bits_uop_fu_code; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_ctrl_br_type = lsu_io_dmem_req_bits_0_bits_uop_ctrl_br_type; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_ctrl_op1_sel = lsu_io_dmem_req_bits_0_bits_uop_ctrl_op1_sel; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_ctrl_op2_sel = lsu_io_dmem_req_bits_0_bits_uop_ctrl_op2_sel; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_ctrl_imm_sel = lsu_io_dmem_req_bits_0_bits_uop_ctrl_imm_sel; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_ctrl_op_fcn = lsu_io_dmem_req_bits_0_bits_uop_ctrl_op_fcn; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_ctrl_fcn_dw = lsu_io_dmem_req_bits_0_bits_uop_ctrl_fcn_dw; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_ctrl_csr_cmd = lsu_io_dmem_req_bits_0_bits_uop_ctrl_csr_cmd; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_ctrl_is_load = lsu_io_dmem_req_bits_0_bits_uop_ctrl_is_load; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_ctrl_is_sta = lsu_io_dmem_req_bits_0_bits_uop_ctrl_is_sta; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_ctrl_is_std = lsu_io_dmem_req_bits_0_bits_uop_ctrl_is_std; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_ctrl_op3_sel = lsu_io_dmem_req_bits_0_bits_uop_ctrl_op3_sel; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_iw_state = lsu_io_dmem_req_bits_0_bits_uop_iw_state; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_iw_p1_poisoned = lsu_io_dmem_req_bits_0_bits_uop_iw_p1_poisoned; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_iw_p2_poisoned = lsu_io_dmem_req_bits_0_bits_uop_iw_p2_poisoned; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_is_br = lsu_io_dmem_req_bits_0_bits_uop_is_br; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_is_jalr = lsu_io_dmem_req_bits_0_bits_uop_is_jalr; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_is_jal = lsu_io_dmem_req_bits_0_bits_uop_is_jal; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_is_sfb = lsu_io_dmem_req_bits_0_bits_uop_is_sfb; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_br_mask = lsu_io_dmem_req_bits_0_bits_uop_br_mask; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_br_tag = lsu_io_dmem_req_bits_0_bits_uop_br_tag; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_ftq_idx = lsu_io_dmem_req_bits_0_bits_uop_ftq_idx; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_edge_inst = lsu_io_dmem_req_bits_0_bits_uop_edge_inst; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_pc_lob = lsu_io_dmem_req_bits_0_bits_uop_pc_lob; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_taken = lsu_io_dmem_req_bits_0_bits_uop_taken; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_imm_packed = lsu_io_dmem_req_bits_0_bits_uop_imm_packed; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_csr_addr = lsu_io_dmem_req_bits_0_bits_uop_csr_addr; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_rob_idx = lsu_io_dmem_req_bits_0_bits_uop_rob_idx; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_ldq_idx = lsu_io_dmem_req_bits_0_bits_uop_ldq_idx; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_stq_idx = lsu_io_dmem_req_bits_0_bits_uop_stq_idx; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_rxq_idx = lsu_io_dmem_req_bits_0_bits_uop_rxq_idx; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_pdst = lsu_io_dmem_req_bits_0_bits_uop_pdst; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_prs1 = lsu_io_dmem_req_bits_0_bits_uop_prs1; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_prs2 = lsu_io_dmem_req_bits_0_bits_uop_prs2; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_prs3 = lsu_io_dmem_req_bits_0_bits_uop_prs3; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_ppred = lsu_io_dmem_req_bits_0_bits_uop_ppred; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_prs1_busy = lsu_io_dmem_req_bits_0_bits_uop_prs1_busy; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_prs2_busy = lsu_io_dmem_req_bits_0_bits_uop_prs2_busy; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_prs3_busy = lsu_io_dmem_req_bits_0_bits_uop_prs3_busy; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_ppred_busy = lsu_io_dmem_req_bits_0_bits_uop_ppred_busy; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_stale_pdst = lsu_io_dmem_req_bits_0_bits_uop_stale_pdst; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_exception = lsu_io_dmem_req_bits_0_bits_uop_exception; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_exc_cause = lsu_io_dmem_req_bits_0_bits_uop_exc_cause; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_bypassable = lsu_io_dmem_req_bits_0_bits_uop_bypassable; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_mem_cmd = lsu_io_dmem_req_bits_0_bits_uop_mem_cmd; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_mem_size = lsu_io_dmem_req_bits_0_bits_uop_mem_size; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_mem_signed = lsu_io_dmem_req_bits_0_bits_uop_mem_signed; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_is_fence = lsu_io_dmem_req_bits_0_bits_uop_is_fence; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_is_fencei = lsu_io_dmem_req_bits_0_bits_uop_is_fencei; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_is_amo = lsu_io_dmem_req_bits_0_bits_uop_is_amo; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_uses_ldq = lsu_io_dmem_req_bits_0_bits_uop_uses_ldq; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_uses_stq = lsu_io_dmem_req_bits_0_bits_uop_uses_stq; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_is_sys_pc2epc = lsu_io_dmem_req_bits_0_bits_uop_is_sys_pc2epc; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_is_unique = lsu_io_dmem_req_bits_0_bits_uop_is_unique; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_flush_on_commit = lsu_io_dmem_req_bits_0_bits_uop_flush_on_commit; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_ldst_is_rs1 = lsu_io_dmem_req_bits_0_bits_uop_ldst_is_rs1; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_ldst = lsu_io_dmem_req_bits_0_bits_uop_ldst; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_lrs1 = lsu_io_dmem_req_bits_0_bits_uop_lrs1; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_lrs2 = lsu_io_dmem_req_bits_0_bits_uop_lrs2; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_lrs3 = lsu_io_dmem_req_bits_0_bits_uop_lrs3; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_ldst_val = lsu_io_dmem_req_bits_0_bits_uop_ldst_val; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_dst_rtype = lsu_io_dmem_req_bits_0_bits_uop_dst_rtype; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_lrs1_rtype = lsu_io_dmem_req_bits_0_bits_uop_lrs1_rtype; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_lrs2_rtype = lsu_io_dmem_req_bits_0_bits_uop_lrs2_rtype; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_frs3_en = lsu_io_dmem_req_bits_0_bits_uop_frs3_en; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_fp_val = lsu_io_dmem_req_bits_0_bits_uop_fp_val; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_fp_single = lsu_io_dmem_req_bits_0_bits_uop_fp_single; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_xcpt_pf_if = lsu_io_dmem_req_bits_0_bits_uop_xcpt_pf_if; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_xcpt_ae_if = lsu_io_dmem_req_bits_0_bits_uop_xcpt_ae_if; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_xcpt_ma_if = lsu_io_dmem_req_bits_0_bits_uop_xcpt_ma_if; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_bp_debug_if = lsu_io_dmem_req_bits_0_bits_uop_bp_debug_if; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_bp_xcpt_if = lsu_io_dmem_req_bits_0_bits_uop_bp_xcpt_if; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_debug_fsrc = lsu_io_dmem_req_bits_0_bits_uop_debug_fsrc; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_uop_debug_tsrc = lsu_io_dmem_req_bits_0_bits_uop_debug_tsrc; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_addr = lsu_io_dmem_req_bits_0_bits_addr; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_data = lsu_io_dmem_req_bits_0_bits_data; // @[tile.scala 239:30]
  assign dcache_io_lsu_req_bits_0_bits_is_hella = lsu_io_dmem_req_bits_0_bits_is_hella; // @[tile.scala 239:30]
  assign dcache_io_lsu_s1_kill_0 = lsu_io_dmem_s1_kill_0; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b1_resolve_mask = lsu_io_dmem_brupdate_b1_resolve_mask; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b1_mispredict_mask = lsu_io_dmem_brupdate_b1_mispredict_mask; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_switch = lsu_io_dmem_brupdate_b2_uop_switch; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_switch_off = lsu_io_dmem_brupdate_b2_uop_switch_off; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_is_unicore = lsu_io_dmem_brupdate_b2_uop_is_unicore; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_shift = lsu_io_dmem_brupdate_b2_uop_shift; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_lrs3_rtype = lsu_io_dmem_brupdate_b2_uop_lrs3_rtype; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_rflag = lsu_io_dmem_brupdate_b2_uop_rflag; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_wflag = lsu_io_dmem_brupdate_b2_uop_wflag; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_prflag = lsu_io_dmem_brupdate_b2_uop_prflag; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_pwflag = lsu_io_dmem_brupdate_b2_uop_pwflag; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_pflag_busy = lsu_io_dmem_brupdate_b2_uop_pflag_busy; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_stale_pflag = lsu_io_dmem_brupdate_b2_uop_stale_pflag; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_op1_sel = lsu_io_dmem_brupdate_b2_uop_op1_sel; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_op2_sel = lsu_io_dmem_brupdate_b2_uop_op2_sel; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_split_num = lsu_io_dmem_brupdate_b2_uop_split_num; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_self_index = lsu_io_dmem_brupdate_b2_uop_self_index; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_rob_inst_idx = lsu_io_dmem_brupdate_b2_uop_rob_inst_idx; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_address_num = lsu_io_dmem_brupdate_b2_uop_address_num; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_uopc = lsu_io_dmem_brupdate_b2_uop_uopc; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_inst = lsu_io_dmem_brupdate_b2_uop_inst; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_debug_inst = lsu_io_dmem_brupdate_b2_uop_debug_inst; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_is_rvc = lsu_io_dmem_brupdate_b2_uop_is_rvc; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_debug_pc = lsu_io_dmem_brupdate_b2_uop_debug_pc; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_iq_type = lsu_io_dmem_brupdate_b2_uop_iq_type; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_fu_code = lsu_io_dmem_brupdate_b2_uop_fu_code; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_ctrl_br_type = lsu_io_dmem_brupdate_b2_uop_ctrl_br_type; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_ctrl_op1_sel = lsu_io_dmem_brupdate_b2_uop_ctrl_op1_sel; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_ctrl_op2_sel = lsu_io_dmem_brupdate_b2_uop_ctrl_op2_sel; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_ctrl_imm_sel = lsu_io_dmem_brupdate_b2_uop_ctrl_imm_sel; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_ctrl_op_fcn = lsu_io_dmem_brupdate_b2_uop_ctrl_op_fcn; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_ctrl_fcn_dw = lsu_io_dmem_brupdate_b2_uop_ctrl_fcn_dw; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_ctrl_csr_cmd = lsu_io_dmem_brupdate_b2_uop_ctrl_csr_cmd; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_ctrl_is_load = lsu_io_dmem_brupdate_b2_uop_ctrl_is_load; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_ctrl_is_sta = lsu_io_dmem_brupdate_b2_uop_ctrl_is_sta; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_ctrl_is_std = lsu_io_dmem_brupdate_b2_uop_ctrl_is_std; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_ctrl_op3_sel = lsu_io_dmem_brupdate_b2_uop_ctrl_op3_sel; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_iw_state = lsu_io_dmem_brupdate_b2_uop_iw_state; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_iw_p1_poisoned = lsu_io_dmem_brupdate_b2_uop_iw_p1_poisoned; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_iw_p2_poisoned = lsu_io_dmem_brupdate_b2_uop_iw_p2_poisoned; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_is_br = lsu_io_dmem_brupdate_b2_uop_is_br; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_is_jalr = lsu_io_dmem_brupdate_b2_uop_is_jalr; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_is_jal = lsu_io_dmem_brupdate_b2_uop_is_jal; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_is_sfb = lsu_io_dmem_brupdate_b2_uop_is_sfb; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_br_mask = lsu_io_dmem_brupdate_b2_uop_br_mask; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_br_tag = lsu_io_dmem_brupdate_b2_uop_br_tag; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_ftq_idx = lsu_io_dmem_brupdate_b2_uop_ftq_idx; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_edge_inst = lsu_io_dmem_brupdate_b2_uop_edge_inst; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_pc_lob = lsu_io_dmem_brupdate_b2_uop_pc_lob; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_taken = lsu_io_dmem_brupdate_b2_uop_taken; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_imm_packed = lsu_io_dmem_brupdate_b2_uop_imm_packed; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_csr_addr = lsu_io_dmem_brupdate_b2_uop_csr_addr; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_rob_idx = lsu_io_dmem_brupdate_b2_uop_rob_idx; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_ldq_idx = lsu_io_dmem_brupdate_b2_uop_ldq_idx; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_stq_idx = lsu_io_dmem_brupdate_b2_uop_stq_idx; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_rxq_idx = lsu_io_dmem_brupdate_b2_uop_rxq_idx; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_pdst = lsu_io_dmem_brupdate_b2_uop_pdst; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_prs1 = lsu_io_dmem_brupdate_b2_uop_prs1; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_prs2 = lsu_io_dmem_brupdate_b2_uop_prs2; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_prs3 = lsu_io_dmem_brupdate_b2_uop_prs3; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_ppred = lsu_io_dmem_brupdate_b2_uop_ppred; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_prs1_busy = lsu_io_dmem_brupdate_b2_uop_prs1_busy; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_prs2_busy = lsu_io_dmem_brupdate_b2_uop_prs2_busy; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_prs3_busy = lsu_io_dmem_brupdate_b2_uop_prs3_busy; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_ppred_busy = lsu_io_dmem_brupdate_b2_uop_ppred_busy; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_stale_pdst = lsu_io_dmem_brupdate_b2_uop_stale_pdst; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_exception = lsu_io_dmem_brupdate_b2_uop_exception; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_exc_cause = lsu_io_dmem_brupdate_b2_uop_exc_cause; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_bypassable = lsu_io_dmem_brupdate_b2_uop_bypassable; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_mem_cmd = lsu_io_dmem_brupdate_b2_uop_mem_cmd; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_mem_size = lsu_io_dmem_brupdate_b2_uop_mem_size; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_mem_signed = lsu_io_dmem_brupdate_b2_uop_mem_signed; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_is_fence = lsu_io_dmem_brupdate_b2_uop_is_fence; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_is_fencei = lsu_io_dmem_brupdate_b2_uop_is_fencei; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_is_amo = lsu_io_dmem_brupdate_b2_uop_is_amo; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_uses_ldq = lsu_io_dmem_brupdate_b2_uop_uses_ldq; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_uses_stq = lsu_io_dmem_brupdate_b2_uop_uses_stq; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_is_sys_pc2epc = lsu_io_dmem_brupdate_b2_uop_is_sys_pc2epc; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_is_unique = lsu_io_dmem_brupdate_b2_uop_is_unique; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_flush_on_commit = lsu_io_dmem_brupdate_b2_uop_flush_on_commit; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_ldst_is_rs1 = lsu_io_dmem_brupdate_b2_uop_ldst_is_rs1; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_ldst = lsu_io_dmem_brupdate_b2_uop_ldst; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_lrs1 = lsu_io_dmem_brupdate_b2_uop_lrs1; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_lrs2 = lsu_io_dmem_brupdate_b2_uop_lrs2; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_lrs3 = lsu_io_dmem_brupdate_b2_uop_lrs3; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_ldst_val = lsu_io_dmem_brupdate_b2_uop_ldst_val; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_dst_rtype = lsu_io_dmem_brupdate_b2_uop_dst_rtype; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_lrs1_rtype = lsu_io_dmem_brupdate_b2_uop_lrs1_rtype; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_lrs2_rtype = lsu_io_dmem_brupdate_b2_uop_lrs2_rtype; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_frs3_en = lsu_io_dmem_brupdate_b2_uop_frs3_en; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_fp_val = lsu_io_dmem_brupdate_b2_uop_fp_val; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_fp_single = lsu_io_dmem_brupdate_b2_uop_fp_single; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_xcpt_pf_if = lsu_io_dmem_brupdate_b2_uop_xcpt_pf_if; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_xcpt_ae_if = lsu_io_dmem_brupdate_b2_uop_xcpt_ae_if; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_xcpt_ma_if = lsu_io_dmem_brupdate_b2_uop_xcpt_ma_if; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_bp_debug_if = lsu_io_dmem_brupdate_b2_uop_bp_debug_if; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_bp_xcpt_if = lsu_io_dmem_brupdate_b2_uop_bp_xcpt_if; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_debug_fsrc = lsu_io_dmem_brupdate_b2_uop_debug_fsrc; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_uop_debug_tsrc = lsu_io_dmem_brupdate_b2_uop_debug_tsrc; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_valid = lsu_io_dmem_brupdate_b2_valid; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_mispredict = lsu_io_dmem_brupdate_b2_mispredict; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_taken = lsu_io_dmem_brupdate_b2_taken; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_cfi_type = lsu_io_dmem_brupdate_b2_cfi_type; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_pc_sel = lsu_io_dmem_brupdate_b2_pc_sel; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_jalr_target = lsu_io_dmem_brupdate_b2_jalr_target; // @[tile.scala 239:30]
  assign dcache_io_lsu_brupdate_b2_target_offset = lsu_io_dmem_brupdate_b2_target_offset; // @[tile.scala 239:30]
  assign dcache_io_lsu_exception = lsu_io_dmem_exception; // @[tile.scala 239:30]
  assign dcache_io_lsu_rob_pnr_idx = lsu_io_dmem_rob_pnr_idx; // @[tile.scala 239:30]
  assign dcache_io_lsu_rob_head_idx = lsu_io_dmem_rob_head_idx; // @[tile.scala 239:30]
  assign dcache_io_lsu_release_ready = lsu_io_dmem_release_ready; // @[tile.scala 239:30]
  assign dcache_io_lsu_force_order = lsu_io_dmem_force_order; // @[tile.scala 239:30]
  assign frontend_clock = clock;
  assign frontend_reset = reset;
  assign frontend_auto_icache_master_out_a_ready = tlMasterXbar_auto_in_1_a_ready; // @[LazyModule.scala 296:16]
  assign frontend_auto_icache_master_out_d_valid = tlMasterXbar_auto_in_1_d_valid; // @[LazyModule.scala 296:16]
  assign frontend_auto_icache_master_out_d_bits_opcode = tlMasterXbar_auto_in_1_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign frontend_auto_icache_master_out_d_bits_param = tlMasterXbar_auto_in_1_d_bits_param; // @[LazyModule.scala 296:16]
  assign frontend_auto_icache_master_out_d_bits_size = tlMasterXbar_auto_in_1_d_bits_size; // @[LazyModule.scala 296:16]
  assign frontend_auto_icache_master_out_d_bits_source = tlMasterXbar_auto_in_1_d_bits_source; // @[LazyModule.scala 296:16]
  assign frontend_auto_icache_master_out_d_bits_sink = tlMasterXbar_auto_in_1_d_bits_sink; // @[LazyModule.scala 296:16]
  assign frontend_auto_icache_master_out_d_bits_denied = tlMasterXbar_auto_in_1_d_bits_denied; // @[LazyModule.scala 296:16]
  assign frontend_auto_icache_master_out_d_bits_data = tlMasterXbar_auto_in_1_d_bits_data; // @[LazyModule.scala 296:16]
  assign frontend_auto_icache_master_out_d_bits_corrupt = tlMasterXbar_auto_in_1_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign frontend_auto_reset_vector_sink_in = broadcast_1_auto_out_1; // @[LazyModule.scala 298:16]
  assign frontend_io_cpu_fetchpacket_ready = core_io_ifu_fetchpacket_ready; // @[tile.scala 177:32]
  assign frontend_io_cpu_get_pc_0_ftq_idx = core_io_ifu_get_pc_0_ftq_idx; // @[tile.scala 177:32]
  assign frontend_io_cpu_get_pc_1_ftq_idx = core_io_ifu_get_pc_1_ftq_idx; // @[tile.scala 177:32]
  assign frontend_io_cpu_get_pc_2_ftq_idx = core_io_ifu_get_pc_2_ftq_idx; // @[tile.scala 177:32]
  assign frontend_io_cpu_get_pc_3_ftq_idx = core_io_ifu_get_pc_3_ftq_idx; // @[tile.scala 177:32]
  assign frontend_io_cpu_debug_ftq_idx_0 = core_io_ifu_debug_ftq_idx_0; // @[tile.scala 177:32]
  assign frontend_io_cpu_debug_ftq_idx_1 = core_io_ifu_debug_ftq_idx_1; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_debug = core_io_ifu_status_debug; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_cease = core_io_ifu_status_cease; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_wfi = core_io_ifu_status_wfi; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_isa = core_io_ifu_status_isa; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_dprv = core_io_ifu_status_dprv; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_prv = core_io_ifu_status_prv; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_sd = core_io_ifu_status_sd; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_zero2 = core_io_ifu_status_zero2; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_sxl = core_io_ifu_status_sxl; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_uxl = core_io_ifu_status_uxl; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_sd_rv32 = core_io_ifu_status_sd_rv32; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_zero1 = core_io_ifu_status_zero1; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_tsr = core_io_ifu_status_tsr; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_tw = core_io_ifu_status_tw; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_tvm = core_io_ifu_status_tvm; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_mxr = core_io_ifu_status_mxr; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_sum = core_io_ifu_status_sum; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_mprv = core_io_ifu_status_mprv; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_xs = core_io_ifu_status_xs; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_fs = core_io_ifu_status_fs; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_mpp = core_io_ifu_status_mpp; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_vs = core_io_ifu_status_vs; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_spp = core_io_ifu_status_spp; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_mpie = core_io_ifu_status_mpie; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_hpie = core_io_ifu_status_hpie; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_spie = core_io_ifu_status_spie; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_upie = core_io_ifu_status_upie; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_mie = core_io_ifu_status_mie; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_hie = core_io_ifu_status_hie; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_sie = core_io_ifu_status_sie; // @[tile.scala 177:32]
  assign frontend_io_cpu_status_uie = core_io_ifu_status_uie; // @[tile.scala 177:32]
  assign frontend_io_cpu_sfence_valid = core_io_ifu_sfence_valid; // @[tile.scala 177:32]
  assign frontend_io_cpu_sfence_bits_rs1 = core_io_ifu_sfence_bits_rs1; // @[tile.scala 177:32]
  assign frontend_io_cpu_sfence_bits_rs2 = core_io_ifu_sfence_bits_rs2; // @[tile.scala 177:32]
  assign frontend_io_cpu_sfence_bits_addr = core_io_ifu_sfence_bits_addr; // @[tile.scala 177:32]
  assign frontend_io_cpu_sfence_bits_asid = core_io_ifu_sfence_bits_asid; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b1_resolve_mask = core_io_ifu_brupdate_b1_resolve_mask; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b1_mispredict_mask = core_io_ifu_brupdate_b1_mispredict_mask; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_switch = core_io_ifu_brupdate_b2_uop_switch; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_switch_off = core_io_ifu_brupdate_b2_uop_switch_off; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_is_unicore = core_io_ifu_brupdate_b2_uop_is_unicore; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_shift = core_io_ifu_brupdate_b2_uop_shift; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_lrs3_rtype = core_io_ifu_brupdate_b2_uop_lrs3_rtype; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_rflag = core_io_ifu_brupdate_b2_uop_rflag; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_wflag = core_io_ifu_brupdate_b2_uop_wflag; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_prflag = core_io_ifu_brupdate_b2_uop_prflag; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_pwflag = core_io_ifu_brupdate_b2_uop_pwflag; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_pflag_busy = core_io_ifu_brupdate_b2_uop_pflag_busy; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_stale_pflag = core_io_ifu_brupdate_b2_uop_stale_pflag; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_op1_sel = core_io_ifu_brupdate_b2_uop_op1_sel; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_op2_sel = core_io_ifu_brupdate_b2_uop_op2_sel; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_split_num = core_io_ifu_brupdate_b2_uop_split_num; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_self_index = core_io_ifu_brupdate_b2_uop_self_index; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_rob_inst_idx = core_io_ifu_brupdate_b2_uop_rob_inst_idx; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_address_num = core_io_ifu_brupdate_b2_uop_address_num; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_uopc = core_io_ifu_brupdate_b2_uop_uopc; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_inst = core_io_ifu_brupdate_b2_uop_inst; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_debug_inst = core_io_ifu_brupdate_b2_uop_debug_inst; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_is_rvc = core_io_ifu_brupdate_b2_uop_is_rvc; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_debug_pc = core_io_ifu_brupdate_b2_uop_debug_pc; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_iq_type = core_io_ifu_brupdate_b2_uop_iq_type; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_fu_code = core_io_ifu_brupdate_b2_uop_fu_code; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_ctrl_br_type = core_io_ifu_brupdate_b2_uop_ctrl_br_type; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_ctrl_op1_sel = core_io_ifu_brupdate_b2_uop_ctrl_op1_sel; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_ctrl_op2_sel = core_io_ifu_brupdate_b2_uop_ctrl_op2_sel; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_ctrl_imm_sel = core_io_ifu_brupdate_b2_uop_ctrl_imm_sel; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_ctrl_op_fcn = core_io_ifu_brupdate_b2_uop_ctrl_op_fcn; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_ctrl_fcn_dw = core_io_ifu_brupdate_b2_uop_ctrl_fcn_dw; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_ctrl_csr_cmd = core_io_ifu_brupdate_b2_uop_ctrl_csr_cmd; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_ctrl_is_load = core_io_ifu_brupdate_b2_uop_ctrl_is_load; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_ctrl_is_sta = core_io_ifu_brupdate_b2_uop_ctrl_is_sta; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_ctrl_is_std = core_io_ifu_brupdate_b2_uop_ctrl_is_std; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_ctrl_op3_sel = core_io_ifu_brupdate_b2_uop_ctrl_op3_sel; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_iw_state = core_io_ifu_brupdate_b2_uop_iw_state; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_iw_p1_poisoned = core_io_ifu_brupdate_b2_uop_iw_p1_poisoned; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_iw_p2_poisoned = core_io_ifu_brupdate_b2_uop_iw_p2_poisoned; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_is_br = core_io_ifu_brupdate_b2_uop_is_br; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_is_jalr = core_io_ifu_brupdate_b2_uop_is_jalr; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_is_jal = core_io_ifu_brupdate_b2_uop_is_jal; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_is_sfb = core_io_ifu_brupdate_b2_uop_is_sfb; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_br_mask = core_io_ifu_brupdate_b2_uop_br_mask; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_br_tag = core_io_ifu_brupdate_b2_uop_br_tag; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_ftq_idx = core_io_ifu_brupdate_b2_uop_ftq_idx; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_edge_inst = core_io_ifu_brupdate_b2_uop_edge_inst; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_pc_lob = core_io_ifu_brupdate_b2_uop_pc_lob; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_taken = core_io_ifu_brupdate_b2_uop_taken; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_imm_packed = core_io_ifu_brupdate_b2_uop_imm_packed; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_csr_addr = core_io_ifu_brupdate_b2_uop_csr_addr; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_rob_idx = core_io_ifu_brupdate_b2_uop_rob_idx; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_ldq_idx = core_io_ifu_brupdate_b2_uop_ldq_idx; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_stq_idx = core_io_ifu_brupdate_b2_uop_stq_idx; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_rxq_idx = core_io_ifu_brupdate_b2_uop_rxq_idx; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_pdst = core_io_ifu_brupdate_b2_uop_pdst; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_prs1 = core_io_ifu_brupdate_b2_uop_prs1; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_prs2 = core_io_ifu_brupdate_b2_uop_prs2; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_prs3 = core_io_ifu_brupdate_b2_uop_prs3; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_ppred = core_io_ifu_brupdate_b2_uop_ppred; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_prs1_busy = core_io_ifu_brupdate_b2_uop_prs1_busy; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_prs2_busy = core_io_ifu_brupdate_b2_uop_prs2_busy; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_prs3_busy = core_io_ifu_brupdate_b2_uop_prs3_busy; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_ppred_busy = core_io_ifu_brupdate_b2_uop_ppred_busy; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_stale_pdst = core_io_ifu_brupdate_b2_uop_stale_pdst; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_exception = core_io_ifu_brupdate_b2_uop_exception; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_exc_cause = core_io_ifu_brupdate_b2_uop_exc_cause; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_bypassable = core_io_ifu_brupdate_b2_uop_bypassable; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_mem_cmd = core_io_ifu_brupdate_b2_uop_mem_cmd; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_mem_size = core_io_ifu_brupdate_b2_uop_mem_size; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_mem_signed = core_io_ifu_brupdate_b2_uop_mem_signed; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_is_fence = core_io_ifu_brupdate_b2_uop_is_fence; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_is_fencei = core_io_ifu_brupdate_b2_uop_is_fencei; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_is_amo = core_io_ifu_brupdate_b2_uop_is_amo; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_uses_ldq = core_io_ifu_brupdate_b2_uop_uses_ldq; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_uses_stq = core_io_ifu_brupdate_b2_uop_uses_stq; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_is_sys_pc2epc = core_io_ifu_brupdate_b2_uop_is_sys_pc2epc; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_is_unique = core_io_ifu_brupdate_b2_uop_is_unique; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_flush_on_commit = core_io_ifu_brupdate_b2_uop_flush_on_commit; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_ldst_is_rs1 = core_io_ifu_brupdate_b2_uop_ldst_is_rs1; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_ldst = core_io_ifu_brupdate_b2_uop_ldst; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_lrs1 = core_io_ifu_brupdate_b2_uop_lrs1; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_lrs2 = core_io_ifu_brupdate_b2_uop_lrs2; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_lrs3 = core_io_ifu_brupdate_b2_uop_lrs3; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_ldst_val = core_io_ifu_brupdate_b2_uop_ldst_val; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_dst_rtype = core_io_ifu_brupdate_b2_uop_dst_rtype; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_lrs1_rtype = core_io_ifu_brupdate_b2_uop_lrs1_rtype; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_lrs2_rtype = core_io_ifu_brupdate_b2_uop_lrs2_rtype; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_frs3_en = core_io_ifu_brupdate_b2_uop_frs3_en; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_fp_val = core_io_ifu_brupdate_b2_uop_fp_val; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_fp_single = core_io_ifu_brupdate_b2_uop_fp_single; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_xcpt_pf_if = core_io_ifu_brupdate_b2_uop_xcpt_pf_if; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_xcpt_ae_if = core_io_ifu_brupdate_b2_uop_xcpt_ae_if; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_xcpt_ma_if = core_io_ifu_brupdate_b2_uop_xcpt_ma_if; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_bp_debug_if = core_io_ifu_brupdate_b2_uop_bp_debug_if; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_bp_xcpt_if = core_io_ifu_brupdate_b2_uop_bp_xcpt_if; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_debug_fsrc = core_io_ifu_brupdate_b2_uop_debug_fsrc; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_uop_debug_tsrc = core_io_ifu_brupdate_b2_uop_debug_tsrc; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_valid = core_io_ifu_brupdate_b2_valid; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_mispredict = core_io_ifu_brupdate_b2_mispredict; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_taken = core_io_ifu_brupdate_b2_taken; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_cfi_type = core_io_ifu_brupdate_b2_cfi_type; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_pc_sel = core_io_ifu_brupdate_b2_pc_sel; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_jalr_target = core_io_ifu_brupdate_b2_jalr_target; // @[tile.scala 177:32]
  assign frontend_io_cpu_brupdate_b2_target_offset = core_io_ifu_brupdate_b2_target_offset; // @[tile.scala 177:32]
  assign frontend_io_cpu_redirect_flush = core_io_ifu_redirect_flush; // @[tile.scala 177:32]
  assign frontend_io_cpu_redirect_val = core_io_ifu_redirect_val; // @[tile.scala 177:32]
  assign frontend_io_cpu_redirect_pc = core_io_ifu_redirect_pc; // @[tile.scala 177:32]
  assign frontend_io_cpu_redirect_ftq_idx = core_io_ifu_redirect_ftq_idx; // @[tile.scala 177:32]
  assign frontend_io_cpu_redirect_ghist_old_history = core_io_ifu_redirect_ghist_old_history; // @[tile.scala 177:32]
  assign frontend_io_cpu_redirect_ghist_current_saw_branch_not_taken =
    core_io_ifu_redirect_ghist_current_saw_branch_not_taken; // @[tile.scala 177:32]
  assign frontend_io_cpu_redirect_ghist_new_saw_branch_not_taken = core_io_ifu_redirect_ghist_new_saw_branch_not_taken; // @[tile.scala 177:32]
  assign frontend_io_cpu_redirect_ghist_new_saw_branch_taken = core_io_ifu_redirect_ghist_new_saw_branch_taken; // @[tile.scala 177:32]
  assign frontend_io_cpu_redirect_ghist_ras_idx = core_io_ifu_redirect_ghist_ras_idx; // @[tile.scala 177:32]
  assign frontend_io_cpu_commit_valid = core_io_ifu_commit_valid; // @[tile.scala 177:32]
  assign frontend_io_cpu_commit_bits = core_io_ifu_commit_bits; // @[tile.scala 177:32]
  assign frontend_io_cpu_flush_icache = core_io_ifu_flush_icache; // @[tile.scala 177:32]
  assign frontend_io_cpu_is_unicore = core_io_ifu_is_unicore; // @[tile.scala 177:32]
  assign frontend_io_ptw_req_ready = ptw_io_requestor_1_req_ready; // @[tile.scala 232:20]
  assign frontend_io_ptw_resp_valid = ptw_io_requestor_1_resp_valid; // @[tile.scala 232:20]
  assign frontend_io_ptw_resp_bits_ae = ptw_io_requestor_1_resp_bits_ae; // @[tile.scala 232:20]
  assign frontend_io_ptw_resp_bits_pte_ppn = ptw_io_requestor_1_resp_bits_pte_ppn; // @[tile.scala 232:20]
  assign frontend_io_ptw_resp_bits_pte_reserved_for_software = ptw_io_requestor_1_resp_bits_pte_reserved_for_software; // @[tile.scala 232:20]
  assign frontend_io_ptw_resp_bits_pte_d = ptw_io_requestor_1_resp_bits_pte_d; // @[tile.scala 232:20]
  assign frontend_io_ptw_resp_bits_pte_a = ptw_io_requestor_1_resp_bits_pte_a; // @[tile.scala 232:20]
  assign frontend_io_ptw_resp_bits_pte_g = ptw_io_requestor_1_resp_bits_pte_g; // @[tile.scala 232:20]
  assign frontend_io_ptw_resp_bits_pte_u = ptw_io_requestor_1_resp_bits_pte_u; // @[tile.scala 232:20]
  assign frontend_io_ptw_resp_bits_pte_x = ptw_io_requestor_1_resp_bits_pte_x; // @[tile.scala 232:20]
  assign frontend_io_ptw_resp_bits_pte_w = ptw_io_requestor_1_resp_bits_pte_w; // @[tile.scala 232:20]
  assign frontend_io_ptw_resp_bits_pte_r = ptw_io_requestor_1_resp_bits_pte_r; // @[tile.scala 232:20]
  assign frontend_io_ptw_resp_bits_pte_v = ptw_io_requestor_1_resp_bits_pte_v; // @[tile.scala 232:20]
  assign frontend_io_ptw_resp_bits_level = ptw_io_requestor_1_resp_bits_level; // @[tile.scala 232:20]
  assign frontend_io_ptw_resp_bits_fragmented_superpage = ptw_io_requestor_1_resp_bits_fragmented_superpage; // @[tile.scala 232:20]
  assign frontend_io_ptw_resp_bits_homogeneous = ptw_io_requestor_1_resp_bits_homogeneous; // @[tile.scala 232:20]
  assign frontend_io_ptw_ptbr_mode = ptw_io_requestor_1_ptbr_mode; // @[tile.scala 232:20]
  assign frontend_io_ptw_ptbr_asid = ptw_io_requestor_1_ptbr_asid; // @[tile.scala 232:20]
  assign frontend_io_ptw_ptbr_ppn = ptw_io_requestor_1_ptbr_ppn; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_debug = ptw_io_requestor_1_status_debug; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_cease = ptw_io_requestor_1_status_cease; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_wfi = ptw_io_requestor_1_status_wfi; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_isa = ptw_io_requestor_1_status_isa; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_dprv = ptw_io_requestor_1_status_dprv; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_prv = ptw_io_requestor_1_status_prv; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_sd = ptw_io_requestor_1_status_sd; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_zero2 = ptw_io_requestor_1_status_zero2; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_sxl = ptw_io_requestor_1_status_sxl; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_uxl = ptw_io_requestor_1_status_uxl; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_sd_rv32 = ptw_io_requestor_1_status_sd_rv32; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_zero1 = ptw_io_requestor_1_status_zero1; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_tsr = ptw_io_requestor_1_status_tsr; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_tw = ptw_io_requestor_1_status_tw; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_tvm = ptw_io_requestor_1_status_tvm; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_mxr = ptw_io_requestor_1_status_mxr; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_sum = ptw_io_requestor_1_status_sum; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_mprv = ptw_io_requestor_1_status_mprv; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_xs = ptw_io_requestor_1_status_xs; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_fs = ptw_io_requestor_1_status_fs; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_mpp = ptw_io_requestor_1_status_mpp; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_vs = ptw_io_requestor_1_status_vs; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_spp = ptw_io_requestor_1_status_spp; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_mpie = ptw_io_requestor_1_status_mpie; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_hpie = ptw_io_requestor_1_status_hpie; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_spie = ptw_io_requestor_1_status_spie; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_upie = ptw_io_requestor_1_status_upie; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_mie = ptw_io_requestor_1_status_mie; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_hie = ptw_io_requestor_1_status_hie; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_sie = ptw_io_requestor_1_status_sie; // @[tile.scala 232:20]
  assign frontend_io_ptw_status_uie = ptw_io_requestor_1_status_uie; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_0_cfg_l = ptw_io_requestor_1_pmp_0_cfg_l; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_0_cfg_res = ptw_io_requestor_1_pmp_0_cfg_res; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_0_cfg_a = ptw_io_requestor_1_pmp_0_cfg_a; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_0_cfg_x = ptw_io_requestor_1_pmp_0_cfg_x; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_0_cfg_w = ptw_io_requestor_1_pmp_0_cfg_w; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_0_cfg_r = ptw_io_requestor_1_pmp_0_cfg_r; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_0_addr = ptw_io_requestor_1_pmp_0_addr; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_0_mask = ptw_io_requestor_1_pmp_0_mask; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_1_cfg_l = ptw_io_requestor_1_pmp_1_cfg_l; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_1_cfg_res = ptw_io_requestor_1_pmp_1_cfg_res; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_1_cfg_a = ptw_io_requestor_1_pmp_1_cfg_a; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_1_cfg_x = ptw_io_requestor_1_pmp_1_cfg_x; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_1_cfg_w = ptw_io_requestor_1_pmp_1_cfg_w; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_1_cfg_r = ptw_io_requestor_1_pmp_1_cfg_r; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_1_addr = ptw_io_requestor_1_pmp_1_addr; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_1_mask = ptw_io_requestor_1_pmp_1_mask; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_2_cfg_l = ptw_io_requestor_1_pmp_2_cfg_l; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_2_cfg_res = ptw_io_requestor_1_pmp_2_cfg_res; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_2_cfg_a = ptw_io_requestor_1_pmp_2_cfg_a; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_2_cfg_x = ptw_io_requestor_1_pmp_2_cfg_x; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_2_cfg_w = ptw_io_requestor_1_pmp_2_cfg_w; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_2_cfg_r = ptw_io_requestor_1_pmp_2_cfg_r; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_2_addr = ptw_io_requestor_1_pmp_2_addr; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_2_mask = ptw_io_requestor_1_pmp_2_mask; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_3_cfg_l = ptw_io_requestor_1_pmp_3_cfg_l; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_3_cfg_res = ptw_io_requestor_1_pmp_3_cfg_res; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_3_cfg_a = ptw_io_requestor_1_pmp_3_cfg_a; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_3_cfg_x = ptw_io_requestor_1_pmp_3_cfg_x; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_3_cfg_w = ptw_io_requestor_1_pmp_3_cfg_w; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_3_cfg_r = ptw_io_requestor_1_pmp_3_cfg_r; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_3_addr = ptw_io_requestor_1_pmp_3_addr; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_3_mask = ptw_io_requestor_1_pmp_3_mask; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_4_cfg_l = ptw_io_requestor_1_pmp_4_cfg_l; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_4_cfg_res = ptw_io_requestor_1_pmp_4_cfg_res; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_4_cfg_a = ptw_io_requestor_1_pmp_4_cfg_a; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_4_cfg_x = ptw_io_requestor_1_pmp_4_cfg_x; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_4_cfg_w = ptw_io_requestor_1_pmp_4_cfg_w; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_4_cfg_r = ptw_io_requestor_1_pmp_4_cfg_r; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_4_addr = ptw_io_requestor_1_pmp_4_addr; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_4_mask = ptw_io_requestor_1_pmp_4_mask; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_5_cfg_l = ptw_io_requestor_1_pmp_5_cfg_l; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_5_cfg_res = ptw_io_requestor_1_pmp_5_cfg_res; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_5_cfg_a = ptw_io_requestor_1_pmp_5_cfg_a; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_5_cfg_x = ptw_io_requestor_1_pmp_5_cfg_x; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_5_cfg_w = ptw_io_requestor_1_pmp_5_cfg_w; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_5_cfg_r = ptw_io_requestor_1_pmp_5_cfg_r; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_5_addr = ptw_io_requestor_1_pmp_5_addr; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_5_mask = ptw_io_requestor_1_pmp_5_mask; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_6_cfg_l = ptw_io_requestor_1_pmp_6_cfg_l; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_6_cfg_res = ptw_io_requestor_1_pmp_6_cfg_res; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_6_cfg_a = ptw_io_requestor_1_pmp_6_cfg_a; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_6_cfg_x = ptw_io_requestor_1_pmp_6_cfg_x; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_6_cfg_w = ptw_io_requestor_1_pmp_6_cfg_w; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_6_cfg_r = ptw_io_requestor_1_pmp_6_cfg_r; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_6_addr = ptw_io_requestor_1_pmp_6_addr; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_6_mask = ptw_io_requestor_1_pmp_6_mask; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_7_cfg_l = ptw_io_requestor_1_pmp_7_cfg_l; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_7_cfg_res = ptw_io_requestor_1_pmp_7_cfg_res; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_7_cfg_a = ptw_io_requestor_1_pmp_7_cfg_a; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_7_cfg_x = ptw_io_requestor_1_pmp_7_cfg_x; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_7_cfg_w = ptw_io_requestor_1_pmp_7_cfg_w; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_7_cfg_r = ptw_io_requestor_1_pmp_7_cfg_r; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_7_addr = ptw_io_requestor_1_pmp_7_addr; // @[tile.scala 232:20]
  assign frontend_io_ptw_pmp_7_mask = ptw_io_requestor_1_pmp_7_mask; // @[tile.scala 232:20]
  assign frontend_io_ptw_customCSRs_csrs_0_wen = ptw_io_requestor_1_customCSRs_csrs_0_wen; // @[tile.scala 232:20]
  assign frontend_io_ptw_customCSRs_csrs_0_wdata = ptw_io_requestor_1_customCSRs_csrs_0_wdata; // @[tile.scala 232:20]
  assign frontend_io_ptw_customCSRs_csrs_0_value = ptw_io_requestor_1_customCSRs_csrs_0_value; // @[tile.scala 232:20]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_hartid = broadcast_auto_out; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign core_io_interrupts_debug = intXbar_auto_int_out_0; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign core_io_interrupts_mtip = intXbar_auto_int_out_2; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign core_io_interrupts_msip = intXbar_auto_int_out_1; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign core_io_interrupts_meip = intXbar_auto_int_out_3; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign core_io_interrupts_seip = intXbar_auto_int_out_4; // @[Nodes.scala 1210:84 LazyModule.scala 296:16]
  assign core_io_ifu_fetchpacket_valid = frontend_io_cpu_fetchpacket_valid; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_valid = frontend_io_cpu_fetchpacket_bits_uops_0_valid; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_switch = frontend_io_cpu_fetchpacket_bits_uops_0_bits_switch; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_switch_off = frontend_io_cpu_fetchpacket_bits_uops_0_bits_switch_off; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_is_unicore = frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_unicore; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_shift = frontend_io_cpu_fetchpacket_bits_uops_0_bits_shift; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_lrs3_rtype = frontend_io_cpu_fetchpacket_bits_uops_0_bits_lrs3_rtype; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_rflag = frontend_io_cpu_fetchpacket_bits_uops_0_bits_rflag; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_wflag = frontend_io_cpu_fetchpacket_bits_uops_0_bits_wflag; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_prflag = frontend_io_cpu_fetchpacket_bits_uops_0_bits_prflag; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_pwflag = frontend_io_cpu_fetchpacket_bits_uops_0_bits_pwflag; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_pflag_busy = frontend_io_cpu_fetchpacket_bits_uops_0_bits_pflag_busy; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_stale_pflag = frontend_io_cpu_fetchpacket_bits_uops_0_bits_stale_pflag
    ; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_op1_sel = frontend_io_cpu_fetchpacket_bits_uops_0_bits_op1_sel; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_op2_sel = frontend_io_cpu_fetchpacket_bits_uops_0_bits_op2_sel; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_split_num = frontend_io_cpu_fetchpacket_bits_uops_0_bits_split_num; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_self_index = frontend_io_cpu_fetchpacket_bits_uops_0_bits_self_index; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_rob_inst_idx =
    frontend_io_cpu_fetchpacket_bits_uops_0_bits_rob_inst_idx; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_address_num = frontend_io_cpu_fetchpacket_bits_uops_0_bits_address_num
    ; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_uopc = frontend_io_cpu_fetchpacket_bits_uops_0_bits_uopc; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_inst = frontend_io_cpu_fetchpacket_bits_uops_0_bits_inst; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_debug_inst = frontend_io_cpu_fetchpacket_bits_uops_0_bits_debug_inst; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_is_rvc = frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_rvc; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_debug_pc = frontend_io_cpu_fetchpacket_bits_uops_0_bits_debug_pc; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_iq_type = frontend_io_cpu_fetchpacket_bits_uops_0_bits_iq_type; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_fu_code = frontend_io_cpu_fetchpacket_bits_uops_0_bits_fu_code; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_br_type =
    frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_br_type; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_op1_sel =
    frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_op1_sel; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_op2_sel =
    frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_op2_sel; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_imm_sel =
    frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_imm_sel; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_op_fcn = frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_op_fcn
    ; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_fcn_dw = frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_fcn_dw
    ; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_csr_cmd =
    frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_csr_cmd; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_is_load =
    frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_is_load; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_is_sta = frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_is_sta
    ; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_is_std = frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_is_std
    ; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_ctrl_op3_sel =
    frontend_io_cpu_fetchpacket_bits_uops_0_bits_ctrl_op3_sel; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_iw_state = frontend_io_cpu_fetchpacket_bits_uops_0_bits_iw_state; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_iw_p1_poisoned =
    frontend_io_cpu_fetchpacket_bits_uops_0_bits_iw_p1_poisoned; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_iw_p2_poisoned =
    frontend_io_cpu_fetchpacket_bits_uops_0_bits_iw_p2_poisoned; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_is_br = frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_br; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_is_jalr = frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_jalr; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_is_jal = frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_jal; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_is_sfb = frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_sfb; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_br_mask = frontend_io_cpu_fetchpacket_bits_uops_0_bits_br_mask; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_br_tag = frontend_io_cpu_fetchpacket_bits_uops_0_bits_br_tag; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_ftq_idx = frontend_io_cpu_fetchpacket_bits_uops_0_bits_ftq_idx; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_edge_inst = frontend_io_cpu_fetchpacket_bits_uops_0_bits_edge_inst; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_pc_lob = frontend_io_cpu_fetchpacket_bits_uops_0_bits_pc_lob; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_taken = frontend_io_cpu_fetchpacket_bits_uops_0_bits_taken; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_imm_packed = frontend_io_cpu_fetchpacket_bits_uops_0_bits_imm_packed; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_csr_addr = frontend_io_cpu_fetchpacket_bits_uops_0_bits_csr_addr; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_rob_idx = frontend_io_cpu_fetchpacket_bits_uops_0_bits_rob_idx; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_ldq_idx = frontend_io_cpu_fetchpacket_bits_uops_0_bits_ldq_idx; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_stq_idx = frontend_io_cpu_fetchpacket_bits_uops_0_bits_stq_idx; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_rxq_idx = frontend_io_cpu_fetchpacket_bits_uops_0_bits_rxq_idx; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_pdst = frontend_io_cpu_fetchpacket_bits_uops_0_bits_pdst; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_prs1 = frontend_io_cpu_fetchpacket_bits_uops_0_bits_prs1; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_prs2 = frontend_io_cpu_fetchpacket_bits_uops_0_bits_prs2; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_prs3 = frontend_io_cpu_fetchpacket_bits_uops_0_bits_prs3; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_ppred = frontend_io_cpu_fetchpacket_bits_uops_0_bits_ppred; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_prs1_busy = frontend_io_cpu_fetchpacket_bits_uops_0_bits_prs1_busy; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_prs2_busy = frontend_io_cpu_fetchpacket_bits_uops_0_bits_prs2_busy; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_prs3_busy = frontend_io_cpu_fetchpacket_bits_uops_0_bits_prs3_busy; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_ppred_busy = frontend_io_cpu_fetchpacket_bits_uops_0_bits_ppred_busy; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_stale_pdst = frontend_io_cpu_fetchpacket_bits_uops_0_bits_stale_pdst; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_exception = frontend_io_cpu_fetchpacket_bits_uops_0_bits_exception; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_exc_cause = frontend_io_cpu_fetchpacket_bits_uops_0_bits_exc_cause; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_bypassable = frontend_io_cpu_fetchpacket_bits_uops_0_bits_bypassable; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_mem_cmd = frontend_io_cpu_fetchpacket_bits_uops_0_bits_mem_cmd; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_mem_size = frontend_io_cpu_fetchpacket_bits_uops_0_bits_mem_size; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_mem_signed = frontend_io_cpu_fetchpacket_bits_uops_0_bits_mem_signed; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_is_fence = frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_fence; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_is_fencei = frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_fencei; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_is_amo = frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_amo; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_uses_ldq = frontend_io_cpu_fetchpacket_bits_uops_0_bits_uses_ldq; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_uses_stq = frontend_io_cpu_fetchpacket_bits_uops_0_bits_uses_stq; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_is_sys_pc2epc =
    frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_sys_pc2epc; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_is_unique = frontend_io_cpu_fetchpacket_bits_uops_0_bits_is_unique; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_flush_on_commit =
    frontend_io_cpu_fetchpacket_bits_uops_0_bits_flush_on_commit; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_ldst_is_rs1 = frontend_io_cpu_fetchpacket_bits_uops_0_bits_ldst_is_rs1
    ; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_ldst = frontend_io_cpu_fetchpacket_bits_uops_0_bits_ldst; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_lrs1 = frontend_io_cpu_fetchpacket_bits_uops_0_bits_lrs1; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_lrs2 = frontend_io_cpu_fetchpacket_bits_uops_0_bits_lrs2; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_lrs3 = frontend_io_cpu_fetchpacket_bits_uops_0_bits_lrs3; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_ldst_val = frontend_io_cpu_fetchpacket_bits_uops_0_bits_ldst_val; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_dst_rtype = frontend_io_cpu_fetchpacket_bits_uops_0_bits_dst_rtype; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_lrs1_rtype = frontend_io_cpu_fetchpacket_bits_uops_0_bits_lrs1_rtype; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_lrs2_rtype = frontend_io_cpu_fetchpacket_bits_uops_0_bits_lrs2_rtype; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_frs3_en = frontend_io_cpu_fetchpacket_bits_uops_0_bits_frs3_en; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_fp_val = frontend_io_cpu_fetchpacket_bits_uops_0_bits_fp_val; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_fp_single = frontend_io_cpu_fetchpacket_bits_uops_0_bits_fp_single; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_xcpt_pf_if = frontend_io_cpu_fetchpacket_bits_uops_0_bits_xcpt_pf_if; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_xcpt_ae_if = frontend_io_cpu_fetchpacket_bits_uops_0_bits_xcpt_ae_if; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_xcpt_ma_if = frontend_io_cpu_fetchpacket_bits_uops_0_bits_xcpt_ma_if; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_bp_debug_if = frontend_io_cpu_fetchpacket_bits_uops_0_bits_bp_debug_if
    ; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_bp_xcpt_if = frontend_io_cpu_fetchpacket_bits_uops_0_bits_bp_xcpt_if; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_debug_fsrc = frontend_io_cpu_fetchpacket_bits_uops_0_bits_debug_fsrc; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_0_bits_debug_tsrc = frontend_io_cpu_fetchpacket_bits_uops_0_bits_debug_tsrc; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_valid = frontend_io_cpu_fetchpacket_bits_uops_1_valid; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_switch = frontend_io_cpu_fetchpacket_bits_uops_1_bits_switch; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_switch_off = frontend_io_cpu_fetchpacket_bits_uops_1_bits_switch_off; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_is_unicore = frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_unicore; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_shift = frontend_io_cpu_fetchpacket_bits_uops_1_bits_shift; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_lrs3_rtype = frontend_io_cpu_fetchpacket_bits_uops_1_bits_lrs3_rtype; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_rflag = frontend_io_cpu_fetchpacket_bits_uops_1_bits_rflag; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_wflag = frontend_io_cpu_fetchpacket_bits_uops_1_bits_wflag; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_prflag = frontend_io_cpu_fetchpacket_bits_uops_1_bits_prflag; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_pwflag = frontend_io_cpu_fetchpacket_bits_uops_1_bits_pwflag; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_pflag_busy = frontend_io_cpu_fetchpacket_bits_uops_1_bits_pflag_busy; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_stale_pflag = frontend_io_cpu_fetchpacket_bits_uops_1_bits_stale_pflag
    ; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_op1_sel = frontend_io_cpu_fetchpacket_bits_uops_1_bits_op1_sel; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_op2_sel = frontend_io_cpu_fetchpacket_bits_uops_1_bits_op2_sel; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_split_num = frontend_io_cpu_fetchpacket_bits_uops_1_bits_split_num; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_self_index = frontend_io_cpu_fetchpacket_bits_uops_1_bits_self_index; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_rob_inst_idx =
    frontend_io_cpu_fetchpacket_bits_uops_1_bits_rob_inst_idx; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_address_num = frontend_io_cpu_fetchpacket_bits_uops_1_bits_address_num
    ; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_uopc = frontend_io_cpu_fetchpacket_bits_uops_1_bits_uopc; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_inst = frontend_io_cpu_fetchpacket_bits_uops_1_bits_inst; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_debug_inst = frontend_io_cpu_fetchpacket_bits_uops_1_bits_debug_inst; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_is_rvc = frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_rvc; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_debug_pc = frontend_io_cpu_fetchpacket_bits_uops_1_bits_debug_pc; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_iq_type = frontend_io_cpu_fetchpacket_bits_uops_1_bits_iq_type; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_fu_code = frontend_io_cpu_fetchpacket_bits_uops_1_bits_fu_code; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_br_type =
    frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_br_type; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_op1_sel =
    frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_op1_sel; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_op2_sel =
    frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_op2_sel; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_imm_sel =
    frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_imm_sel; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_op_fcn = frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_op_fcn
    ; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_fcn_dw = frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_fcn_dw
    ; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_csr_cmd =
    frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_csr_cmd; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_is_load =
    frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_is_load; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_is_sta = frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_is_sta
    ; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_is_std = frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_is_std
    ; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_ctrl_op3_sel =
    frontend_io_cpu_fetchpacket_bits_uops_1_bits_ctrl_op3_sel; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_iw_state = frontend_io_cpu_fetchpacket_bits_uops_1_bits_iw_state; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_iw_p1_poisoned =
    frontend_io_cpu_fetchpacket_bits_uops_1_bits_iw_p1_poisoned; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_iw_p2_poisoned =
    frontend_io_cpu_fetchpacket_bits_uops_1_bits_iw_p2_poisoned; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_is_br = frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_br; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_is_jalr = frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_jalr; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_is_jal = frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_jal; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_is_sfb = frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_sfb; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_br_mask = frontend_io_cpu_fetchpacket_bits_uops_1_bits_br_mask; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_br_tag = frontend_io_cpu_fetchpacket_bits_uops_1_bits_br_tag; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_ftq_idx = frontend_io_cpu_fetchpacket_bits_uops_1_bits_ftq_idx; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_edge_inst = frontend_io_cpu_fetchpacket_bits_uops_1_bits_edge_inst; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_pc_lob = frontend_io_cpu_fetchpacket_bits_uops_1_bits_pc_lob; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_taken = frontend_io_cpu_fetchpacket_bits_uops_1_bits_taken; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_imm_packed = frontend_io_cpu_fetchpacket_bits_uops_1_bits_imm_packed; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_csr_addr = frontend_io_cpu_fetchpacket_bits_uops_1_bits_csr_addr; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_rob_idx = frontend_io_cpu_fetchpacket_bits_uops_1_bits_rob_idx; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_ldq_idx = frontend_io_cpu_fetchpacket_bits_uops_1_bits_ldq_idx; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_stq_idx = frontend_io_cpu_fetchpacket_bits_uops_1_bits_stq_idx; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_rxq_idx = frontend_io_cpu_fetchpacket_bits_uops_1_bits_rxq_idx; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_pdst = frontend_io_cpu_fetchpacket_bits_uops_1_bits_pdst; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_prs1 = frontend_io_cpu_fetchpacket_bits_uops_1_bits_prs1; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_prs2 = frontend_io_cpu_fetchpacket_bits_uops_1_bits_prs2; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_prs3 = frontend_io_cpu_fetchpacket_bits_uops_1_bits_prs3; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_ppred = frontend_io_cpu_fetchpacket_bits_uops_1_bits_ppred; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_prs1_busy = frontend_io_cpu_fetchpacket_bits_uops_1_bits_prs1_busy; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_prs2_busy = frontend_io_cpu_fetchpacket_bits_uops_1_bits_prs2_busy; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_prs3_busy = frontend_io_cpu_fetchpacket_bits_uops_1_bits_prs3_busy; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_ppred_busy = frontend_io_cpu_fetchpacket_bits_uops_1_bits_ppred_busy; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_stale_pdst = frontend_io_cpu_fetchpacket_bits_uops_1_bits_stale_pdst; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_exception = frontend_io_cpu_fetchpacket_bits_uops_1_bits_exception; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_exc_cause = frontend_io_cpu_fetchpacket_bits_uops_1_bits_exc_cause; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_bypassable = frontend_io_cpu_fetchpacket_bits_uops_1_bits_bypassable; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_mem_cmd = frontend_io_cpu_fetchpacket_bits_uops_1_bits_mem_cmd; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_mem_size = frontend_io_cpu_fetchpacket_bits_uops_1_bits_mem_size; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_mem_signed = frontend_io_cpu_fetchpacket_bits_uops_1_bits_mem_signed; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_is_fence = frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_fence; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_is_fencei = frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_fencei; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_is_amo = frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_amo; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_uses_ldq = frontend_io_cpu_fetchpacket_bits_uops_1_bits_uses_ldq; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_uses_stq = frontend_io_cpu_fetchpacket_bits_uops_1_bits_uses_stq; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_is_sys_pc2epc =
    frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_sys_pc2epc; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_is_unique = frontend_io_cpu_fetchpacket_bits_uops_1_bits_is_unique; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_flush_on_commit =
    frontend_io_cpu_fetchpacket_bits_uops_1_bits_flush_on_commit; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_ldst_is_rs1 = frontend_io_cpu_fetchpacket_bits_uops_1_bits_ldst_is_rs1
    ; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_ldst = frontend_io_cpu_fetchpacket_bits_uops_1_bits_ldst; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_lrs1 = frontend_io_cpu_fetchpacket_bits_uops_1_bits_lrs1; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_lrs2 = frontend_io_cpu_fetchpacket_bits_uops_1_bits_lrs2; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_lrs3 = frontend_io_cpu_fetchpacket_bits_uops_1_bits_lrs3; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_ldst_val = frontend_io_cpu_fetchpacket_bits_uops_1_bits_ldst_val; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_dst_rtype = frontend_io_cpu_fetchpacket_bits_uops_1_bits_dst_rtype; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_lrs1_rtype = frontend_io_cpu_fetchpacket_bits_uops_1_bits_lrs1_rtype; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_lrs2_rtype = frontend_io_cpu_fetchpacket_bits_uops_1_bits_lrs2_rtype; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_frs3_en = frontend_io_cpu_fetchpacket_bits_uops_1_bits_frs3_en; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_fp_val = frontend_io_cpu_fetchpacket_bits_uops_1_bits_fp_val; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_fp_single = frontend_io_cpu_fetchpacket_bits_uops_1_bits_fp_single; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_xcpt_pf_if = frontend_io_cpu_fetchpacket_bits_uops_1_bits_xcpt_pf_if; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_xcpt_ae_if = frontend_io_cpu_fetchpacket_bits_uops_1_bits_xcpt_ae_if; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_xcpt_ma_if = frontend_io_cpu_fetchpacket_bits_uops_1_bits_xcpt_ma_if; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_bp_debug_if = frontend_io_cpu_fetchpacket_bits_uops_1_bits_bp_debug_if
    ; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_bp_xcpt_if = frontend_io_cpu_fetchpacket_bits_uops_1_bits_bp_xcpt_if; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_debug_fsrc = frontend_io_cpu_fetchpacket_bits_uops_1_bits_debug_fsrc; // @[tile.scala 177:32]
  assign core_io_ifu_fetchpacket_bits_uops_1_bits_debug_tsrc = frontend_io_cpu_fetchpacket_bits_uops_1_bits_debug_tsrc; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_0_entry_cfi_idx_valid = frontend_io_cpu_get_pc_0_entry_cfi_idx_valid; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_0_entry_cfi_idx_bits = frontend_io_cpu_get_pc_0_entry_cfi_idx_bits; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_0_entry_cfi_taken = frontend_io_cpu_get_pc_0_entry_cfi_taken; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_0_entry_cfi_mispredicted = frontend_io_cpu_get_pc_0_entry_cfi_mispredicted; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_0_entry_cfi_type = frontend_io_cpu_get_pc_0_entry_cfi_type; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_0_entry_br_mask = frontend_io_cpu_get_pc_0_entry_br_mask; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_0_entry_cfi_is_call = frontend_io_cpu_get_pc_0_entry_cfi_is_call; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_0_entry_cfi_is_ret = frontend_io_cpu_get_pc_0_entry_cfi_is_ret; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_0_entry_cfi_npc_plus4 = frontend_io_cpu_get_pc_0_entry_cfi_npc_plus4; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_0_entry_ras_top = frontend_io_cpu_get_pc_0_entry_ras_top; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_0_entry_ras_idx = frontend_io_cpu_get_pc_0_entry_ras_idx; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_0_entry_start_bank = frontend_io_cpu_get_pc_0_entry_start_bank; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_0_ghist_old_history = frontend_io_cpu_get_pc_0_ghist_old_history; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_0_ghist_current_saw_branch_not_taken =
    frontend_io_cpu_get_pc_0_ghist_current_saw_branch_not_taken; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_0_ghist_new_saw_branch_not_taken = frontend_io_cpu_get_pc_0_ghist_new_saw_branch_not_taken; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_0_ghist_new_saw_branch_taken = frontend_io_cpu_get_pc_0_ghist_new_saw_branch_taken; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_0_ghist_ras_idx = frontend_io_cpu_get_pc_0_ghist_ras_idx; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_0_pc = frontend_io_cpu_get_pc_0_pc; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_0_com_pc = frontend_io_cpu_get_pc_0_com_pc; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_0_next_val = frontend_io_cpu_get_pc_0_next_val; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_0_next_pc = frontend_io_cpu_get_pc_0_next_pc; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_1_entry_cfi_idx_valid = frontend_io_cpu_get_pc_1_entry_cfi_idx_valid; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_1_entry_cfi_idx_bits = frontend_io_cpu_get_pc_1_entry_cfi_idx_bits; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_1_entry_cfi_taken = frontend_io_cpu_get_pc_1_entry_cfi_taken; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_1_entry_cfi_mispredicted = frontend_io_cpu_get_pc_1_entry_cfi_mispredicted; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_1_entry_cfi_type = frontend_io_cpu_get_pc_1_entry_cfi_type; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_1_entry_br_mask = frontend_io_cpu_get_pc_1_entry_br_mask; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_1_entry_cfi_is_call = frontend_io_cpu_get_pc_1_entry_cfi_is_call; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_1_entry_cfi_is_ret = frontend_io_cpu_get_pc_1_entry_cfi_is_ret; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_1_entry_cfi_npc_plus4 = frontend_io_cpu_get_pc_1_entry_cfi_npc_plus4; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_1_entry_ras_top = frontend_io_cpu_get_pc_1_entry_ras_top; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_1_entry_ras_idx = frontend_io_cpu_get_pc_1_entry_ras_idx; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_1_entry_start_bank = frontend_io_cpu_get_pc_1_entry_start_bank; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_1_ghist_old_history = frontend_io_cpu_get_pc_1_ghist_old_history; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_1_ghist_current_saw_branch_not_taken =
    frontend_io_cpu_get_pc_1_ghist_current_saw_branch_not_taken; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_1_ghist_new_saw_branch_not_taken = frontend_io_cpu_get_pc_1_ghist_new_saw_branch_not_taken; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_1_ghist_new_saw_branch_taken = frontend_io_cpu_get_pc_1_ghist_new_saw_branch_taken; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_1_ghist_ras_idx = frontend_io_cpu_get_pc_1_ghist_ras_idx; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_1_pc = frontend_io_cpu_get_pc_1_pc; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_1_com_pc = frontend_io_cpu_get_pc_1_com_pc; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_1_next_val = frontend_io_cpu_get_pc_1_next_val; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_1_next_pc = frontend_io_cpu_get_pc_1_next_pc; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_2_entry_cfi_idx_valid = frontend_io_cpu_get_pc_2_entry_cfi_idx_valid; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_2_entry_cfi_idx_bits = frontend_io_cpu_get_pc_2_entry_cfi_idx_bits; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_2_entry_cfi_taken = frontend_io_cpu_get_pc_2_entry_cfi_taken; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_2_entry_cfi_mispredicted = frontend_io_cpu_get_pc_2_entry_cfi_mispredicted; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_2_entry_cfi_type = frontend_io_cpu_get_pc_2_entry_cfi_type; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_2_entry_br_mask = frontend_io_cpu_get_pc_2_entry_br_mask; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_2_entry_cfi_is_call = frontend_io_cpu_get_pc_2_entry_cfi_is_call; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_2_entry_cfi_is_ret = frontend_io_cpu_get_pc_2_entry_cfi_is_ret; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_2_entry_cfi_npc_plus4 = frontend_io_cpu_get_pc_2_entry_cfi_npc_plus4; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_2_entry_ras_top = frontend_io_cpu_get_pc_2_entry_ras_top; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_2_entry_ras_idx = frontend_io_cpu_get_pc_2_entry_ras_idx; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_2_entry_start_bank = frontend_io_cpu_get_pc_2_entry_start_bank; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_2_ghist_old_history = frontend_io_cpu_get_pc_2_ghist_old_history; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_2_ghist_current_saw_branch_not_taken =
    frontend_io_cpu_get_pc_2_ghist_current_saw_branch_not_taken; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_2_ghist_new_saw_branch_not_taken = frontend_io_cpu_get_pc_2_ghist_new_saw_branch_not_taken; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_2_ghist_new_saw_branch_taken = frontend_io_cpu_get_pc_2_ghist_new_saw_branch_taken; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_2_ghist_ras_idx = frontend_io_cpu_get_pc_2_ghist_ras_idx; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_2_pc = frontend_io_cpu_get_pc_2_pc; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_2_com_pc = frontend_io_cpu_get_pc_2_com_pc; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_2_next_val = frontend_io_cpu_get_pc_2_next_val; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_2_next_pc = frontend_io_cpu_get_pc_2_next_pc; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_3_entry_cfi_idx_valid = frontend_io_cpu_get_pc_3_entry_cfi_idx_valid; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_3_entry_cfi_idx_bits = frontend_io_cpu_get_pc_3_entry_cfi_idx_bits; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_3_entry_cfi_taken = frontend_io_cpu_get_pc_3_entry_cfi_taken; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_3_entry_cfi_mispredicted = frontend_io_cpu_get_pc_3_entry_cfi_mispredicted; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_3_entry_cfi_type = frontend_io_cpu_get_pc_3_entry_cfi_type; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_3_entry_br_mask = frontend_io_cpu_get_pc_3_entry_br_mask; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_3_entry_cfi_is_call = frontend_io_cpu_get_pc_3_entry_cfi_is_call; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_3_entry_cfi_is_ret = frontend_io_cpu_get_pc_3_entry_cfi_is_ret; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_3_entry_cfi_npc_plus4 = frontend_io_cpu_get_pc_3_entry_cfi_npc_plus4; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_3_entry_ras_top = frontend_io_cpu_get_pc_3_entry_ras_top; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_3_entry_ras_idx = frontend_io_cpu_get_pc_3_entry_ras_idx; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_3_entry_start_bank = frontend_io_cpu_get_pc_3_entry_start_bank; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_3_ghist_old_history = frontend_io_cpu_get_pc_3_ghist_old_history; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_3_ghist_current_saw_branch_not_taken =
    frontend_io_cpu_get_pc_3_ghist_current_saw_branch_not_taken; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_3_ghist_new_saw_branch_not_taken = frontend_io_cpu_get_pc_3_ghist_new_saw_branch_not_taken; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_3_ghist_new_saw_branch_taken = frontend_io_cpu_get_pc_3_ghist_new_saw_branch_taken; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_3_ghist_ras_idx = frontend_io_cpu_get_pc_3_ghist_ras_idx; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_3_pc = frontend_io_cpu_get_pc_3_pc; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_3_com_pc = frontend_io_cpu_get_pc_3_com_pc; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_3_next_val = frontend_io_cpu_get_pc_3_next_val; // @[tile.scala 177:32]
  assign core_io_ifu_get_pc_3_next_pc = frontend_io_cpu_get_pc_3_next_pc; // @[tile.scala 177:32]
  assign core_io_ifu_debug_fetch_pc_0 = frontend_io_cpu_debug_fetch_pc_0; // @[tile.scala 177:32]
  assign core_io_ifu_debug_fetch_pc_1 = frontend_io_cpu_debug_fetch_pc_1; // @[tile.scala 177:32]
  assign core_io_ifu_perf_acquire = frontend_io_cpu_perf_acquire; // @[tile.scala 177:32]
  assign core_io_ifu_perf_tlbMiss = frontend_io_cpu_perf_tlbMiss; // @[tile.scala 177:32]
  assign core_io_ptw_perf_l2miss = ptw_io_dpath_perf_l2miss; // @[tile.scala 231:15]
  assign core_io_ptw_perf_l2hit = ptw_io_dpath_perf_l2hit; // @[tile.scala 231:15]
  assign core_io_ptw_perf_pte_miss = ptw_io_dpath_perf_pte_miss; // @[tile.scala 231:15]
  assign core_io_ptw_perf_pte_hit = ptw_io_dpath_perf_pte_hit; // @[tile.scala 231:15]
  assign core_io_ptw_clock_enabled = ptw_io_dpath_clock_enabled; // @[tile.scala 231:15]
  assign core_io_rocc_cmd_ready = 1'h0;
  assign core_io_rocc_resp_valid = 1'h0;
  assign core_io_rocc_resp_bits_rd = 5'h0;
  assign core_io_rocc_resp_bits_data = 64'h0;
  assign core_io_rocc_mem_req_valid = 1'h0;
  assign core_io_rocc_mem_req_bits_addr = 40'h0;
  assign core_io_rocc_mem_req_bits_tag = 7'h0;
  assign core_io_rocc_mem_req_bits_cmd = 5'h0;
  assign core_io_rocc_mem_req_bits_size = 2'h0;
  assign core_io_rocc_mem_req_bits_signed = 1'h0;
  assign core_io_rocc_mem_req_bits_dprv = 2'h0;
  assign core_io_rocc_mem_req_bits_phys = 1'h0;
  assign core_io_rocc_mem_req_bits_no_alloc = 1'h0;
  assign core_io_rocc_mem_req_bits_no_xcpt = 1'h0;
  assign core_io_rocc_mem_req_bits_data = 64'h0;
  assign core_io_rocc_mem_req_bits_mask = 8'h0;
  assign core_io_rocc_mem_s1_kill = 1'h0;
  assign core_io_rocc_mem_s1_data_data = 64'h0;
  assign core_io_rocc_mem_s1_data_mask = 8'h0;
  assign core_io_rocc_mem_s2_kill = 1'h0;
  assign core_io_rocc_mem_keep_clock_enabled = 1'h0;
  assign core_io_rocc_busy = 1'h0;
  assign core_io_rocc_interrupt = 1'h0;
  assign core_io_lsu_exe_0_iresp_valid = lsu_io_core_exe_0_iresp_valid; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_switch = lsu_io_core_exe_0_iresp_bits_uop_switch; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_switch_off = lsu_io_core_exe_0_iresp_bits_uop_switch_off; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_is_unicore = lsu_io_core_exe_0_iresp_bits_uop_is_unicore; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_shift = lsu_io_core_exe_0_iresp_bits_uop_shift; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_lrs3_rtype = lsu_io_core_exe_0_iresp_bits_uop_lrs3_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_rflag = lsu_io_core_exe_0_iresp_bits_uop_rflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_wflag = lsu_io_core_exe_0_iresp_bits_uop_wflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_prflag = lsu_io_core_exe_0_iresp_bits_uop_prflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_pwflag = lsu_io_core_exe_0_iresp_bits_uop_pwflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_pflag_busy = lsu_io_core_exe_0_iresp_bits_uop_pflag_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_stale_pflag = lsu_io_core_exe_0_iresp_bits_uop_stale_pflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_op1_sel = lsu_io_core_exe_0_iresp_bits_uop_op1_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_op2_sel = lsu_io_core_exe_0_iresp_bits_uop_op2_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_split_num = lsu_io_core_exe_0_iresp_bits_uop_split_num; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_self_index = lsu_io_core_exe_0_iresp_bits_uop_self_index; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_rob_inst_idx = lsu_io_core_exe_0_iresp_bits_uop_rob_inst_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_address_num = lsu_io_core_exe_0_iresp_bits_uop_address_num; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_uopc = lsu_io_core_exe_0_iresp_bits_uop_uopc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_inst = lsu_io_core_exe_0_iresp_bits_uop_inst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_debug_inst = lsu_io_core_exe_0_iresp_bits_uop_debug_inst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_is_rvc = lsu_io_core_exe_0_iresp_bits_uop_is_rvc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_debug_pc = lsu_io_core_exe_0_iresp_bits_uop_debug_pc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_iq_type = lsu_io_core_exe_0_iresp_bits_uop_iq_type; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_fu_code = lsu_io_core_exe_0_iresp_bits_uop_fu_code; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_ctrl_br_type = lsu_io_core_exe_0_iresp_bits_uop_ctrl_br_type; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_ctrl_op1_sel = lsu_io_core_exe_0_iresp_bits_uop_ctrl_op1_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_ctrl_op2_sel = lsu_io_core_exe_0_iresp_bits_uop_ctrl_op2_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_ctrl_imm_sel = lsu_io_core_exe_0_iresp_bits_uop_ctrl_imm_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_ctrl_op_fcn = lsu_io_core_exe_0_iresp_bits_uop_ctrl_op_fcn; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_ctrl_fcn_dw = lsu_io_core_exe_0_iresp_bits_uop_ctrl_fcn_dw; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_ctrl_csr_cmd = lsu_io_core_exe_0_iresp_bits_uop_ctrl_csr_cmd; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_ctrl_is_load = lsu_io_core_exe_0_iresp_bits_uop_ctrl_is_load; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_ctrl_is_sta = lsu_io_core_exe_0_iresp_bits_uop_ctrl_is_sta; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_ctrl_is_std = lsu_io_core_exe_0_iresp_bits_uop_ctrl_is_std; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_ctrl_op3_sel = lsu_io_core_exe_0_iresp_bits_uop_ctrl_op3_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_iw_state = lsu_io_core_exe_0_iresp_bits_uop_iw_state; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_iw_p1_poisoned = lsu_io_core_exe_0_iresp_bits_uop_iw_p1_poisoned; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_iw_p2_poisoned = lsu_io_core_exe_0_iresp_bits_uop_iw_p2_poisoned; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_is_br = lsu_io_core_exe_0_iresp_bits_uop_is_br; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_is_jalr = lsu_io_core_exe_0_iresp_bits_uop_is_jalr; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_is_jal = lsu_io_core_exe_0_iresp_bits_uop_is_jal; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_is_sfb = lsu_io_core_exe_0_iresp_bits_uop_is_sfb; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_br_mask = lsu_io_core_exe_0_iresp_bits_uop_br_mask; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_br_tag = lsu_io_core_exe_0_iresp_bits_uop_br_tag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_ftq_idx = lsu_io_core_exe_0_iresp_bits_uop_ftq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_edge_inst = lsu_io_core_exe_0_iresp_bits_uop_edge_inst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_pc_lob = lsu_io_core_exe_0_iresp_bits_uop_pc_lob; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_taken = lsu_io_core_exe_0_iresp_bits_uop_taken; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_imm_packed = lsu_io_core_exe_0_iresp_bits_uop_imm_packed; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_csr_addr = lsu_io_core_exe_0_iresp_bits_uop_csr_addr; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_rob_idx = lsu_io_core_exe_0_iresp_bits_uop_rob_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_ldq_idx = lsu_io_core_exe_0_iresp_bits_uop_ldq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_stq_idx = lsu_io_core_exe_0_iresp_bits_uop_stq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_rxq_idx = lsu_io_core_exe_0_iresp_bits_uop_rxq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_pdst = lsu_io_core_exe_0_iresp_bits_uop_pdst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_prs1 = lsu_io_core_exe_0_iresp_bits_uop_prs1; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_prs2 = lsu_io_core_exe_0_iresp_bits_uop_prs2; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_prs3 = lsu_io_core_exe_0_iresp_bits_uop_prs3; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_ppred = lsu_io_core_exe_0_iresp_bits_uop_ppred; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_prs1_busy = lsu_io_core_exe_0_iresp_bits_uop_prs1_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_prs2_busy = lsu_io_core_exe_0_iresp_bits_uop_prs2_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_prs3_busy = lsu_io_core_exe_0_iresp_bits_uop_prs3_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_ppred_busy = lsu_io_core_exe_0_iresp_bits_uop_ppred_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_stale_pdst = lsu_io_core_exe_0_iresp_bits_uop_stale_pdst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_exception = lsu_io_core_exe_0_iresp_bits_uop_exception; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_exc_cause = lsu_io_core_exe_0_iresp_bits_uop_exc_cause; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_bypassable = lsu_io_core_exe_0_iresp_bits_uop_bypassable; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_mem_cmd = lsu_io_core_exe_0_iresp_bits_uop_mem_cmd; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_mem_size = lsu_io_core_exe_0_iresp_bits_uop_mem_size; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_mem_signed = lsu_io_core_exe_0_iresp_bits_uop_mem_signed; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_is_fence = lsu_io_core_exe_0_iresp_bits_uop_is_fence; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_is_fencei = lsu_io_core_exe_0_iresp_bits_uop_is_fencei; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_is_amo = lsu_io_core_exe_0_iresp_bits_uop_is_amo; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_uses_ldq = lsu_io_core_exe_0_iresp_bits_uop_uses_ldq; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_uses_stq = lsu_io_core_exe_0_iresp_bits_uop_uses_stq; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_is_sys_pc2epc = lsu_io_core_exe_0_iresp_bits_uop_is_sys_pc2epc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_is_unique = lsu_io_core_exe_0_iresp_bits_uop_is_unique; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_flush_on_commit = lsu_io_core_exe_0_iresp_bits_uop_flush_on_commit; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_ldst_is_rs1 = lsu_io_core_exe_0_iresp_bits_uop_ldst_is_rs1; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_ldst = lsu_io_core_exe_0_iresp_bits_uop_ldst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_lrs1 = lsu_io_core_exe_0_iresp_bits_uop_lrs1; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_lrs2 = lsu_io_core_exe_0_iresp_bits_uop_lrs2; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_lrs3 = lsu_io_core_exe_0_iresp_bits_uop_lrs3; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_ldst_val = lsu_io_core_exe_0_iresp_bits_uop_ldst_val; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_dst_rtype = lsu_io_core_exe_0_iresp_bits_uop_dst_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_lrs1_rtype = lsu_io_core_exe_0_iresp_bits_uop_lrs1_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_lrs2_rtype = lsu_io_core_exe_0_iresp_bits_uop_lrs2_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_frs3_en = lsu_io_core_exe_0_iresp_bits_uop_frs3_en; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_fp_val = lsu_io_core_exe_0_iresp_bits_uop_fp_val; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_fp_single = lsu_io_core_exe_0_iresp_bits_uop_fp_single; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_xcpt_pf_if = lsu_io_core_exe_0_iresp_bits_uop_xcpt_pf_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_xcpt_ae_if = lsu_io_core_exe_0_iresp_bits_uop_xcpt_ae_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_xcpt_ma_if = lsu_io_core_exe_0_iresp_bits_uop_xcpt_ma_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_bp_debug_if = lsu_io_core_exe_0_iresp_bits_uop_bp_debug_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_bp_xcpt_if = lsu_io_core_exe_0_iresp_bits_uop_bp_xcpt_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_debug_fsrc = lsu_io_core_exe_0_iresp_bits_uop_debug_fsrc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_uop_debug_tsrc = lsu_io_core_exe_0_iresp_bits_uop_debug_tsrc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_data = lsu_io_core_exe_0_iresp_bits_data; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_predicated = lsu_io_core_exe_0_iresp_bits_predicated; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_valid = lsu_io_core_exe_0_iresp_bits_fflags_valid; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_switch = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_switch; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_switch_off =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_switch_off; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_unicore =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_unicore; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_shift = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_shift; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs3_rtype =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_lrs3_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_rflag = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_rflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_wflag = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_wflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_prflag = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_prflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_pwflag = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_pwflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_pflag_busy =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_pflag_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_stale_pflag =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_stale_pflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_op1_sel = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_op1_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_op2_sel = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_op2_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_split_num = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_split_num
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_self_index =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_self_index; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_rob_inst_idx =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_rob_inst_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_address_num =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_address_num; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_uopc = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_uopc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_inst = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_inst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_debug_inst =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_debug_inst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_rvc = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_rvc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_debug_pc = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_debug_pc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_iq_type = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_iq_type; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_fu_code = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_fu_code; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_br_type =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_br_type; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_op1_sel =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_op1_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_op2_sel =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_op2_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_imm_sel =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_imm_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_op_fcn =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_op_fcn; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_fcn_dw =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_fcn_dw; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_csr_cmd =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_csr_cmd; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_load =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_load; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_sta =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_sta; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_std =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_is_std; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ctrl_op3_sel =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ctrl_op3_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_iw_state = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_iw_state; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_iw_p1_poisoned =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_iw_p1_poisoned; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_iw_p2_poisoned =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_iw_p2_poisoned; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_br = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_br; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_jalr = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_jalr; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_jal = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_jal; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_sfb = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_sfb; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_br_mask = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_br_mask; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_br_tag = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_br_tag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ftq_idx = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ftq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_edge_inst = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_edge_inst
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_pc_lob = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_pc_lob; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_taken = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_taken; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_imm_packed =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_imm_packed; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_csr_addr = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_csr_addr; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_rob_idx = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_rob_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ldq_idx = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ldq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_stq_idx = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_stq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_rxq_idx = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_rxq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_pdst = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_pdst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs1 = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_prs1; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs2 = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_prs2; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs3 = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_prs3; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ppred = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ppred; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs1_busy = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_prs1_busy
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs2_busy = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_prs2_busy
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_prs3_busy = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_prs3_busy
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ppred_busy =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ppred_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_stale_pdst =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_stale_pdst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_exception = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_exception
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_exc_cause = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_exc_cause
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_bypassable =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_bypassable; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_mem_cmd = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_mem_cmd; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_mem_size = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_mem_size; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_mem_signed =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_mem_signed; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_fence = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_fence; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_fencei = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_fencei
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_amo = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_amo; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_uses_ldq = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_uses_ldq; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_uses_stq = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_uses_stq; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_sys_pc2epc =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_sys_pc2epc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_is_unique = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_is_unique
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_flush_on_commit =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_flush_on_commit; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ldst_is_rs1 =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ldst_is_rs1; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ldst = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ldst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs1 = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_lrs1; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs2 = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_lrs2; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs3 = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_lrs3; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_ldst_val = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_ldst_val; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_dst_rtype = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_dst_rtype
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs1_rtype =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_lrs1_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_lrs2_rtype =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_lrs2_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_frs3_en = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_frs3_en; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_fp_val = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_fp_val; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_fp_single = lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_fp_single
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_xcpt_pf_if =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_xcpt_pf_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_xcpt_ae_if =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_xcpt_ae_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_xcpt_ma_if =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_xcpt_ma_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_bp_debug_if =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_bp_debug_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_bp_xcpt_if =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_bp_xcpt_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_debug_fsrc =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_debug_fsrc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_uop_debug_tsrc =
    lsu_io_core_exe_0_iresp_bits_fflags_bits_uop_debug_tsrc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflags_bits_flags = lsu_io_core_exe_0_iresp_bits_fflags_bits_flags; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_flagdata = lsu_io_core_exe_0_iresp_bits_flagdata; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_valid = lsu_io_core_exe_0_iresp_bits_fflagdata_valid; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_switch = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_switch
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_switch_off =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_switch_off; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_unicore =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_unicore; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_shift = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_shift; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs3_rtype =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs3_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_rflag = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_rflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_wflag = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_wflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prflag = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_prflag
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_pwflag = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_pwflag
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_pflag_busy =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_pflag_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_stale_pflag =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_stale_pflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_op1_sel =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_op1_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_op2_sel =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_op2_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_split_num =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_split_num; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_self_index =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_self_index; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_rob_inst_idx =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_rob_inst_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_address_num =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_address_num; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_uopc = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_uopc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_inst = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_inst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_debug_inst =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_debug_inst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_rvc = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_rvc
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_debug_pc =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_debug_pc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_iq_type =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_iq_type; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_fu_code =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_fu_code; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_br_type =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_br_type; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op1_sel =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op1_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op2_sel =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op2_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_imm_sel =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_imm_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op_fcn =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op_fcn; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_fcn_dw =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_fcn_dw; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_csr_cmd =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_csr_cmd; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_load =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_load; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_sta =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_sta; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_std =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_is_std; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op3_sel =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ctrl_op3_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_iw_state =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_iw_state; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_iw_p1_poisoned =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_iw_p1_poisoned; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_iw_p2_poisoned =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_iw_p2_poisoned; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_br = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_br; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_jalr =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_jalr; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_jal = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_jal
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_sfb = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_sfb
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_br_mask =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_br_mask; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_br_tag = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_br_tag
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ftq_idx =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ftq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_edge_inst =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_edge_inst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_pc_lob = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_pc_lob
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_taken = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_taken; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_imm_packed =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_imm_packed; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_csr_addr =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_csr_addr; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_rob_idx =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_rob_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ldq_idx =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ldq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_stq_idx =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_stq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_rxq_idx =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_rxq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_pdst = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_pdst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs1 = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs1; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs2 = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs2; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs3 = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs3; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ppred = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ppred; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs1_busy =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs1_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs2_busy =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs2_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_prs3_busy =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_prs3_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ppred_busy =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ppred_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_stale_pdst =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_stale_pdst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_exception =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_exception; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_exc_cause =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_exc_cause; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_bypassable =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_bypassable; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_mem_cmd =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_mem_cmd; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_mem_size =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_mem_size; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_mem_signed =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_mem_signed; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_fence =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_fence; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_fencei =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_fencei; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_amo = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_amo
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_uses_ldq =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_uses_ldq; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_uses_stq =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_uses_stq; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_sys_pc2epc =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_sys_pc2epc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_is_unique =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_is_unique; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_flush_on_commit =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_flush_on_commit; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ldst_is_rs1 =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ldst_is_rs1; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ldst = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ldst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs1 = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs1; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs2 = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs2; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs3 = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs3; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_ldst_val =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_ldst_val; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_dst_rtype =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_dst_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs1_rtype =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs1_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_lrs2_rtype =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_lrs2_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_frs3_en =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_frs3_en; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_fp_val = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_fp_val
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_fp_single =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_fp_single; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_pf_if =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_pf_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_ae_if =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_ae_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_ma_if =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_xcpt_ma_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_bp_debug_if =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_bp_debug_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_bp_xcpt_if =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_bp_xcpt_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_debug_fsrc =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_debug_fsrc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_uop_debug_tsrc =
    lsu_io_core_exe_0_iresp_bits_fflagdata_bits_uop_debug_tsrc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_iresp_bits_fflagdata_bits_fflag = lsu_io_core_exe_0_iresp_bits_fflagdata_bits_fflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_valid = lsu_io_core_exe_0_fresp_valid; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_switch = lsu_io_core_exe_0_fresp_bits_uop_switch; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_switch_off = lsu_io_core_exe_0_fresp_bits_uop_switch_off; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_is_unicore = lsu_io_core_exe_0_fresp_bits_uop_is_unicore; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_shift = lsu_io_core_exe_0_fresp_bits_uop_shift; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_lrs3_rtype = lsu_io_core_exe_0_fresp_bits_uop_lrs3_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_rflag = lsu_io_core_exe_0_fresp_bits_uop_rflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_wflag = lsu_io_core_exe_0_fresp_bits_uop_wflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_prflag = lsu_io_core_exe_0_fresp_bits_uop_prflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_pwflag = lsu_io_core_exe_0_fresp_bits_uop_pwflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_pflag_busy = lsu_io_core_exe_0_fresp_bits_uop_pflag_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_stale_pflag = lsu_io_core_exe_0_fresp_bits_uop_stale_pflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_op1_sel = lsu_io_core_exe_0_fresp_bits_uop_op1_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_op2_sel = lsu_io_core_exe_0_fresp_bits_uop_op2_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_split_num = lsu_io_core_exe_0_fresp_bits_uop_split_num; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_self_index = lsu_io_core_exe_0_fresp_bits_uop_self_index; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_rob_inst_idx = lsu_io_core_exe_0_fresp_bits_uop_rob_inst_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_address_num = lsu_io_core_exe_0_fresp_bits_uop_address_num; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_uopc = lsu_io_core_exe_0_fresp_bits_uop_uopc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_inst = lsu_io_core_exe_0_fresp_bits_uop_inst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_debug_inst = lsu_io_core_exe_0_fresp_bits_uop_debug_inst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_is_rvc = lsu_io_core_exe_0_fresp_bits_uop_is_rvc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_debug_pc = lsu_io_core_exe_0_fresp_bits_uop_debug_pc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_iq_type = lsu_io_core_exe_0_fresp_bits_uop_iq_type; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_fu_code = lsu_io_core_exe_0_fresp_bits_uop_fu_code; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_ctrl_br_type = lsu_io_core_exe_0_fresp_bits_uop_ctrl_br_type; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_ctrl_op1_sel = lsu_io_core_exe_0_fresp_bits_uop_ctrl_op1_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_ctrl_op2_sel = lsu_io_core_exe_0_fresp_bits_uop_ctrl_op2_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_ctrl_imm_sel = lsu_io_core_exe_0_fresp_bits_uop_ctrl_imm_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_ctrl_op_fcn = lsu_io_core_exe_0_fresp_bits_uop_ctrl_op_fcn; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_ctrl_fcn_dw = lsu_io_core_exe_0_fresp_bits_uop_ctrl_fcn_dw; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_ctrl_csr_cmd = lsu_io_core_exe_0_fresp_bits_uop_ctrl_csr_cmd; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_ctrl_is_load = lsu_io_core_exe_0_fresp_bits_uop_ctrl_is_load; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_ctrl_is_sta = lsu_io_core_exe_0_fresp_bits_uop_ctrl_is_sta; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_ctrl_is_std = lsu_io_core_exe_0_fresp_bits_uop_ctrl_is_std; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_ctrl_op3_sel = lsu_io_core_exe_0_fresp_bits_uop_ctrl_op3_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_iw_state = lsu_io_core_exe_0_fresp_bits_uop_iw_state; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_iw_p1_poisoned = lsu_io_core_exe_0_fresp_bits_uop_iw_p1_poisoned; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_iw_p2_poisoned = lsu_io_core_exe_0_fresp_bits_uop_iw_p2_poisoned; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_is_br = lsu_io_core_exe_0_fresp_bits_uop_is_br; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_is_jalr = lsu_io_core_exe_0_fresp_bits_uop_is_jalr; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_is_jal = lsu_io_core_exe_0_fresp_bits_uop_is_jal; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_is_sfb = lsu_io_core_exe_0_fresp_bits_uop_is_sfb; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_br_mask = lsu_io_core_exe_0_fresp_bits_uop_br_mask; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_br_tag = lsu_io_core_exe_0_fresp_bits_uop_br_tag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_ftq_idx = lsu_io_core_exe_0_fresp_bits_uop_ftq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_edge_inst = lsu_io_core_exe_0_fresp_bits_uop_edge_inst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_pc_lob = lsu_io_core_exe_0_fresp_bits_uop_pc_lob; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_taken = lsu_io_core_exe_0_fresp_bits_uop_taken; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_imm_packed = lsu_io_core_exe_0_fresp_bits_uop_imm_packed; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_csr_addr = lsu_io_core_exe_0_fresp_bits_uop_csr_addr; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_rob_idx = lsu_io_core_exe_0_fresp_bits_uop_rob_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_ldq_idx = lsu_io_core_exe_0_fresp_bits_uop_ldq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_stq_idx = lsu_io_core_exe_0_fresp_bits_uop_stq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_rxq_idx = lsu_io_core_exe_0_fresp_bits_uop_rxq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_pdst = lsu_io_core_exe_0_fresp_bits_uop_pdst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_prs1 = lsu_io_core_exe_0_fresp_bits_uop_prs1; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_prs2 = lsu_io_core_exe_0_fresp_bits_uop_prs2; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_prs3 = lsu_io_core_exe_0_fresp_bits_uop_prs3; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_ppred = lsu_io_core_exe_0_fresp_bits_uop_ppred; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_prs1_busy = lsu_io_core_exe_0_fresp_bits_uop_prs1_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_prs2_busy = lsu_io_core_exe_0_fresp_bits_uop_prs2_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_prs3_busy = lsu_io_core_exe_0_fresp_bits_uop_prs3_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_ppred_busy = lsu_io_core_exe_0_fresp_bits_uop_ppred_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_stale_pdst = lsu_io_core_exe_0_fresp_bits_uop_stale_pdst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_exception = lsu_io_core_exe_0_fresp_bits_uop_exception; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_exc_cause = lsu_io_core_exe_0_fresp_bits_uop_exc_cause; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_bypassable = lsu_io_core_exe_0_fresp_bits_uop_bypassable; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_mem_cmd = lsu_io_core_exe_0_fresp_bits_uop_mem_cmd; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_mem_size = lsu_io_core_exe_0_fresp_bits_uop_mem_size; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_mem_signed = lsu_io_core_exe_0_fresp_bits_uop_mem_signed; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_is_fence = lsu_io_core_exe_0_fresp_bits_uop_is_fence; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_is_fencei = lsu_io_core_exe_0_fresp_bits_uop_is_fencei; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_is_amo = lsu_io_core_exe_0_fresp_bits_uop_is_amo; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_uses_ldq = lsu_io_core_exe_0_fresp_bits_uop_uses_ldq; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_uses_stq = lsu_io_core_exe_0_fresp_bits_uop_uses_stq; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_is_sys_pc2epc = lsu_io_core_exe_0_fresp_bits_uop_is_sys_pc2epc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_is_unique = lsu_io_core_exe_0_fresp_bits_uop_is_unique; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_flush_on_commit = lsu_io_core_exe_0_fresp_bits_uop_flush_on_commit; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_ldst_is_rs1 = lsu_io_core_exe_0_fresp_bits_uop_ldst_is_rs1; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_ldst = lsu_io_core_exe_0_fresp_bits_uop_ldst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_lrs1 = lsu_io_core_exe_0_fresp_bits_uop_lrs1; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_lrs2 = lsu_io_core_exe_0_fresp_bits_uop_lrs2; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_lrs3 = lsu_io_core_exe_0_fresp_bits_uop_lrs3; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_ldst_val = lsu_io_core_exe_0_fresp_bits_uop_ldst_val; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_dst_rtype = lsu_io_core_exe_0_fresp_bits_uop_dst_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_lrs1_rtype = lsu_io_core_exe_0_fresp_bits_uop_lrs1_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_lrs2_rtype = lsu_io_core_exe_0_fresp_bits_uop_lrs2_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_frs3_en = lsu_io_core_exe_0_fresp_bits_uop_frs3_en; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_fp_val = lsu_io_core_exe_0_fresp_bits_uop_fp_val; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_fp_single = lsu_io_core_exe_0_fresp_bits_uop_fp_single; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_xcpt_pf_if = lsu_io_core_exe_0_fresp_bits_uop_xcpt_pf_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_xcpt_ae_if = lsu_io_core_exe_0_fresp_bits_uop_xcpt_ae_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_xcpt_ma_if = lsu_io_core_exe_0_fresp_bits_uop_xcpt_ma_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_bp_debug_if = lsu_io_core_exe_0_fresp_bits_uop_bp_debug_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_bp_xcpt_if = lsu_io_core_exe_0_fresp_bits_uop_bp_xcpt_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_debug_fsrc = lsu_io_core_exe_0_fresp_bits_uop_debug_fsrc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_uop_debug_tsrc = lsu_io_core_exe_0_fresp_bits_uop_debug_tsrc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_data = lsu_io_core_exe_0_fresp_bits_data; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_predicated = lsu_io_core_exe_0_fresp_bits_predicated; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_valid = lsu_io_core_exe_0_fresp_bits_fflags_valid; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_switch = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_switch; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_switch_off =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_switch_off; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_unicore =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_unicore; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_shift = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_shift; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs3_rtype =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_lrs3_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_rflag = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_rflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_wflag = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_wflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_prflag = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_prflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_pwflag = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_pwflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_pflag_busy =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_pflag_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_stale_pflag =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_stale_pflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_op1_sel = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_op1_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_op2_sel = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_op2_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_split_num = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_split_num
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_self_index =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_self_index; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_rob_inst_idx =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_rob_inst_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_address_num =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_address_num; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_uopc = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_uopc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_inst = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_inst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_debug_inst =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_debug_inst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_rvc = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_rvc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_debug_pc = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_debug_pc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_iq_type = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_iq_type; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_fu_code = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_fu_code; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_br_type =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_br_type; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_op1_sel =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_op1_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_op2_sel =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_op2_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_imm_sel =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_imm_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_op_fcn =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_op_fcn; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_fcn_dw =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_fcn_dw; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_csr_cmd =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_csr_cmd; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_load =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_load; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_sta =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_sta; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_std =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_is_std; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ctrl_op3_sel =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ctrl_op3_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_iw_state = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_iw_state; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_iw_p1_poisoned =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_iw_p1_poisoned; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_iw_p2_poisoned =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_iw_p2_poisoned; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_br = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_br; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_jalr = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_jalr; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_jal = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_jal; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_sfb = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_sfb; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_br_mask = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_br_mask; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_br_tag = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_br_tag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ftq_idx = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ftq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_edge_inst = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_edge_inst
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_pc_lob = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_pc_lob; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_taken = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_taken; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_imm_packed =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_imm_packed; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_csr_addr = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_csr_addr; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_rob_idx = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_rob_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ldq_idx = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ldq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_stq_idx = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_stq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_rxq_idx = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_rxq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_pdst = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_pdst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs1 = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_prs1; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs2 = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_prs2; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs3 = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_prs3; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ppred = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ppred; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs1_busy = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_prs1_busy
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs2_busy = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_prs2_busy
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_prs3_busy = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_prs3_busy
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ppred_busy =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ppred_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_stale_pdst =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_stale_pdst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_exception = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_exception
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_exc_cause = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_exc_cause
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_bypassable =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_bypassable; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_mem_cmd = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_mem_cmd; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_mem_size = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_mem_size; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_mem_signed =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_mem_signed; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_fence = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_fence; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_fencei = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_fencei
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_amo = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_amo; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_uses_ldq = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_uses_ldq; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_uses_stq = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_uses_stq; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_sys_pc2epc =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_sys_pc2epc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_is_unique = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_is_unique
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_flush_on_commit =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_flush_on_commit; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ldst_is_rs1 =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ldst_is_rs1; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ldst = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ldst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs1 = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_lrs1; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs2 = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_lrs2; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs3 = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_lrs3; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_ldst_val = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_ldst_val; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_dst_rtype = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_dst_rtype
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs1_rtype =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_lrs1_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_lrs2_rtype =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_lrs2_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_frs3_en = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_frs3_en; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_fp_val = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_fp_val; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_fp_single = lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_fp_single
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_xcpt_pf_if =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_xcpt_pf_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_xcpt_ae_if =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_xcpt_ae_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_xcpt_ma_if =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_xcpt_ma_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_bp_debug_if =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_bp_debug_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_bp_xcpt_if =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_bp_xcpt_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_debug_fsrc =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_debug_fsrc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_uop_debug_tsrc =
    lsu_io_core_exe_0_fresp_bits_fflags_bits_uop_debug_tsrc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflags_bits_flags = lsu_io_core_exe_0_fresp_bits_fflags_bits_flags; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_flagdata = lsu_io_core_exe_0_fresp_bits_flagdata; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_valid = lsu_io_core_exe_0_fresp_bits_fflagdata_valid; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_switch = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_switch
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_switch_off =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_switch_off; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_unicore =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_unicore; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_shift = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_shift; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs3_rtype =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs3_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_rflag = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_rflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_wflag = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_wflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prflag = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_prflag
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_pwflag = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_pwflag
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_pflag_busy =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_pflag_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_stale_pflag =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_stale_pflag; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_op1_sel =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_op1_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_op2_sel =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_op2_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_split_num =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_split_num; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_self_index =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_self_index; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_rob_inst_idx =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_rob_inst_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_address_num =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_address_num; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_uopc = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_uopc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_inst = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_inst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_debug_inst =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_debug_inst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_rvc = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_rvc
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_debug_pc =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_debug_pc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_iq_type =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_iq_type; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_fu_code =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_fu_code; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_br_type =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_br_type; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op1_sel =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op1_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op2_sel =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op2_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_imm_sel =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_imm_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op_fcn =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op_fcn; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_fcn_dw =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_fcn_dw; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_csr_cmd =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_csr_cmd; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_load =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_load; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_sta =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_sta; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_std =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_is_std; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op3_sel =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ctrl_op3_sel; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_iw_state =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_iw_state; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_iw_p1_poisoned =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_iw_p1_poisoned; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_iw_p2_poisoned =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_iw_p2_poisoned; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_br = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_br; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_jalr =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_jalr; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_jal = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_jal
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_sfb = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_sfb
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_br_mask =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_br_mask; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_br_tag = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_br_tag
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ftq_idx =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ftq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_edge_inst =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_edge_inst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_pc_lob = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_pc_lob
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_taken = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_taken; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_imm_packed =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_imm_packed; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_csr_addr =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_csr_addr; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_rob_idx =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_rob_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ldq_idx =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ldq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_stq_idx =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_stq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_rxq_idx =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_rxq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_pdst = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_pdst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs1 = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs1; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs2 = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs2; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs3 = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs3; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ppred = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ppred; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs1_busy =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs1_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs2_busy =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs2_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_prs3_busy =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_prs3_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ppred_busy =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ppred_busy; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_stale_pdst =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_stale_pdst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_exception =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_exception; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_exc_cause =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_exc_cause; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_bypassable =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_bypassable; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_mem_cmd =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_mem_cmd; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_mem_size =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_mem_size; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_mem_signed =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_mem_signed; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_fence =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_fence; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_fencei =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_fencei; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_amo = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_amo
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_uses_ldq =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_uses_ldq; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_uses_stq =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_uses_stq; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_sys_pc2epc =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_sys_pc2epc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_is_unique =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_is_unique; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_flush_on_commit =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_flush_on_commit; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ldst_is_rs1 =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ldst_is_rs1; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ldst = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ldst; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs1 = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs1; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs2 = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs2; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs3 = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs3; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_ldst_val =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_ldst_val; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_dst_rtype =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_dst_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs1_rtype =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs1_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_lrs2_rtype =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_lrs2_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_frs3_en =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_frs3_en; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_fp_val = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_fp_val
    ; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_fp_single =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_fp_single; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_pf_if =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_pf_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_ae_if =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_ae_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_ma_if =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_xcpt_ma_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_bp_debug_if =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_bp_debug_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_bp_xcpt_if =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_bp_xcpt_if; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_debug_fsrc =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_debug_fsrc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_uop_debug_tsrc =
    lsu_io_core_exe_0_fresp_bits_fflagdata_bits_uop_debug_tsrc; // @[tile.scala 178:15]
  assign core_io_lsu_exe_0_fresp_bits_fflagdata_bits_fflag = lsu_io_core_exe_0_fresp_bits_fflagdata_bits_fflag; // @[tile.scala 178:15]
  assign core_io_lsu_dis_ldq_idx_0 = lsu_io_core_dis_ldq_idx_0; // @[tile.scala 178:15]
  assign core_io_lsu_dis_ldq_idx_1 = lsu_io_core_dis_ldq_idx_1; // @[tile.scala 178:15]
  assign core_io_lsu_dis_stq_idx_0 = lsu_io_core_dis_stq_idx_0; // @[tile.scala 178:15]
  assign core_io_lsu_dis_stq_idx_1 = lsu_io_core_dis_stq_idx_1; // @[tile.scala 178:15]
  assign core_io_lsu_ldq_full_0 = lsu_io_core_ldq_full_0; // @[tile.scala 178:15]
  assign core_io_lsu_ldq_full_1 = lsu_io_core_ldq_full_1; // @[tile.scala 178:15]
  assign core_io_lsu_stq_full_0 = lsu_io_core_stq_full_0; // @[tile.scala 178:15]
  assign core_io_lsu_stq_full_1 = lsu_io_core_stq_full_1; // @[tile.scala 178:15]
  assign core_io_lsu_fp_stdata_ready = lsu_io_core_fp_stdata_ready; // @[tile.scala 178:15]
  assign core_io_lsu_clr_bsy_0_valid = lsu_io_core_clr_bsy_0_valid; // @[tile.scala 178:15]
  assign core_io_lsu_clr_bsy_0_bits = lsu_io_core_clr_bsy_0_bits; // @[tile.scala 178:15]
  assign core_io_lsu_clr_bsy_1_valid = lsu_io_core_clr_bsy_1_valid; // @[tile.scala 178:15]
  assign core_io_lsu_clr_bsy_1_bits = lsu_io_core_clr_bsy_1_bits; // @[tile.scala 178:15]
  assign core_io_lsu_clr_unsafe_0_valid = lsu_io_core_clr_unsafe_0_valid; // @[tile.scala 178:15]
  assign core_io_lsu_clr_unsafe_0_bits = lsu_io_core_clr_unsafe_0_bits; // @[tile.scala 178:15]
  assign core_io_lsu_clr_bsy_first_idx_0 = lsu_io_core_clr_bsy_first_idx_0; // @[tile.scala 178:15]
  assign core_io_lsu_clr_bsy_first_idx_1 = lsu_io_core_clr_bsy_first_idx_1; // @[tile.scala 178:15]
  assign core_io_lsu_clr_bsy_self_idx_0 = lsu_io_core_clr_bsy_self_idx_0; // @[tile.scala 178:15]
  assign core_io_lsu_clr_bsy_self_idx_1 = lsu_io_core_clr_bsy_self_idx_1; // @[tile.scala 178:15]
  assign core_io_lsu_spec_ld_wakeup_0_valid = lsu_io_core_spec_ld_wakeup_0_valid; // @[tile.scala 178:15]
  assign core_io_lsu_spec_ld_wakeup_0_bits = lsu_io_core_spec_ld_wakeup_0_bits; // @[tile.scala 178:15]
  assign core_io_lsu_ld_miss = lsu_io_core_ld_miss; // @[tile.scala 178:15]
  assign core_io_lsu_fencei_rdy = lsu_io_core_fencei_rdy; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_valid = lsu_io_core_lxcpt_valid; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_switch = lsu_io_core_lxcpt_bits_uop_switch; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_switch_off = lsu_io_core_lxcpt_bits_uop_switch_off; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_is_unicore = lsu_io_core_lxcpt_bits_uop_is_unicore; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_shift = lsu_io_core_lxcpt_bits_uop_shift; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_lrs3_rtype = lsu_io_core_lxcpt_bits_uop_lrs3_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_rflag = lsu_io_core_lxcpt_bits_uop_rflag; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_wflag = lsu_io_core_lxcpt_bits_uop_wflag; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_prflag = lsu_io_core_lxcpt_bits_uop_prflag; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_pwflag = lsu_io_core_lxcpt_bits_uop_pwflag; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_pflag_busy = lsu_io_core_lxcpt_bits_uop_pflag_busy; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_stale_pflag = lsu_io_core_lxcpt_bits_uop_stale_pflag; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_op1_sel = lsu_io_core_lxcpt_bits_uop_op1_sel; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_op2_sel = lsu_io_core_lxcpt_bits_uop_op2_sel; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_split_num = lsu_io_core_lxcpt_bits_uop_split_num; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_self_index = lsu_io_core_lxcpt_bits_uop_self_index; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_rob_inst_idx = lsu_io_core_lxcpt_bits_uop_rob_inst_idx; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_address_num = lsu_io_core_lxcpt_bits_uop_address_num; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_uopc = lsu_io_core_lxcpt_bits_uop_uopc; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_inst = lsu_io_core_lxcpt_bits_uop_inst; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_debug_inst = lsu_io_core_lxcpt_bits_uop_debug_inst; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_is_rvc = lsu_io_core_lxcpt_bits_uop_is_rvc; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_debug_pc = lsu_io_core_lxcpt_bits_uop_debug_pc; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_iq_type = lsu_io_core_lxcpt_bits_uop_iq_type; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_fu_code = lsu_io_core_lxcpt_bits_uop_fu_code; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_ctrl_br_type = lsu_io_core_lxcpt_bits_uop_ctrl_br_type; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_ctrl_op1_sel = lsu_io_core_lxcpt_bits_uop_ctrl_op1_sel; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_ctrl_op2_sel = lsu_io_core_lxcpt_bits_uop_ctrl_op2_sel; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_ctrl_imm_sel = lsu_io_core_lxcpt_bits_uop_ctrl_imm_sel; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_ctrl_op_fcn = lsu_io_core_lxcpt_bits_uop_ctrl_op_fcn; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_ctrl_fcn_dw = lsu_io_core_lxcpt_bits_uop_ctrl_fcn_dw; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_ctrl_csr_cmd = lsu_io_core_lxcpt_bits_uop_ctrl_csr_cmd; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_ctrl_is_load = lsu_io_core_lxcpt_bits_uop_ctrl_is_load; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_ctrl_is_sta = lsu_io_core_lxcpt_bits_uop_ctrl_is_sta; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_ctrl_is_std = lsu_io_core_lxcpt_bits_uop_ctrl_is_std; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_ctrl_op3_sel = lsu_io_core_lxcpt_bits_uop_ctrl_op3_sel; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_iw_state = lsu_io_core_lxcpt_bits_uop_iw_state; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_iw_p1_poisoned = lsu_io_core_lxcpt_bits_uop_iw_p1_poisoned; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_iw_p2_poisoned = lsu_io_core_lxcpt_bits_uop_iw_p2_poisoned; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_is_br = lsu_io_core_lxcpt_bits_uop_is_br; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_is_jalr = lsu_io_core_lxcpt_bits_uop_is_jalr; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_is_jal = lsu_io_core_lxcpt_bits_uop_is_jal; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_is_sfb = lsu_io_core_lxcpt_bits_uop_is_sfb; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_br_mask = lsu_io_core_lxcpt_bits_uop_br_mask; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_br_tag = lsu_io_core_lxcpt_bits_uop_br_tag; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_ftq_idx = lsu_io_core_lxcpt_bits_uop_ftq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_edge_inst = lsu_io_core_lxcpt_bits_uop_edge_inst; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_pc_lob = lsu_io_core_lxcpt_bits_uop_pc_lob; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_taken = lsu_io_core_lxcpt_bits_uop_taken; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_imm_packed = lsu_io_core_lxcpt_bits_uop_imm_packed; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_csr_addr = lsu_io_core_lxcpt_bits_uop_csr_addr; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_rob_idx = lsu_io_core_lxcpt_bits_uop_rob_idx; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_ldq_idx = lsu_io_core_lxcpt_bits_uop_ldq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_stq_idx = lsu_io_core_lxcpt_bits_uop_stq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_rxq_idx = lsu_io_core_lxcpt_bits_uop_rxq_idx; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_pdst = lsu_io_core_lxcpt_bits_uop_pdst; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_prs1 = lsu_io_core_lxcpt_bits_uop_prs1; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_prs2 = lsu_io_core_lxcpt_bits_uop_prs2; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_prs3 = lsu_io_core_lxcpt_bits_uop_prs3; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_ppred = lsu_io_core_lxcpt_bits_uop_ppred; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_prs1_busy = lsu_io_core_lxcpt_bits_uop_prs1_busy; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_prs2_busy = lsu_io_core_lxcpt_bits_uop_prs2_busy; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_prs3_busy = lsu_io_core_lxcpt_bits_uop_prs3_busy; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_ppred_busy = lsu_io_core_lxcpt_bits_uop_ppred_busy; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_stale_pdst = lsu_io_core_lxcpt_bits_uop_stale_pdst; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_exception = lsu_io_core_lxcpt_bits_uop_exception; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_exc_cause = lsu_io_core_lxcpt_bits_uop_exc_cause; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_bypassable = lsu_io_core_lxcpt_bits_uop_bypassable; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_mem_cmd = lsu_io_core_lxcpt_bits_uop_mem_cmd; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_mem_size = lsu_io_core_lxcpt_bits_uop_mem_size; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_mem_signed = lsu_io_core_lxcpt_bits_uop_mem_signed; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_is_fence = lsu_io_core_lxcpt_bits_uop_is_fence; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_is_fencei = lsu_io_core_lxcpt_bits_uop_is_fencei; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_is_amo = lsu_io_core_lxcpt_bits_uop_is_amo; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_uses_ldq = lsu_io_core_lxcpt_bits_uop_uses_ldq; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_uses_stq = lsu_io_core_lxcpt_bits_uop_uses_stq; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_is_sys_pc2epc = lsu_io_core_lxcpt_bits_uop_is_sys_pc2epc; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_is_unique = lsu_io_core_lxcpt_bits_uop_is_unique; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_flush_on_commit = lsu_io_core_lxcpt_bits_uop_flush_on_commit; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_ldst_is_rs1 = lsu_io_core_lxcpt_bits_uop_ldst_is_rs1; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_ldst = lsu_io_core_lxcpt_bits_uop_ldst; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_lrs1 = lsu_io_core_lxcpt_bits_uop_lrs1; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_lrs2 = lsu_io_core_lxcpt_bits_uop_lrs2; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_lrs3 = lsu_io_core_lxcpt_bits_uop_lrs3; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_ldst_val = lsu_io_core_lxcpt_bits_uop_ldst_val; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_dst_rtype = lsu_io_core_lxcpt_bits_uop_dst_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_lrs1_rtype = lsu_io_core_lxcpt_bits_uop_lrs1_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_lrs2_rtype = lsu_io_core_lxcpt_bits_uop_lrs2_rtype; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_frs3_en = lsu_io_core_lxcpt_bits_uop_frs3_en; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_fp_val = lsu_io_core_lxcpt_bits_uop_fp_val; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_fp_single = lsu_io_core_lxcpt_bits_uop_fp_single; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_xcpt_pf_if = lsu_io_core_lxcpt_bits_uop_xcpt_pf_if; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_xcpt_ae_if = lsu_io_core_lxcpt_bits_uop_xcpt_ae_if; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_xcpt_ma_if = lsu_io_core_lxcpt_bits_uop_xcpt_ma_if; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_bp_debug_if = lsu_io_core_lxcpt_bits_uop_bp_debug_if; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_bp_xcpt_if = lsu_io_core_lxcpt_bits_uop_bp_xcpt_if; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_debug_fsrc = lsu_io_core_lxcpt_bits_uop_debug_fsrc; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_uop_debug_tsrc = lsu_io_core_lxcpt_bits_uop_debug_tsrc; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_cause = lsu_io_core_lxcpt_bits_cause; // @[tile.scala 178:15]
  assign core_io_lsu_lxcpt_bits_badvaddr = lsu_io_core_lxcpt_bits_badvaddr; // @[tile.scala 178:15]
  assign core_io_lsu_perf_acquire = lsu_io_core_perf_acquire; // @[tile.scala 178:15]
  assign core_io_lsu_perf_release = lsu_io_core_perf_release; // @[tile.scala 178:15]
  assign core_io_lsu_perf_tlbMiss = lsu_io_core_perf_tlbMiss; // @[tile.scala 178:15]
  assign core_io_ptw_tlb_req_ready = ptw_io_requestor_2_req_ready; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_resp_valid = ptw_io_requestor_2_resp_valid; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_resp_bits_ae = ptw_io_requestor_2_resp_bits_ae; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_resp_bits_pte_ppn = ptw_io_requestor_2_resp_bits_pte_ppn; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_resp_bits_pte_reserved_for_software = ptw_io_requestor_2_resp_bits_pte_reserved_for_software; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_resp_bits_pte_d = ptw_io_requestor_2_resp_bits_pte_d; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_resp_bits_pte_a = ptw_io_requestor_2_resp_bits_pte_a; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_resp_bits_pte_g = ptw_io_requestor_2_resp_bits_pte_g; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_resp_bits_pte_u = ptw_io_requestor_2_resp_bits_pte_u; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_resp_bits_pte_x = ptw_io_requestor_2_resp_bits_pte_x; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_resp_bits_pte_w = ptw_io_requestor_2_resp_bits_pte_w; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_resp_bits_pte_r = ptw_io_requestor_2_resp_bits_pte_r; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_resp_bits_pte_v = ptw_io_requestor_2_resp_bits_pte_v; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_resp_bits_level = ptw_io_requestor_2_resp_bits_level; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_resp_bits_fragmented_superpage = ptw_io_requestor_2_resp_bits_fragmented_superpage; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_resp_bits_homogeneous = ptw_io_requestor_2_resp_bits_homogeneous; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_ptbr_mode = ptw_io_requestor_2_ptbr_mode; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_ptbr_asid = ptw_io_requestor_2_ptbr_asid; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_ptbr_ppn = ptw_io_requestor_2_ptbr_ppn; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_debug = ptw_io_requestor_2_status_debug; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_cease = ptw_io_requestor_2_status_cease; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_wfi = ptw_io_requestor_2_status_wfi; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_isa = ptw_io_requestor_2_status_isa; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_dprv = ptw_io_requestor_2_status_dprv; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_prv = ptw_io_requestor_2_status_prv; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_sd = ptw_io_requestor_2_status_sd; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_zero2 = ptw_io_requestor_2_status_zero2; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_sxl = ptw_io_requestor_2_status_sxl; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_uxl = ptw_io_requestor_2_status_uxl; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_sd_rv32 = ptw_io_requestor_2_status_sd_rv32; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_zero1 = ptw_io_requestor_2_status_zero1; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_tsr = ptw_io_requestor_2_status_tsr; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_tw = ptw_io_requestor_2_status_tw; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_tvm = ptw_io_requestor_2_status_tvm; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_mxr = ptw_io_requestor_2_status_mxr; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_sum = ptw_io_requestor_2_status_sum; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_mprv = ptw_io_requestor_2_status_mprv; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_xs = ptw_io_requestor_2_status_xs; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_fs = ptw_io_requestor_2_status_fs; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_mpp = ptw_io_requestor_2_status_mpp; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_vs = ptw_io_requestor_2_status_vs; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_spp = ptw_io_requestor_2_status_spp; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_mpie = ptw_io_requestor_2_status_mpie; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_hpie = ptw_io_requestor_2_status_hpie; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_spie = ptw_io_requestor_2_status_spie; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_upie = ptw_io_requestor_2_status_upie; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_mie = ptw_io_requestor_2_status_mie; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_hie = ptw_io_requestor_2_status_hie; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_sie = ptw_io_requestor_2_status_sie; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_status_uie = ptw_io_requestor_2_status_uie; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_0_cfg_l = ptw_io_requestor_2_pmp_0_cfg_l; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_0_cfg_res = ptw_io_requestor_2_pmp_0_cfg_res; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_0_cfg_a = ptw_io_requestor_2_pmp_0_cfg_a; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_0_cfg_x = ptw_io_requestor_2_pmp_0_cfg_x; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_0_cfg_w = ptw_io_requestor_2_pmp_0_cfg_w; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_0_cfg_r = ptw_io_requestor_2_pmp_0_cfg_r; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_0_addr = ptw_io_requestor_2_pmp_0_addr; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_0_mask = ptw_io_requestor_2_pmp_0_mask; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_1_cfg_l = ptw_io_requestor_2_pmp_1_cfg_l; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_1_cfg_res = ptw_io_requestor_2_pmp_1_cfg_res; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_1_cfg_a = ptw_io_requestor_2_pmp_1_cfg_a; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_1_cfg_x = ptw_io_requestor_2_pmp_1_cfg_x; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_1_cfg_w = ptw_io_requestor_2_pmp_1_cfg_w; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_1_cfg_r = ptw_io_requestor_2_pmp_1_cfg_r; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_1_addr = ptw_io_requestor_2_pmp_1_addr; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_1_mask = ptw_io_requestor_2_pmp_1_mask; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_2_cfg_l = ptw_io_requestor_2_pmp_2_cfg_l; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_2_cfg_res = ptw_io_requestor_2_pmp_2_cfg_res; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_2_cfg_a = ptw_io_requestor_2_pmp_2_cfg_a; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_2_cfg_x = ptw_io_requestor_2_pmp_2_cfg_x; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_2_cfg_w = ptw_io_requestor_2_pmp_2_cfg_w; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_2_cfg_r = ptw_io_requestor_2_pmp_2_cfg_r; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_2_addr = ptw_io_requestor_2_pmp_2_addr; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_2_mask = ptw_io_requestor_2_pmp_2_mask; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_3_cfg_l = ptw_io_requestor_2_pmp_3_cfg_l; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_3_cfg_res = ptw_io_requestor_2_pmp_3_cfg_res; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_3_cfg_a = ptw_io_requestor_2_pmp_3_cfg_a; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_3_cfg_x = ptw_io_requestor_2_pmp_3_cfg_x; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_3_cfg_w = ptw_io_requestor_2_pmp_3_cfg_w; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_3_cfg_r = ptw_io_requestor_2_pmp_3_cfg_r; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_3_addr = ptw_io_requestor_2_pmp_3_addr; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_3_mask = ptw_io_requestor_2_pmp_3_mask; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_4_cfg_l = ptw_io_requestor_2_pmp_4_cfg_l; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_4_cfg_res = ptw_io_requestor_2_pmp_4_cfg_res; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_4_cfg_a = ptw_io_requestor_2_pmp_4_cfg_a; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_4_cfg_x = ptw_io_requestor_2_pmp_4_cfg_x; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_4_cfg_w = ptw_io_requestor_2_pmp_4_cfg_w; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_4_cfg_r = ptw_io_requestor_2_pmp_4_cfg_r; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_4_addr = ptw_io_requestor_2_pmp_4_addr; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_4_mask = ptw_io_requestor_2_pmp_4_mask; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_5_cfg_l = ptw_io_requestor_2_pmp_5_cfg_l; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_5_cfg_res = ptw_io_requestor_2_pmp_5_cfg_res; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_5_cfg_a = ptw_io_requestor_2_pmp_5_cfg_a; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_5_cfg_x = ptw_io_requestor_2_pmp_5_cfg_x; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_5_cfg_w = ptw_io_requestor_2_pmp_5_cfg_w; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_5_cfg_r = ptw_io_requestor_2_pmp_5_cfg_r; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_5_addr = ptw_io_requestor_2_pmp_5_addr; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_5_mask = ptw_io_requestor_2_pmp_5_mask; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_6_cfg_l = ptw_io_requestor_2_pmp_6_cfg_l; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_6_cfg_res = ptw_io_requestor_2_pmp_6_cfg_res; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_6_cfg_a = ptw_io_requestor_2_pmp_6_cfg_a; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_6_cfg_x = ptw_io_requestor_2_pmp_6_cfg_x; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_6_cfg_w = ptw_io_requestor_2_pmp_6_cfg_w; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_6_cfg_r = ptw_io_requestor_2_pmp_6_cfg_r; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_6_addr = ptw_io_requestor_2_pmp_6_addr; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_6_mask = ptw_io_requestor_2_pmp_6_mask; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_7_cfg_l = ptw_io_requestor_2_pmp_7_cfg_l; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_7_cfg_res = ptw_io_requestor_2_pmp_7_cfg_res; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_7_cfg_a = ptw_io_requestor_2_pmp_7_cfg_a; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_7_cfg_x = ptw_io_requestor_2_pmp_7_cfg_x; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_7_cfg_w = ptw_io_requestor_2_pmp_7_cfg_w; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_7_cfg_r = ptw_io_requestor_2_pmp_7_cfg_r; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_7_addr = ptw_io_requestor_2_pmp_7_addr; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_pmp_7_mask = ptw_io_requestor_2_pmp_7_mask; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_customCSRs_csrs_0_wen = ptw_io_requestor_2_customCSRs_csrs_0_wen; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_customCSRs_csrs_0_wdata = ptw_io_requestor_2_customCSRs_csrs_0_wdata; // @[tile.scala 232:20]
  assign core_io_ptw_tlb_customCSRs_csrs_0_value = ptw_io_requestor_2_customCSRs_csrs_0_value; // @[tile.scala 232:20]
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign lsu_io_ptw_req_ready = ptw_io_requestor_0_req_ready; // @[tile.scala 232:20]
  assign lsu_io_ptw_resp_valid = ptw_io_requestor_0_resp_valid; // @[tile.scala 232:20]
  assign lsu_io_ptw_resp_bits_ae = ptw_io_requestor_0_resp_bits_ae; // @[tile.scala 232:20]
  assign lsu_io_ptw_resp_bits_pte_ppn = ptw_io_requestor_0_resp_bits_pte_ppn; // @[tile.scala 232:20]
  assign lsu_io_ptw_resp_bits_pte_reserved_for_software = ptw_io_requestor_0_resp_bits_pte_reserved_for_software; // @[tile.scala 232:20]
  assign lsu_io_ptw_resp_bits_pte_d = ptw_io_requestor_0_resp_bits_pte_d; // @[tile.scala 232:20]
  assign lsu_io_ptw_resp_bits_pte_a = ptw_io_requestor_0_resp_bits_pte_a; // @[tile.scala 232:20]
  assign lsu_io_ptw_resp_bits_pte_g = ptw_io_requestor_0_resp_bits_pte_g; // @[tile.scala 232:20]
  assign lsu_io_ptw_resp_bits_pte_u = ptw_io_requestor_0_resp_bits_pte_u; // @[tile.scala 232:20]
  assign lsu_io_ptw_resp_bits_pte_x = ptw_io_requestor_0_resp_bits_pte_x; // @[tile.scala 232:20]
  assign lsu_io_ptw_resp_bits_pte_w = ptw_io_requestor_0_resp_bits_pte_w; // @[tile.scala 232:20]
  assign lsu_io_ptw_resp_bits_pte_r = ptw_io_requestor_0_resp_bits_pte_r; // @[tile.scala 232:20]
  assign lsu_io_ptw_resp_bits_pte_v = ptw_io_requestor_0_resp_bits_pte_v; // @[tile.scala 232:20]
  assign lsu_io_ptw_resp_bits_level = ptw_io_requestor_0_resp_bits_level; // @[tile.scala 232:20]
  assign lsu_io_ptw_resp_bits_fragmented_superpage = ptw_io_requestor_0_resp_bits_fragmented_superpage; // @[tile.scala 232:20]
  assign lsu_io_ptw_resp_bits_homogeneous = ptw_io_requestor_0_resp_bits_homogeneous; // @[tile.scala 232:20]
  assign lsu_io_ptw_ptbr_mode = ptw_io_requestor_0_ptbr_mode; // @[tile.scala 232:20]
  assign lsu_io_ptw_ptbr_asid = ptw_io_requestor_0_ptbr_asid; // @[tile.scala 232:20]
  assign lsu_io_ptw_ptbr_ppn = ptw_io_requestor_0_ptbr_ppn; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_debug = ptw_io_requestor_0_status_debug; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_cease = ptw_io_requestor_0_status_cease; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_wfi = ptw_io_requestor_0_status_wfi; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_isa = ptw_io_requestor_0_status_isa; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_dprv = ptw_io_requestor_0_status_dprv; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_prv = ptw_io_requestor_0_status_prv; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_sd = ptw_io_requestor_0_status_sd; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_zero2 = ptw_io_requestor_0_status_zero2; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_sxl = ptw_io_requestor_0_status_sxl; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_uxl = ptw_io_requestor_0_status_uxl; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_sd_rv32 = ptw_io_requestor_0_status_sd_rv32; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_zero1 = ptw_io_requestor_0_status_zero1; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_tsr = ptw_io_requestor_0_status_tsr; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_tw = ptw_io_requestor_0_status_tw; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_tvm = ptw_io_requestor_0_status_tvm; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_mxr = ptw_io_requestor_0_status_mxr; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_sum = ptw_io_requestor_0_status_sum; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_mprv = ptw_io_requestor_0_status_mprv; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_xs = ptw_io_requestor_0_status_xs; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_fs = ptw_io_requestor_0_status_fs; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_mpp = ptw_io_requestor_0_status_mpp; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_vs = ptw_io_requestor_0_status_vs; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_spp = ptw_io_requestor_0_status_spp; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_mpie = ptw_io_requestor_0_status_mpie; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_hpie = ptw_io_requestor_0_status_hpie; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_spie = ptw_io_requestor_0_status_spie; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_upie = ptw_io_requestor_0_status_upie; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_mie = ptw_io_requestor_0_status_mie; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_hie = ptw_io_requestor_0_status_hie; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_sie = ptw_io_requestor_0_status_sie; // @[tile.scala 232:20]
  assign lsu_io_ptw_status_uie = ptw_io_requestor_0_status_uie; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_0_cfg_l = ptw_io_requestor_0_pmp_0_cfg_l; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_0_cfg_res = ptw_io_requestor_0_pmp_0_cfg_res; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_0_cfg_a = ptw_io_requestor_0_pmp_0_cfg_a; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_0_cfg_x = ptw_io_requestor_0_pmp_0_cfg_x; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_0_cfg_w = ptw_io_requestor_0_pmp_0_cfg_w; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_0_cfg_r = ptw_io_requestor_0_pmp_0_cfg_r; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_0_addr = ptw_io_requestor_0_pmp_0_addr; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_0_mask = ptw_io_requestor_0_pmp_0_mask; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_1_cfg_l = ptw_io_requestor_0_pmp_1_cfg_l; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_1_cfg_res = ptw_io_requestor_0_pmp_1_cfg_res; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_1_cfg_a = ptw_io_requestor_0_pmp_1_cfg_a; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_1_cfg_x = ptw_io_requestor_0_pmp_1_cfg_x; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_1_cfg_w = ptw_io_requestor_0_pmp_1_cfg_w; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_1_cfg_r = ptw_io_requestor_0_pmp_1_cfg_r; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_1_addr = ptw_io_requestor_0_pmp_1_addr; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_1_mask = ptw_io_requestor_0_pmp_1_mask; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_2_cfg_l = ptw_io_requestor_0_pmp_2_cfg_l; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_2_cfg_res = ptw_io_requestor_0_pmp_2_cfg_res; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_2_cfg_a = ptw_io_requestor_0_pmp_2_cfg_a; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_2_cfg_x = ptw_io_requestor_0_pmp_2_cfg_x; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_2_cfg_w = ptw_io_requestor_0_pmp_2_cfg_w; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_2_cfg_r = ptw_io_requestor_0_pmp_2_cfg_r; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_2_addr = ptw_io_requestor_0_pmp_2_addr; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_2_mask = ptw_io_requestor_0_pmp_2_mask; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_3_cfg_l = ptw_io_requestor_0_pmp_3_cfg_l; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_3_cfg_res = ptw_io_requestor_0_pmp_3_cfg_res; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_3_cfg_a = ptw_io_requestor_0_pmp_3_cfg_a; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_3_cfg_x = ptw_io_requestor_0_pmp_3_cfg_x; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_3_cfg_w = ptw_io_requestor_0_pmp_3_cfg_w; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_3_cfg_r = ptw_io_requestor_0_pmp_3_cfg_r; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_3_addr = ptw_io_requestor_0_pmp_3_addr; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_3_mask = ptw_io_requestor_0_pmp_3_mask; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_4_cfg_l = ptw_io_requestor_0_pmp_4_cfg_l; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_4_cfg_res = ptw_io_requestor_0_pmp_4_cfg_res; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_4_cfg_a = ptw_io_requestor_0_pmp_4_cfg_a; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_4_cfg_x = ptw_io_requestor_0_pmp_4_cfg_x; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_4_cfg_w = ptw_io_requestor_0_pmp_4_cfg_w; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_4_cfg_r = ptw_io_requestor_0_pmp_4_cfg_r; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_4_addr = ptw_io_requestor_0_pmp_4_addr; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_4_mask = ptw_io_requestor_0_pmp_4_mask; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_5_cfg_l = ptw_io_requestor_0_pmp_5_cfg_l; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_5_cfg_res = ptw_io_requestor_0_pmp_5_cfg_res; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_5_cfg_a = ptw_io_requestor_0_pmp_5_cfg_a; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_5_cfg_x = ptw_io_requestor_0_pmp_5_cfg_x; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_5_cfg_w = ptw_io_requestor_0_pmp_5_cfg_w; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_5_cfg_r = ptw_io_requestor_0_pmp_5_cfg_r; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_5_addr = ptw_io_requestor_0_pmp_5_addr; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_5_mask = ptw_io_requestor_0_pmp_5_mask; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_6_cfg_l = ptw_io_requestor_0_pmp_6_cfg_l; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_6_cfg_res = ptw_io_requestor_0_pmp_6_cfg_res; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_6_cfg_a = ptw_io_requestor_0_pmp_6_cfg_a; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_6_cfg_x = ptw_io_requestor_0_pmp_6_cfg_x; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_6_cfg_w = ptw_io_requestor_0_pmp_6_cfg_w; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_6_cfg_r = ptw_io_requestor_0_pmp_6_cfg_r; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_6_addr = ptw_io_requestor_0_pmp_6_addr; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_6_mask = ptw_io_requestor_0_pmp_6_mask; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_7_cfg_l = ptw_io_requestor_0_pmp_7_cfg_l; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_7_cfg_res = ptw_io_requestor_0_pmp_7_cfg_res; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_7_cfg_a = ptw_io_requestor_0_pmp_7_cfg_a; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_7_cfg_x = ptw_io_requestor_0_pmp_7_cfg_x; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_7_cfg_w = ptw_io_requestor_0_pmp_7_cfg_w; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_7_cfg_r = ptw_io_requestor_0_pmp_7_cfg_r; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_7_addr = ptw_io_requestor_0_pmp_7_addr; // @[tile.scala 232:20]
  assign lsu_io_ptw_pmp_7_mask = ptw_io_requestor_0_pmp_7_mask; // @[tile.scala 232:20]
  assign lsu_io_ptw_customCSRs_csrs_0_wen = ptw_io_requestor_0_customCSRs_csrs_0_wen; // @[tile.scala 232:20]
  assign lsu_io_ptw_customCSRs_csrs_0_wdata = ptw_io_requestor_0_customCSRs_csrs_0_wdata; // @[tile.scala 232:20]
  assign lsu_io_ptw_customCSRs_csrs_0_value = ptw_io_requestor_0_customCSRs_csrs_0_value; // @[tile.scala 232:20]
  assign lsu_io_core_exe_0_req_valid = core_io_lsu_exe_0_req_valid; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_switch = core_io_lsu_exe_0_req_bits_uop_switch; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_switch_off = core_io_lsu_exe_0_req_bits_uop_switch_off; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_is_unicore = core_io_lsu_exe_0_req_bits_uop_is_unicore; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_shift = core_io_lsu_exe_0_req_bits_uop_shift; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_lrs3_rtype = core_io_lsu_exe_0_req_bits_uop_lrs3_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_rflag = core_io_lsu_exe_0_req_bits_uop_rflag; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_wflag = core_io_lsu_exe_0_req_bits_uop_wflag; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_prflag = core_io_lsu_exe_0_req_bits_uop_prflag; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_pwflag = core_io_lsu_exe_0_req_bits_uop_pwflag; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_pflag_busy = core_io_lsu_exe_0_req_bits_uop_pflag_busy; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_stale_pflag = core_io_lsu_exe_0_req_bits_uop_stale_pflag; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_op1_sel = core_io_lsu_exe_0_req_bits_uop_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_op2_sel = core_io_lsu_exe_0_req_bits_uop_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_split_num = core_io_lsu_exe_0_req_bits_uop_split_num; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_self_index = core_io_lsu_exe_0_req_bits_uop_self_index; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_rob_inst_idx = core_io_lsu_exe_0_req_bits_uop_rob_inst_idx; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_address_num = core_io_lsu_exe_0_req_bits_uop_address_num; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_uopc = core_io_lsu_exe_0_req_bits_uop_uopc; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_inst = core_io_lsu_exe_0_req_bits_uop_inst; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_debug_inst = core_io_lsu_exe_0_req_bits_uop_debug_inst; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_is_rvc = core_io_lsu_exe_0_req_bits_uop_is_rvc; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_debug_pc = core_io_lsu_exe_0_req_bits_uop_debug_pc; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_iq_type = core_io_lsu_exe_0_req_bits_uop_iq_type; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_fu_code = core_io_lsu_exe_0_req_bits_uop_fu_code; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_ctrl_br_type = core_io_lsu_exe_0_req_bits_uop_ctrl_br_type; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_ctrl_op1_sel = core_io_lsu_exe_0_req_bits_uop_ctrl_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_ctrl_op2_sel = core_io_lsu_exe_0_req_bits_uop_ctrl_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_ctrl_imm_sel = core_io_lsu_exe_0_req_bits_uop_ctrl_imm_sel; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_ctrl_op_fcn = core_io_lsu_exe_0_req_bits_uop_ctrl_op_fcn; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_ctrl_fcn_dw = core_io_lsu_exe_0_req_bits_uop_ctrl_fcn_dw; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_ctrl_csr_cmd = core_io_lsu_exe_0_req_bits_uop_ctrl_csr_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_ctrl_is_load = core_io_lsu_exe_0_req_bits_uop_ctrl_is_load; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_ctrl_is_sta = core_io_lsu_exe_0_req_bits_uop_ctrl_is_sta; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_ctrl_is_std = core_io_lsu_exe_0_req_bits_uop_ctrl_is_std; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_ctrl_op3_sel = core_io_lsu_exe_0_req_bits_uop_ctrl_op3_sel; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_iw_state = core_io_lsu_exe_0_req_bits_uop_iw_state; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_iw_p1_poisoned = core_io_lsu_exe_0_req_bits_uop_iw_p1_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_iw_p2_poisoned = core_io_lsu_exe_0_req_bits_uop_iw_p2_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_is_br = core_io_lsu_exe_0_req_bits_uop_is_br; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_is_jalr = core_io_lsu_exe_0_req_bits_uop_is_jalr; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_is_jal = core_io_lsu_exe_0_req_bits_uop_is_jal; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_is_sfb = core_io_lsu_exe_0_req_bits_uop_is_sfb; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_br_mask = core_io_lsu_exe_0_req_bits_uop_br_mask; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_br_tag = core_io_lsu_exe_0_req_bits_uop_br_tag; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_ftq_idx = core_io_lsu_exe_0_req_bits_uop_ftq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_edge_inst = core_io_lsu_exe_0_req_bits_uop_edge_inst; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_pc_lob = core_io_lsu_exe_0_req_bits_uop_pc_lob; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_taken = core_io_lsu_exe_0_req_bits_uop_taken; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_imm_packed = core_io_lsu_exe_0_req_bits_uop_imm_packed; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_csr_addr = core_io_lsu_exe_0_req_bits_uop_csr_addr; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_rob_idx = core_io_lsu_exe_0_req_bits_uop_rob_idx; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_ldq_idx = core_io_lsu_exe_0_req_bits_uop_ldq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_stq_idx = core_io_lsu_exe_0_req_bits_uop_stq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_rxq_idx = core_io_lsu_exe_0_req_bits_uop_rxq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_pdst = core_io_lsu_exe_0_req_bits_uop_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_prs1 = core_io_lsu_exe_0_req_bits_uop_prs1; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_prs2 = core_io_lsu_exe_0_req_bits_uop_prs2; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_prs3 = core_io_lsu_exe_0_req_bits_uop_prs3; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_ppred = core_io_lsu_exe_0_req_bits_uop_ppred; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_prs1_busy = core_io_lsu_exe_0_req_bits_uop_prs1_busy; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_prs2_busy = core_io_lsu_exe_0_req_bits_uop_prs2_busy; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_prs3_busy = core_io_lsu_exe_0_req_bits_uop_prs3_busy; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_ppred_busy = core_io_lsu_exe_0_req_bits_uop_ppred_busy; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_stale_pdst = core_io_lsu_exe_0_req_bits_uop_stale_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_exception = core_io_lsu_exe_0_req_bits_uop_exception; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_exc_cause = core_io_lsu_exe_0_req_bits_uop_exc_cause; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_bypassable = core_io_lsu_exe_0_req_bits_uop_bypassable; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_mem_cmd = core_io_lsu_exe_0_req_bits_uop_mem_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_mem_size = core_io_lsu_exe_0_req_bits_uop_mem_size; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_mem_signed = core_io_lsu_exe_0_req_bits_uop_mem_signed; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_is_fence = core_io_lsu_exe_0_req_bits_uop_is_fence; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_is_fencei = core_io_lsu_exe_0_req_bits_uop_is_fencei; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_is_amo = core_io_lsu_exe_0_req_bits_uop_is_amo; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_uses_ldq = core_io_lsu_exe_0_req_bits_uop_uses_ldq; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_uses_stq = core_io_lsu_exe_0_req_bits_uop_uses_stq; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_is_sys_pc2epc = core_io_lsu_exe_0_req_bits_uop_is_sys_pc2epc; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_is_unique = core_io_lsu_exe_0_req_bits_uop_is_unique; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_flush_on_commit = core_io_lsu_exe_0_req_bits_uop_flush_on_commit; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_ldst_is_rs1 = core_io_lsu_exe_0_req_bits_uop_ldst_is_rs1; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_ldst = core_io_lsu_exe_0_req_bits_uop_ldst; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_lrs1 = core_io_lsu_exe_0_req_bits_uop_lrs1; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_lrs2 = core_io_lsu_exe_0_req_bits_uop_lrs2; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_lrs3 = core_io_lsu_exe_0_req_bits_uop_lrs3; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_ldst_val = core_io_lsu_exe_0_req_bits_uop_ldst_val; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_dst_rtype = core_io_lsu_exe_0_req_bits_uop_dst_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_lrs1_rtype = core_io_lsu_exe_0_req_bits_uop_lrs1_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_lrs2_rtype = core_io_lsu_exe_0_req_bits_uop_lrs2_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_frs3_en = core_io_lsu_exe_0_req_bits_uop_frs3_en; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_fp_val = core_io_lsu_exe_0_req_bits_uop_fp_val; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_fp_single = core_io_lsu_exe_0_req_bits_uop_fp_single; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_xcpt_pf_if = core_io_lsu_exe_0_req_bits_uop_xcpt_pf_if; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_xcpt_ae_if = core_io_lsu_exe_0_req_bits_uop_xcpt_ae_if; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_xcpt_ma_if = core_io_lsu_exe_0_req_bits_uop_xcpt_ma_if; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_bp_debug_if = core_io_lsu_exe_0_req_bits_uop_bp_debug_if; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_bp_xcpt_if = core_io_lsu_exe_0_req_bits_uop_bp_xcpt_if; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_debug_fsrc = core_io_lsu_exe_0_req_bits_uop_debug_fsrc; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_uop_debug_tsrc = core_io_lsu_exe_0_req_bits_uop_debug_tsrc; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_predicated = core_io_lsu_exe_0_req_bits_predicated; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_data = core_io_lsu_exe_0_req_bits_data; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_valid = core_io_lsu_exe_0_req_bits_fflags_valid; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_switch = core_io_lsu_exe_0_req_bits_fflags_bits_uop_switch; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_switch_off = core_io_lsu_exe_0_req_bits_fflags_bits_uop_switch_off; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_unicore = core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_unicore; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_shift = core_io_lsu_exe_0_req_bits_fflags_bits_uop_shift; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_lrs3_rtype = core_io_lsu_exe_0_req_bits_fflags_bits_uop_lrs3_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_rflag = core_io_lsu_exe_0_req_bits_fflags_bits_uop_rflag; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_wflag = core_io_lsu_exe_0_req_bits_fflags_bits_uop_wflag; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_prflag = core_io_lsu_exe_0_req_bits_fflags_bits_uop_prflag; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_pwflag = core_io_lsu_exe_0_req_bits_fflags_bits_uop_pwflag; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_pflag_busy = core_io_lsu_exe_0_req_bits_fflags_bits_uop_pflag_busy; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_stale_pflag = core_io_lsu_exe_0_req_bits_fflags_bits_uop_stale_pflag
    ; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_op1_sel = core_io_lsu_exe_0_req_bits_fflags_bits_uop_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_op2_sel = core_io_lsu_exe_0_req_bits_fflags_bits_uop_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_split_num = core_io_lsu_exe_0_req_bits_fflags_bits_uop_split_num; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_self_index = core_io_lsu_exe_0_req_bits_fflags_bits_uop_self_index; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_rob_inst_idx =
    core_io_lsu_exe_0_req_bits_fflags_bits_uop_rob_inst_idx; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_address_num = core_io_lsu_exe_0_req_bits_fflags_bits_uop_address_num
    ; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_uopc = core_io_lsu_exe_0_req_bits_fflags_bits_uop_uopc; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_inst = core_io_lsu_exe_0_req_bits_fflags_bits_uop_inst; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_debug_inst = core_io_lsu_exe_0_req_bits_fflags_bits_uop_debug_inst; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_rvc = core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_rvc; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_debug_pc = core_io_lsu_exe_0_req_bits_fflags_bits_uop_debug_pc; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_iq_type = core_io_lsu_exe_0_req_bits_fflags_bits_uop_iq_type; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_fu_code = core_io_lsu_exe_0_req_bits_fflags_bits_uop_fu_code; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_br_type =
    core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_br_type; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_op1_sel =
    core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_op2_sel =
    core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_imm_sel =
    core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_imm_sel; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_op_fcn = core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_op_fcn
    ; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_fcn_dw = core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_fcn_dw
    ; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_csr_cmd =
    core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_csr_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_is_load =
    core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_is_load; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_is_sta = core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_is_sta
    ; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_is_std = core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_is_std
    ; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_ctrl_op3_sel =
    core_io_lsu_exe_0_req_bits_fflags_bits_uop_ctrl_op3_sel; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_iw_state = core_io_lsu_exe_0_req_bits_fflags_bits_uop_iw_state; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_iw_p1_poisoned =
    core_io_lsu_exe_0_req_bits_fflags_bits_uop_iw_p1_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_iw_p2_poisoned =
    core_io_lsu_exe_0_req_bits_fflags_bits_uop_iw_p2_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_br = core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_br; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_jalr = core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_jalr; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_jal = core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_jal; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_sfb = core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_sfb; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_br_mask = core_io_lsu_exe_0_req_bits_fflags_bits_uop_br_mask; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_br_tag = core_io_lsu_exe_0_req_bits_fflags_bits_uop_br_tag; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_ftq_idx = core_io_lsu_exe_0_req_bits_fflags_bits_uop_ftq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_edge_inst = core_io_lsu_exe_0_req_bits_fflags_bits_uop_edge_inst; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_pc_lob = core_io_lsu_exe_0_req_bits_fflags_bits_uop_pc_lob; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_taken = core_io_lsu_exe_0_req_bits_fflags_bits_uop_taken; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_imm_packed = core_io_lsu_exe_0_req_bits_fflags_bits_uop_imm_packed; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_csr_addr = core_io_lsu_exe_0_req_bits_fflags_bits_uop_csr_addr; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_rob_idx = core_io_lsu_exe_0_req_bits_fflags_bits_uop_rob_idx; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_ldq_idx = core_io_lsu_exe_0_req_bits_fflags_bits_uop_ldq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_stq_idx = core_io_lsu_exe_0_req_bits_fflags_bits_uop_stq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_rxq_idx = core_io_lsu_exe_0_req_bits_fflags_bits_uop_rxq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_pdst = core_io_lsu_exe_0_req_bits_fflags_bits_uop_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_prs1 = core_io_lsu_exe_0_req_bits_fflags_bits_uop_prs1; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_prs2 = core_io_lsu_exe_0_req_bits_fflags_bits_uop_prs2; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_prs3 = core_io_lsu_exe_0_req_bits_fflags_bits_uop_prs3; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_ppred = core_io_lsu_exe_0_req_bits_fflags_bits_uop_ppred; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_prs1_busy = core_io_lsu_exe_0_req_bits_fflags_bits_uop_prs1_busy; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_prs2_busy = core_io_lsu_exe_0_req_bits_fflags_bits_uop_prs2_busy; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_prs3_busy = core_io_lsu_exe_0_req_bits_fflags_bits_uop_prs3_busy; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_ppred_busy = core_io_lsu_exe_0_req_bits_fflags_bits_uop_ppred_busy; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_stale_pdst = core_io_lsu_exe_0_req_bits_fflags_bits_uop_stale_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_exception = core_io_lsu_exe_0_req_bits_fflags_bits_uop_exception; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_exc_cause = core_io_lsu_exe_0_req_bits_fflags_bits_uop_exc_cause; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_bypassable = core_io_lsu_exe_0_req_bits_fflags_bits_uop_bypassable; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_mem_cmd = core_io_lsu_exe_0_req_bits_fflags_bits_uop_mem_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_mem_size = core_io_lsu_exe_0_req_bits_fflags_bits_uop_mem_size; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_mem_signed = core_io_lsu_exe_0_req_bits_fflags_bits_uop_mem_signed; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_fence = core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_fence; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_fencei = core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_fencei; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_amo = core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_amo; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_uses_ldq = core_io_lsu_exe_0_req_bits_fflags_bits_uop_uses_ldq; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_uses_stq = core_io_lsu_exe_0_req_bits_fflags_bits_uop_uses_stq; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_sys_pc2epc =
    core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_sys_pc2epc; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_is_unique = core_io_lsu_exe_0_req_bits_fflags_bits_uop_is_unique; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_flush_on_commit =
    core_io_lsu_exe_0_req_bits_fflags_bits_uop_flush_on_commit; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_ldst_is_rs1 = core_io_lsu_exe_0_req_bits_fflags_bits_uop_ldst_is_rs1
    ; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_ldst = core_io_lsu_exe_0_req_bits_fflags_bits_uop_ldst; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_lrs1 = core_io_lsu_exe_0_req_bits_fflags_bits_uop_lrs1; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_lrs2 = core_io_lsu_exe_0_req_bits_fflags_bits_uop_lrs2; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_lrs3 = core_io_lsu_exe_0_req_bits_fflags_bits_uop_lrs3; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_ldst_val = core_io_lsu_exe_0_req_bits_fflags_bits_uop_ldst_val; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_dst_rtype = core_io_lsu_exe_0_req_bits_fflags_bits_uop_dst_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_lrs1_rtype = core_io_lsu_exe_0_req_bits_fflags_bits_uop_lrs1_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_lrs2_rtype = core_io_lsu_exe_0_req_bits_fflags_bits_uop_lrs2_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_frs3_en = core_io_lsu_exe_0_req_bits_fflags_bits_uop_frs3_en; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_fp_val = core_io_lsu_exe_0_req_bits_fflags_bits_uop_fp_val; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_fp_single = core_io_lsu_exe_0_req_bits_fflags_bits_uop_fp_single; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_xcpt_pf_if = core_io_lsu_exe_0_req_bits_fflags_bits_uop_xcpt_pf_if; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_xcpt_ae_if = core_io_lsu_exe_0_req_bits_fflags_bits_uop_xcpt_ae_if; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_xcpt_ma_if = core_io_lsu_exe_0_req_bits_fflags_bits_uop_xcpt_ma_if; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_bp_debug_if = core_io_lsu_exe_0_req_bits_fflags_bits_uop_bp_debug_if
    ; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_bp_xcpt_if = core_io_lsu_exe_0_req_bits_fflags_bits_uop_bp_xcpt_if; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_debug_fsrc = core_io_lsu_exe_0_req_bits_fflags_bits_uop_debug_fsrc; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_uop_debug_tsrc = core_io_lsu_exe_0_req_bits_fflags_bits_uop_debug_tsrc; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflags_bits_flags = core_io_lsu_exe_0_req_bits_fflags_bits_flags; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_addr = core_io_lsu_exe_0_req_bits_addr; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_mxcpt_valid = core_io_lsu_exe_0_req_bits_mxcpt_valid; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_mxcpt_bits = core_io_lsu_exe_0_req_bits_mxcpt_bits; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_sfence_valid = core_io_lsu_exe_0_req_bits_sfence_valid; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_sfence_bits_rs1 = core_io_lsu_exe_0_req_bits_sfence_bits_rs1; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_sfence_bits_rs2 = core_io_lsu_exe_0_req_bits_sfence_bits_rs2; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_sfence_bits_addr = core_io_lsu_exe_0_req_bits_sfence_bits_addr; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_sfence_bits_asid = core_io_lsu_exe_0_req_bits_sfence_bits_asid; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_flagdata = core_io_lsu_exe_0_req_bits_flagdata; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_valid = core_io_lsu_exe_0_req_bits_fflagdata_valid; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_switch = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_switch; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_switch_off =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_switch_off; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_unicore =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_unicore; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_shift = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_shift; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_lrs3_rtype =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs3_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_rflag = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_rflag; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_wflag = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_wflag; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_prflag = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_prflag; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_pwflag = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_pwflag; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_pflag_busy =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_pflag_busy; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_stale_pflag =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_stale_pflag; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_op1_sel = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_op2_sel = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_split_num =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_split_num; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_self_index =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_self_index; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_rob_inst_idx =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_rob_inst_idx; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_address_num =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_address_num; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_uopc = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_uopc; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_inst = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_inst; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_debug_inst =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_debug_inst; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_rvc = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_rvc; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_debug_pc = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_debug_pc
    ; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_iq_type = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_iq_type; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_fu_code = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_fu_code; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_br_type =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_br_type; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_op1_sel =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_op2_sel =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_imm_sel =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_imm_sel; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_op_fcn =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_op_fcn; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_fcn_dw =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_fcn_dw; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_csr_cmd =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_csr_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_load =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_load; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_sta =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_sta; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_std =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_is_std; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ctrl_op3_sel =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ctrl_op3_sel; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_iw_state = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_iw_state
    ; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_iw_p1_poisoned =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_iw_p1_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_iw_p2_poisoned =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_iw_p2_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_br = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_br; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_jalr = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_jalr; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_jal = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_jal; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_sfb = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_sfb; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_br_mask = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_br_mask; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_br_tag = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_br_tag; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ftq_idx = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ftq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_edge_inst =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_edge_inst; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_pc_lob = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_pc_lob; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_taken = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_taken; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_imm_packed =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_imm_packed; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_csr_addr = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_csr_addr
    ; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_rob_idx = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_rob_idx; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ldq_idx = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ldq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_stq_idx = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_stq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_rxq_idx = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_rxq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_pdst = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_prs1 = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs1; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_prs2 = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs2; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_prs3 = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs3; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ppred = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ppred; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_prs1_busy =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs1_busy; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_prs2_busy =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs2_busy; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_prs3_busy =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_prs3_busy; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ppred_busy =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ppred_busy; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_stale_pdst =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_stale_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_exception =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_exception; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_exc_cause =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_exc_cause; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_bypassable =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_bypassable; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_mem_cmd = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_mem_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_mem_size = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_mem_size
    ; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_mem_signed =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_mem_signed; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_fence = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_fence
    ; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_fencei =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_fencei; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_amo = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_amo; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_uses_ldq = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_uses_ldq
    ; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_uses_stq = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_uses_stq
    ; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_sys_pc2epc =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_sys_pc2epc; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_is_unique =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_is_unique; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_flush_on_commit =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_flush_on_commit; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ldst_is_rs1 =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ldst_is_rs1; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ldst = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ldst; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_lrs1 = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs1; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_lrs2 = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs2; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_lrs3 = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs3; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_ldst_val = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_ldst_val
    ; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_dst_rtype =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_dst_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_lrs1_rtype =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs1_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_lrs2_rtype =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_lrs2_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_frs3_en = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_frs3_en; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_fp_val = core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_fp_val; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_fp_single =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_fp_single; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_xcpt_pf_if =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_xcpt_pf_if; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_xcpt_ae_if =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_xcpt_ae_if; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_xcpt_ma_if =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_xcpt_ma_if; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_bp_debug_if =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_bp_debug_if; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_bp_xcpt_if =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_bp_xcpt_if; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_debug_fsrc =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_debug_fsrc; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_uop_debug_tsrc =
    core_io_lsu_exe_0_req_bits_fflagdata_bits_uop_debug_tsrc; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_req_bits_fflagdata_bits_fflag = core_io_lsu_exe_0_req_bits_fflagdata_bits_fflag; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_iresp_ready = core_io_lsu_exe_0_iresp_ready; // @[tile.scala 178:15]
  assign lsu_io_core_exe_0_fresp_ready = core_io_lsu_exe_0_fresp_ready; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_valid = core_io_lsu_dis_uops_0_valid; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_switch = core_io_lsu_dis_uops_0_bits_switch; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_switch_off = core_io_lsu_dis_uops_0_bits_switch_off; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_is_unicore = core_io_lsu_dis_uops_0_bits_is_unicore; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_shift = core_io_lsu_dis_uops_0_bits_shift; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_lrs3_rtype = core_io_lsu_dis_uops_0_bits_lrs3_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_rflag = core_io_lsu_dis_uops_0_bits_rflag; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_wflag = core_io_lsu_dis_uops_0_bits_wflag; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_prflag = core_io_lsu_dis_uops_0_bits_prflag; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_pwflag = core_io_lsu_dis_uops_0_bits_pwflag; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_pflag_busy = core_io_lsu_dis_uops_0_bits_pflag_busy; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_stale_pflag = core_io_lsu_dis_uops_0_bits_stale_pflag; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_op1_sel = core_io_lsu_dis_uops_0_bits_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_op2_sel = core_io_lsu_dis_uops_0_bits_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_split_num = core_io_lsu_dis_uops_0_bits_split_num; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_self_index = core_io_lsu_dis_uops_0_bits_self_index; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_rob_inst_idx = core_io_lsu_dis_uops_0_bits_rob_inst_idx; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_address_num = core_io_lsu_dis_uops_0_bits_address_num; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_uopc = core_io_lsu_dis_uops_0_bits_uopc; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_inst = core_io_lsu_dis_uops_0_bits_inst; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_debug_inst = core_io_lsu_dis_uops_0_bits_debug_inst; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_is_rvc = core_io_lsu_dis_uops_0_bits_is_rvc; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_debug_pc = core_io_lsu_dis_uops_0_bits_debug_pc; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_iq_type = core_io_lsu_dis_uops_0_bits_iq_type; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_fu_code = core_io_lsu_dis_uops_0_bits_fu_code; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_ctrl_br_type = core_io_lsu_dis_uops_0_bits_ctrl_br_type; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_ctrl_op1_sel = core_io_lsu_dis_uops_0_bits_ctrl_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_ctrl_op2_sel = core_io_lsu_dis_uops_0_bits_ctrl_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_ctrl_imm_sel = core_io_lsu_dis_uops_0_bits_ctrl_imm_sel; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_ctrl_op_fcn = core_io_lsu_dis_uops_0_bits_ctrl_op_fcn; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_ctrl_fcn_dw = core_io_lsu_dis_uops_0_bits_ctrl_fcn_dw; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_ctrl_csr_cmd = core_io_lsu_dis_uops_0_bits_ctrl_csr_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_ctrl_is_load = core_io_lsu_dis_uops_0_bits_ctrl_is_load; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_ctrl_is_sta = core_io_lsu_dis_uops_0_bits_ctrl_is_sta; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_ctrl_is_std = core_io_lsu_dis_uops_0_bits_ctrl_is_std; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_ctrl_op3_sel = core_io_lsu_dis_uops_0_bits_ctrl_op3_sel; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_iw_state = core_io_lsu_dis_uops_0_bits_iw_state; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_iw_p1_poisoned = core_io_lsu_dis_uops_0_bits_iw_p1_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_iw_p2_poisoned = core_io_lsu_dis_uops_0_bits_iw_p2_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_is_br = core_io_lsu_dis_uops_0_bits_is_br; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_is_jalr = core_io_lsu_dis_uops_0_bits_is_jalr; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_is_jal = core_io_lsu_dis_uops_0_bits_is_jal; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_is_sfb = core_io_lsu_dis_uops_0_bits_is_sfb; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_br_mask = core_io_lsu_dis_uops_0_bits_br_mask; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_br_tag = core_io_lsu_dis_uops_0_bits_br_tag; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_ftq_idx = core_io_lsu_dis_uops_0_bits_ftq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_edge_inst = core_io_lsu_dis_uops_0_bits_edge_inst; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_pc_lob = core_io_lsu_dis_uops_0_bits_pc_lob; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_taken = core_io_lsu_dis_uops_0_bits_taken; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_imm_packed = core_io_lsu_dis_uops_0_bits_imm_packed; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_csr_addr = core_io_lsu_dis_uops_0_bits_csr_addr; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_rob_idx = core_io_lsu_dis_uops_0_bits_rob_idx; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_ldq_idx = core_io_lsu_dis_uops_0_bits_ldq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_stq_idx = core_io_lsu_dis_uops_0_bits_stq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_rxq_idx = core_io_lsu_dis_uops_0_bits_rxq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_pdst = core_io_lsu_dis_uops_0_bits_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_prs1 = core_io_lsu_dis_uops_0_bits_prs1; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_prs2 = core_io_lsu_dis_uops_0_bits_prs2; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_prs3 = core_io_lsu_dis_uops_0_bits_prs3; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_ppred = core_io_lsu_dis_uops_0_bits_ppred; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_prs1_busy = core_io_lsu_dis_uops_0_bits_prs1_busy; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_prs2_busy = core_io_lsu_dis_uops_0_bits_prs2_busy; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_prs3_busy = core_io_lsu_dis_uops_0_bits_prs3_busy; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_ppred_busy = core_io_lsu_dis_uops_0_bits_ppred_busy; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_stale_pdst = core_io_lsu_dis_uops_0_bits_stale_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_exception = core_io_lsu_dis_uops_0_bits_exception; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_exc_cause = core_io_lsu_dis_uops_0_bits_exc_cause; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_bypassable = core_io_lsu_dis_uops_0_bits_bypassable; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_mem_cmd = core_io_lsu_dis_uops_0_bits_mem_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_mem_size = core_io_lsu_dis_uops_0_bits_mem_size; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_mem_signed = core_io_lsu_dis_uops_0_bits_mem_signed; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_is_fence = core_io_lsu_dis_uops_0_bits_is_fence; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_is_fencei = core_io_lsu_dis_uops_0_bits_is_fencei; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_is_amo = core_io_lsu_dis_uops_0_bits_is_amo; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_uses_ldq = core_io_lsu_dis_uops_0_bits_uses_ldq; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_uses_stq = core_io_lsu_dis_uops_0_bits_uses_stq; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_is_sys_pc2epc = core_io_lsu_dis_uops_0_bits_is_sys_pc2epc; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_is_unique = core_io_lsu_dis_uops_0_bits_is_unique; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_flush_on_commit = core_io_lsu_dis_uops_0_bits_flush_on_commit; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_ldst_is_rs1 = core_io_lsu_dis_uops_0_bits_ldst_is_rs1; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_ldst = core_io_lsu_dis_uops_0_bits_ldst; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_lrs1 = core_io_lsu_dis_uops_0_bits_lrs1; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_lrs2 = core_io_lsu_dis_uops_0_bits_lrs2; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_lrs3 = core_io_lsu_dis_uops_0_bits_lrs3; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_ldst_val = core_io_lsu_dis_uops_0_bits_ldst_val; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_dst_rtype = core_io_lsu_dis_uops_0_bits_dst_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_lrs1_rtype = core_io_lsu_dis_uops_0_bits_lrs1_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_lrs2_rtype = core_io_lsu_dis_uops_0_bits_lrs2_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_frs3_en = core_io_lsu_dis_uops_0_bits_frs3_en; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_fp_val = core_io_lsu_dis_uops_0_bits_fp_val; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_fp_single = core_io_lsu_dis_uops_0_bits_fp_single; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_xcpt_pf_if = core_io_lsu_dis_uops_0_bits_xcpt_pf_if; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_xcpt_ae_if = core_io_lsu_dis_uops_0_bits_xcpt_ae_if; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_xcpt_ma_if = core_io_lsu_dis_uops_0_bits_xcpt_ma_if; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_bp_debug_if = core_io_lsu_dis_uops_0_bits_bp_debug_if; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_bp_xcpt_if = core_io_lsu_dis_uops_0_bits_bp_xcpt_if; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_debug_fsrc = core_io_lsu_dis_uops_0_bits_debug_fsrc; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_0_bits_debug_tsrc = core_io_lsu_dis_uops_0_bits_debug_tsrc; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_valid = core_io_lsu_dis_uops_1_valid; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_switch = core_io_lsu_dis_uops_1_bits_switch; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_switch_off = core_io_lsu_dis_uops_1_bits_switch_off; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_is_unicore = core_io_lsu_dis_uops_1_bits_is_unicore; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_shift = core_io_lsu_dis_uops_1_bits_shift; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_lrs3_rtype = core_io_lsu_dis_uops_1_bits_lrs3_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_rflag = core_io_lsu_dis_uops_1_bits_rflag; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_wflag = core_io_lsu_dis_uops_1_bits_wflag; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_prflag = core_io_lsu_dis_uops_1_bits_prflag; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_pwflag = core_io_lsu_dis_uops_1_bits_pwflag; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_pflag_busy = core_io_lsu_dis_uops_1_bits_pflag_busy; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_stale_pflag = core_io_lsu_dis_uops_1_bits_stale_pflag; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_op1_sel = core_io_lsu_dis_uops_1_bits_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_op2_sel = core_io_lsu_dis_uops_1_bits_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_split_num = core_io_lsu_dis_uops_1_bits_split_num; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_self_index = core_io_lsu_dis_uops_1_bits_self_index; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_rob_inst_idx = core_io_lsu_dis_uops_1_bits_rob_inst_idx; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_address_num = core_io_lsu_dis_uops_1_bits_address_num; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_uopc = core_io_lsu_dis_uops_1_bits_uopc; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_inst = core_io_lsu_dis_uops_1_bits_inst; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_debug_inst = core_io_lsu_dis_uops_1_bits_debug_inst; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_is_rvc = core_io_lsu_dis_uops_1_bits_is_rvc; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_debug_pc = core_io_lsu_dis_uops_1_bits_debug_pc; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_iq_type = core_io_lsu_dis_uops_1_bits_iq_type; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_fu_code = core_io_lsu_dis_uops_1_bits_fu_code; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_ctrl_br_type = core_io_lsu_dis_uops_1_bits_ctrl_br_type; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_ctrl_op1_sel = core_io_lsu_dis_uops_1_bits_ctrl_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_ctrl_op2_sel = core_io_lsu_dis_uops_1_bits_ctrl_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_ctrl_imm_sel = core_io_lsu_dis_uops_1_bits_ctrl_imm_sel; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_ctrl_op_fcn = core_io_lsu_dis_uops_1_bits_ctrl_op_fcn; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_ctrl_fcn_dw = core_io_lsu_dis_uops_1_bits_ctrl_fcn_dw; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_ctrl_csr_cmd = core_io_lsu_dis_uops_1_bits_ctrl_csr_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_ctrl_is_load = core_io_lsu_dis_uops_1_bits_ctrl_is_load; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_ctrl_is_sta = core_io_lsu_dis_uops_1_bits_ctrl_is_sta; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_ctrl_is_std = core_io_lsu_dis_uops_1_bits_ctrl_is_std; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_ctrl_op3_sel = core_io_lsu_dis_uops_1_bits_ctrl_op3_sel; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_iw_state = core_io_lsu_dis_uops_1_bits_iw_state; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_iw_p1_poisoned = core_io_lsu_dis_uops_1_bits_iw_p1_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_iw_p2_poisoned = core_io_lsu_dis_uops_1_bits_iw_p2_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_is_br = core_io_lsu_dis_uops_1_bits_is_br; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_is_jalr = core_io_lsu_dis_uops_1_bits_is_jalr; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_is_jal = core_io_lsu_dis_uops_1_bits_is_jal; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_is_sfb = core_io_lsu_dis_uops_1_bits_is_sfb; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_br_mask = core_io_lsu_dis_uops_1_bits_br_mask; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_br_tag = core_io_lsu_dis_uops_1_bits_br_tag; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_ftq_idx = core_io_lsu_dis_uops_1_bits_ftq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_edge_inst = core_io_lsu_dis_uops_1_bits_edge_inst; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_pc_lob = core_io_lsu_dis_uops_1_bits_pc_lob; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_taken = core_io_lsu_dis_uops_1_bits_taken; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_imm_packed = core_io_lsu_dis_uops_1_bits_imm_packed; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_csr_addr = core_io_lsu_dis_uops_1_bits_csr_addr; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_rob_idx = core_io_lsu_dis_uops_1_bits_rob_idx; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_ldq_idx = core_io_lsu_dis_uops_1_bits_ldq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_stq_idx = core_io_lsu_dis_uops_1_bits_stq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_rxq_idx = core_io_lsu_dis_uops_1_bits_rxq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_pdst = core_io_lsu_dis_uops_1_bits_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_prs1 = core_io_lsu_dis_uops_1_bits_prs1; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_prs2 = core_io_lsu_dis_uops_1_bits_prs2; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_prs3 = core_io_lsu_dis_uops_1_bits_prs3; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_ppred = core_io_lsu_dis_uops_1_bits_ppred; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_prs1_busy = core_io_lsu_dis_uops_1_bits_prs1_busy; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_prs2_busy = core_io_lsu_dis_uops_1_bits_prs2_busy; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_prs3_busy = core_io_lsu_dis_uops_1_bits_prs3_busy; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_ppred_busy = core_io_lsu_dis_uops_1_bits_ppred_busy; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_stale_pdst = core_io_lsu_dis_uops_1_bits_stale_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_exception = core_io_lsu_dis_uops_1_bits_exception; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_exc_cause = core_io_lsu_dis_uops_1_bits_exc_cause; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_bypassable = core_io_lsu_dis_uops_1_bits_bypassable; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_mem_cmd = core_io_lsu_dis_uops_1_bits_mem_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_mem_size = core_io_lsu_dis_uops_1_bits_mem_size; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_mem_signed = core_io_lsu_dis_uops_1_bits_mem_signed; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_is_fence = core_io_lsu_dis_uops_1_bits_is_fence; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_is_fencei = core_io_lsu_dis_uops_1_bits_is_fencei; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_is_amo = core_io_lsu_dis_uops_1_bits_is_amo; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_uses_ldq = core_io_lsu_dis_uops_1_bits_uses_ldq; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_uses_stq = core_io_lsu_dis_uops_1_bits_uses_stq; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_is_sys_pc2epc = core_io_lsu_dis_uops_1_bits_is_sys_pc2epc; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_is_unique = core_io_lsu_dis_uops_1_bits_is_unique; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_flush_on_commit = core_io_lsu_dis_uops_1_bits_flush_on_commit; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_ldst_is_rs1 = core_io_lsu_dis_uops_1_bits_ldst_is_rs1; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_ldst = core_io_lsu_dis_uops_1_bits_ldst; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_lrs1 = core_io_lsu_dis_uops_1_bits_lrs1; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_lrs2 = core_io_lsu_dis_uops_1_bits_lrs2; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_lrs3 = core_io_lsu_dis_uops_1_bits_lrs3; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_ldst_val = core_io_lsu_dis_uops_1_bits_ldst_val; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_dst_rtype = core_io_lsu_dis_uops_1_bits_dst_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_lrs1_rtype = core_io_lsu_dis_uops_1_bits_lrs1_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_lrs2_rtype = core_io_lsu_dis_uops_1_bits_lrs2_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_frs3_en = core_io_lsu_dis_uops_1_bits_frs3_en; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_fp_val = core_io_lsu_dis_uops_1_bits_fp_val; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_fp_single = core_io_lsu_dis_uops_1_bits_fp_single; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_xcpt_pf_if = core_io_lsu_dis_uops_1_bits_xcpt_pf_if; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_xcpt_ae_if = core_io_lsu_dis_uops_1_bits_xcpt_ae_if; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_xcpt_ma_if = core_io_lsu_dis_uops_1_bits_xcpt_ma_if; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_bp_debug_if = core_io_lsu_dis_uops_1_bits_bp_debug_if; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_bp_xcpt_if = core_io_lsu_dis_uops_1_bits_bp_xcpt_if; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_debug_fsrc = core_io_lsu_dis_uops_1_bits_debug_fsrc; // @[tile.scala 178:15]
  assign lsu_io_core_dis_uops_1_bits_debug_tsrc = core_io_lsu_dis_uops_1_bits_debug_tsrc; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_valid = core_io_lsu_fp_stdata_valid; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_switch = core_io_lsu_fp_stdata_bits_uop_switch; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_switch_off = core_io_lsu_fp_stdata_bits_uop_switch_off; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_is_unicore = core_io_lsu_fp_stdata_bits_uop_is_unicore; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_shift = core_io_lsu_fp_stdata_bits_uop_shift; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_lrs3_rtype = core_io_lsu_fp_stdata_bits_uop_lrs3_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_rflag = core_io_lsu_fp_stdata_bits_uop_rflag; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_wflag = core_io_lsu_fp_stdata_bits_uop_wflag; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_prflag = core_io_lsu_fp_stdata_bits_uop_prflag; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_pwflag = core_io_lsu_fp_stdata_bits_uop_pwflag; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_pflag_busy = core_io_lsu_fp_stdata_bits_uop_pflag_busy; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_stale_pflag = core_io_lsu_fp_stdata_bits_uop_stale_pflag; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_op1_sel = core_io_lsu_fp_stdata_bits_uop_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_op2_sel = core_io_lsu_fp_stdata_bits_uop_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_split_num = core_io_lsu_fp_stdata_bits_uop_split_num; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_self_index = core_io_lsu_fp_stdata_bits_uop_self_index; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_rob_inst_idx = core_io_lsu_fp_stdata_bits_uop_rob_inst_idx; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_address_num = core_io_lsu_fp_stdata_bits_uop_address_num; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_uopc = core_io_lsu_fp_stdata_bits_uop_uopc; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_inst = core_io_lsu_fp_stdata_bits_uop_inst; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_debug_inst = core_io_lsu_fp_stdata_bits_uop_debug_inst; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_is_rvc = core_io_lsu_fp_stdata_bits_uop_is_rvc; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_debug_pc = core_io_lsu_fp_stdata_bits_uop_debug_pc; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_iq_type = core_io_lsu_fp_stdata_bits_uop_iq_type; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_fu_code = core_io_lsu_fp_stdata_bits_uop_fu_code; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_ctrl_br_type = core_io_lsu_fp_stdata_bits_uop_ctrl_br_type; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_ctrl_op1_sel = core_io_lsu_fp_stdata_bits_uop_ctrl_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_ctrl_op2_sel = core_io_lsu_fp_stdata_bits_uop_ctrl_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_ctrl_imm_sel = core_io_lsu_fp_stdata_bits_uop_ctrl_imm_sel; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_ctrl_op_fcn = core_io_lsu_fp_stdata_bits_uop_ctrl_op_fcn; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_ctrl_fcn_dw = core_io_lsu_fp_stdata_bits_uop_ctrl_fcn_dw; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_ctrl_csr_cmd = core_io_lsu_fp_stdata_bits_uop_ctrl_csr_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_ctrl_is_load = core_io_lsu_fp_stdata_bits_uop_ctrl_is_load; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_ctrl_is_sta = core_io_lsu_fp_stdata_bits_uop_ctrl_is_sta; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_ctrl_is_std = core_io_lsu_fp_stdata_bits_uop_ctrl_is_std; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_ctrl_op3_sel = core_io_lsu_fp_stdata_bits_uop_ctrl_op3_sel; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_iw_state = core_io_lsu_fp_stdata_bits_uop_iw_state; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_iw_p1_poisoned = core_io_lsu_fp_stdata_bits_uop_iw_p1_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_iw_p2_poisoned = core_io_lsu_fp_stdata_bits_uop_iw_p2_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_is_br = core_io_lsu_fp_stdata_bits_uop_is_br; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_is_jalr = core_io_lsu_fp_stdata_bits_uop_is_jalr; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_is_jal = core_io_lsu_fp_stdata_bits_uop_is_jal; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_is_sfb = core_io_lsu_fp_stdata_bits_uop_is_sfb; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_br_mask = core_io_lsu_fp_stdata_bits_uop_br_mask; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_br_tag = core_io_lsu_fp_stdata_bits_uop_br_tag; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_ftq_idx = core_io_lsu_fp_stdata_bits_uop_ftq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_edge_inst = core_io_lsu_fp_stdata_bits_uop_edge_inst; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_pc_lob = core_io_lsu_fp_stdata_bits_uop_pc_lob; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_taken = core_io_lsu_fp_stdata_bits_uop_taken; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_imm_packed = core_io_lsu_fp_stdata_bits_uop_imm_packed; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_csr_addr = core_io_lsu_fp_stdata_bits_uop_csr_addr; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_rob_idx = core_io_lsu_fp_stdata_bits_uop_rob_idx; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_ldq_idx = core_io_lsu_fp_stdata_bits_uop_ldq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_stq_idx = core_io_lsu_fp_stdata_bits_uop_stq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_rxq_idx = core_io_lsu_fp_stdata_bits_uop_rxq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_pdst = core_io_lsu_fp_stdata_bits_uop_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_prs1 = core_io_lsu_fp_stdata_bits_uop_prs1; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_prs2 = core_io_lsu_fp_stdata_bits_uop_prs2; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_prs3 = core_io_lsu_fp_stdata_bits_uop_prs3; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_ppred = core_io_lsu_fp_stdata_bits_uop_ppred; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_prs1_busy = core_io_lsu_fp_stdata_bits_uop_prs1_busy; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_prs2_busy = core_io_lsu_fp_stdata_bits_uop_prs2_busy; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_prs3_busy = core_io_lsu_fp_stdata_bits_uop_prs3_busy; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_ppred_busy = core_io_lsu_fp_stdata_bits_uop_ppred_busy; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_stale_pdst = core_io_lsu_fp_stdata_bits_uop_stale_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_exception = core_io_lsu_fp_stdata_bits_uop_exception; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_exc_cause = core_io_lsu_fp_stdata_bits_uop_exc_cause; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_bypassable = core_io_lsu_fp_stdata_bits_uop_bypassable; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_mem_cmd = core_io_lsu_fp_stdata_bits_uop_mem_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_mem_size = core_io_lsu_fp_stdata_bits_uop_mem_size; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_mem_signed = core_io_lsu_fp_stdata_bits_uop_mem_signed; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_is_fence = core_io_lsu_fp_stdata_bits_uop_is_fence; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_is_fencei = core_io_lsu_fp_stdata_bits_uop_is_fencei; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_is_amo = core_io_lsu_fp_stdata_bits_uop_is_amo; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_uses_ldq = core_io_lsu_fp_stdata_bits_uop_uses_ldq; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_uses_stq = core_io_lsu_fp_stdata_bits_uop_uses_stq; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_is_sys_pc2epc = core_io_lsu_fp_stdata_bits_uop_is_sys_pc2epc; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_is_unique = core_io_lsu_fp_stdata_bits_uop_is_unique; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_flush_on_commit = core_io_lsu_fp_stdata_bits_uop_flush_on_commit; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_ldst_is_rs1 = core_io_lsu_fp_stdata_bits_uop_ldst_is_rs1; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_ldst = core_io_lsu_fp_stdata_bits_uop_ldst; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_lrs1 = core_io_lsu_fp_stdata_bits_uop_lrs1; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_lrs2 = core_io_lsu_fp_stdata_bits_uop_lrs2; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_lrs3 = core_io_lsu_fp_stdata_bits_uop_lrs3; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_ldst_val = core_io_lsu_fp_stdata_bits_uop_ldst_val; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_dst_rtype = core_io_lsu_fp_stdata_bits_uop_dst_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_lrs1_rtype = core_io_lsu_fp_stdata_bits_uop_lrs1_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_lrs2_rtype = core_io_lsu_fp_stdata_bits_uop_lrs2_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_frs3_en = core_io_lsu_fp_stdata_bits_uop_frs3_en; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_fp_val = core_io_lsu_fp_stdata_bits_uop_fp_val; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_fp_single = core_io_lsu_fp_stdata_bits_uop_fp_single; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_xcpt_pf_if = core_io_lsu_fp_stdata_bits_uop_xcpt_pf_if; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_xcpt_ae_if = core_io_lsu_fp_stdata_bits_uop_xcpt_ae_if; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_xcpt_ma_if = core_io_lsu_fp_stdata_bits_uop_xcpt_ma_if; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_bp_debug_if = core_io_lsu_fp_stdata_bits_uop_bp_debug_if; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_bp_xcpt_if = core_io_lsu_fp_stdata_bits_uop_bp_xcpt_if; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_debug_fsrc = core_io_lsu_fp_stdata_bits_uop_debug_fsrc; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_uop_debug_tsrc = core_io_lsu_fp_stdata_bits_uop_debug_tsrc; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_data = core_io_lsu_fp_stdata_bits_data; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_predicated = core_io_lsu_fp_stdata_bits_predicated; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_valid = core_io_lsu_fp_stdata_bits_fflags_valid; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_switch = core_io_lsu_fp_stdata_bits_fflags_bits_uop_switch; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_switch_off = core_io_lsu_fp_stdata_bits_fflags_bits_uop_switch_off; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_unicore = core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_unicore; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_shift = core_io_lsu_fp_stdata_bits_fflags_bits_uop_shift; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_lrs3_rtype = core_io_lsu_fp_stdata_bits_fflags_bits_uop_lrs3_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_rflag = core_io_lsu_fp_stdata_bits_fflags_bits_uop_rflag; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_wflag = core_io_lsu_fp_stdata_bits_fflags_bits_uop_wflag; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_prflag = core_io_lsu_fp_stdata_bits_fflags_bits_uop_prflag; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_pwflag = core_io_lsu_fp_stdata_bits_fflags_bits_uop_pwflag; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_pflag_busy = core_io_lsu_fp_stdata_bits_fflags_bits_uop_pflag_busy; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_stale_pflag = core_io_lsu_fp_stdata_bits_fflags_bits_uop_stale_pflag
    ; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_op1_sel = core_io_lsu_fp_stdata_bits_fflags_bits_uop_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_op2_sel = core_io_lsu_fp_stdata_bits_fflags_bits_uop_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_split_num = core_io_lsu_fp_stdata_bits_fflags_bits_uop_split_num; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_self_index = core_io_lsu_fp_stdata_bits_fflags_bits_uop_self_index; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_rob_inst_idx =
    core_io_lsu_fp_stdata_bits_fflags_bits_uop_rob_inst_idx; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_address_num = core_io_lsu_fp_stdata_bits_fflags_bits_uop_address_num
    ; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_uopc = core_io_lsu_fp_stdata_bits_fflags_bits_uop_uopc; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_inst = core_io_lsu_fp_stdata_bits_fflags_bits_uop_inst; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_debug_inst = core_io_lsu_fp_stdata_bits_fflags_bits_uop_debug_inst; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_rvc = core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_rvc; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_debug_pc = core_io_lsu_fp_stdata_bits_fflags_bits_uop_debug_pc; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_iq_type = core_io_lsu_fp_stdata_bits_fflags_bits_uop_iq_type; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_fu_code = core_io_lsu_fp_stdata_bits_fflags_bits_uop_fu_code; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_br_type =
    core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_br_type; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_op1_sel =
    core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_op2_sel =
    core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_imm_sel =
    core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_imm_sel; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_op_fcn = core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_op_fcn
    ; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_fcn_dw = core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_fcn_dw
    ; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_csr_cmd =
    core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_csr_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_is_load =
    core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_is_load; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_is_sta = core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_is_sta
    ; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_is_std = core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_is_std
    ; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_ctrl_op3_sel =
    core_io_lsu_fp_stdata_bits_fflags_bits_uop_ctrl_op3_sel; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_iw_state = core_io_lsu_fp_stdata_bits_fflags_bits_uop_iw_state; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_iw_p1_poisoned =
    core_io_lsu_fp_stdata_bits_fflags_bits_uop_iw_p1_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_iw_p2_poisoned =
    core_io_lsu_fp_stdata_bits_fflags_bits_uop_iw_p2_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_br = core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_br; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_jalr = core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_jalr; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_jal = core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_jal; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_sfb = core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_sfb; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_br_mask = core_io_lsu_fp_stdata_bits_fflags_bits_uop_br_mask; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_br_tag = core_io_lsu_fp_stdata_bits_fflags_bits_uop_br_tag; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_ftq_idx = core_io_lsu_fp_stdata_bits_fflags_bits_uop_ftq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_edge_inst = core_io_lsu_fp_stdata_bits_fflags_bits_uop_edge_inst; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_pc_lob = core_io_lsu_fp_stdata_bits_fflags_bits_uop_pc_lob; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_taken = core_io_lsu_fp_stdata_bits_fflags_bits_uop_taken; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_imm_packed = core_io_lsu_fp_stdata_bits_fflags_bits_uop_imm_packed; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_csr_addr = core_io_lsu_fp_stdata_bits_fflags_bits_uop_csr_addr; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_rob_idx = core_io_lsu_fp_stdata_bits_fflags_bits_uop_rob_idx; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_ldq_idx = core_io_lsu_fp_stdata_bits_fflags_bits_uop_ldq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_stq_idx = core_io_lsu_fp_stdata_bits_fflags_bits_uop_stq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_rxq_idx = core_io_lsu_fp_stdata_bits_fflags_bits_uop_rxq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_pdst = core_io_lsu_fp_stdata_bits_fflags_bits_uop_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_prs1 = core_io_lsu_fp_stdata_bits_fflags_bits_uop_prs1; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_prs2 = core_io_lsu_fp_stdata_bits_fflags_bits_uop_prs2; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_prs3 = core_io_lsu_fp_stdata_bits_fflags_bits_uop_prs3; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_ppred = core_io_lsu_fp_stdata_bits_fflags_bits_uop_ppred; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_prs1_busy = core_io_lsu_fp_stdata_bits_fflags_bits_uop_prs1_busy; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_prs2_busy = core_io_lsu_fp_stdata_bits_fflags_bits_uop_prs2_busy; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_prs3_busy = core_io_lsu_fp_stdata_bits_fflags_bits_uop_prs3_busy; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_ppred_busy = core_io_lsu_fp_stdata_bits_fflags_bits_uop_ppred_busy; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_stale_pdst = core_io_lsu_fp_stdata_bits_fflags_bits_uop_stale_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_exception = core_io_lsu_fp_stdata_bits_fflags_bits_uop_exception; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_exc_cause = core_io_lsu_fp_stdata_bits_fflags_bits_uop_exc_cause; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_bypassable = core_io_lsu_fp_stdata_bits_fflags_bits_uop_bypassable; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_mem_cmd = core_io_lsu_fp_stdata_bits_fflags_bits_uop_mem_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_mem_size = core_io_lsu_fp_stdata_bits_fflags_bits_uop_mem_size; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_mem_signed = core_io_lsu_fp_stdata_bits_fflags_bits_uop_mem_signed; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_fence = core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_fence; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_fencei = core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_fencei; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_amo = core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_amo; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_uses_ldq = core_io_lsu_fp_stdata_bits_fflags_bits_uop_uses_ldq; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_uses_stq = core_io_lsu_fp_stdata_bits_fflags_bits_uop_uses_stq; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_sys_pc2epc =
    core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_sys_pc2epc; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_is_unique = core_io_lsu_fp_stdata_bits_fflags_bits_uop_is_unique; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_flush_on_commit =
    core_io_lsu_fp_stdata_bits_fflags_bits_uop_flush_on_commit; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_ldst_is_rs1 = core_io_lsu_fp_stdata_bits_fflags_bits_uop_ldst_is_rs1
    ; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_ldst = core_io_lsu_fp_stdata_bits_fflags_bits_uop_ldst; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_lrs1 = core_io_lsu_fp_stdata_bits_fflags_bits_uop_lrs1; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_lrs2 = core_io_lsu_fp_stdata_bits_fflags_bits_uop_lrs2; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_lrs3 = core_io_lsu_fp_stdata_bits_fflags_bits_uop_lrs3; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_ldst_val = core_io_lsu_fp_stdata_bits_fflags_bits_uop_ldst_val; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_dst_rtype = core_io_lsu_fp_stdata_bits_fflags_bits_uop_dst_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_lrs1_rtype = core_io_lsu_fp_stdata_bits_fflags_bits_uop_lrs1_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_lrs2_rtype = core_io_lsu_fp_stdata_bits_fflags_bits_uop_lrs2_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_frs3_en = core_io_lsu_fp_stdata_bits_fflags_bits_uop_frs3_en; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_fp_val = core_io_lsu_fp_stdata_bits_fflags_bits_uop_fp_val; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_fp_single = core_io_lsu_fp_stdata_bits_fflags_bits_uop_fp_single; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_xcpt_pf_if = core_io_lsu_fp_stdata_bits_fflags_bits_uop_xcpt_pf_if; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_xcpt_ae_if = core_io_lsu_fp_stdata_bits_fflags_bits_uop_xcpt_ae_if; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_xcpt_ma_if = core_io_lsu_fp_stdata_bits_fflags_bits_uop_xcpt_ma_if; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_bp_debug_if = core_io_lsu_fp_stdata_bits_fflags_bits_uop_bp_debug_if
    ; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_bp_xcpt_if = core_io_lsu_fp_stdata_bits_fflags_bits_uop_bp_xcpt_if; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_debug_fsrc = core_io_lsu_fp_stdata_bits_fflags_bits_uop_debug_fsrc; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_uop_debug_tsrc = core_io_lsu_fp_stdata_bits_fflags_bits_uop_debug_tsrc; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflags_bits_flags = core_io_lsu_fp_stdata_bits_fflags_bits_flags; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_flagdata = core_io_lsu_fp_stdata_bits_flagdata; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_valid = core_io_lsu_fp_stdata_bits_fflagdata_valid; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_switch = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_switch; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_switch_off =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_switch_off; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_unicore =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_unicore; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_shift = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_shift; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_lrs3_rtype =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs3_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_rflag = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_rflag; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_wflag = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_wflag; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_prflag = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_prflag; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_pwflag = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_pwflag; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_pflag_busy =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_pflag_busy; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_stale_pflag =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_stale_pflag; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_op1_sel = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_op2_sel = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_split_num =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_split_num; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_self_index =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_self_index; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_rob_inst_idx =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_rob_inst_idx; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_address_num =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_address_num; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_uopc = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_uopc; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_inst = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_inst; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_debug_inst =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_debug_inst; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_rvc = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_rvc; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_debug_pc = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_debug_pc
    ; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_iq_type = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_iq_type; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_fu_code = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_fu_code; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_br_type =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_br_type; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_op1_sel =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_op2_sel =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_imm_sel =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_imm_sel; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_op_fcn =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_op_fcn; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_fcn_dw =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_fcn_dw; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_csr_cmd =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_csr_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_load =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_load; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_sta =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_sta; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_std =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_is_std; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ctrl_op3_sel =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ctrl_op3_sel; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_iw_state = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_iw_state
    ; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_iw_p1_poisoned =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_iw_p1_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_iw_p2_poisoned =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_iw_p2_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_br = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_br; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_jalr = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_jalr; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_jal = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_jal; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_sfb = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_sfb; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_br_mask = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_br_mask; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_br_tag = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_br_tag; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ftq_idx = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ftq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_edge_inst =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_edge_inst; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_pc_lob = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_pc_lob; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_taken = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_taken; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_imm_packed =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_imm_packed; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_csr_addr = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_csr_addr
    ; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_rob_idx = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_rob_idx; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ldq_idx = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ldq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_stq_idx = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_stq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_rxq_idx = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_rxq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_pdst = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_prs1 = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs1; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_prs2 = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs2; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_prs3 = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs3; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ppred = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ppred; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_prs1_busy =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs1_busy; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_prs2_busy =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs2_busy; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_prs3_busy =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_prs3_busy; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ppred_busy =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ppred_busy; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_stale_pdst =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_stale_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_exception =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_exception; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_exc_cause =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_exc_cause; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_bypassable =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_bypassable; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_mem_cmd = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_mem_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_mem_size = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_mem_size
    ; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_mem_signed =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_mem_signed; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_fence = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_fence
    ; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_fencei =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_fencei; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_amo = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_amo; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_uses_ldq = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_uses_ldq
    ; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_uses_stq = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_uses_stq
    ; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_sys_pc2epc =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_sys_pc2epc; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_is_unique =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_is_unique; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_flush_on_commit =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_flush_on_commit; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ldst_is_rs1 =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ldst_is_rs1; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ldst = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ldst; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_lrs1 = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs1; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_lrs2 = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs2; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_lrs3 = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs3; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_ldst_val = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_ldst_val
    ; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_dst_rtype =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_dst_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_lrs1_rtype =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs1_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_lrs2_rtype =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_lrs2_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_frs3_en = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_frs3_en; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_fp_val = core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_fp_val; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_fp_single =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_fp_single; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_xcpt_pf_if =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_xcpt_pf_if; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_xcpt_ae_if =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_xcpt_ae_if; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_xcpt_ma_if =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_xcpt_ma_if; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_bp_debug_if =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_bp_debug_if; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_bp_xcpt_if =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_bp_xcpt_if; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_debug_fsrc =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_debug_fsrc; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_uop_debug_tsrc =
    core_io_lsu_fp_stdata_bits_fflagdata_bits_uop_debug_tsrc; // @[tile.scala 178:15]
  assign lsu_io_core_fp_stdata_bits_fflagdata_bits_fflag = core_io_lsu_fp_stdata_bits_fflagdata_bits_fflag; // @[tile.scala 178:15]
  assign lsu_io_core_commit_valids_0 = core_io_lsu_commit_valids_0; // @[tile.scala 178:15]
  assign lsu_io_core_commit_valids_1 = core_io_lsu_commit_valids_1; // @[tile.scala 178:15]
  assign lsu_io_core_commit_arch_valids_0 = core_io_lsu_commit_arch_valids_0; // @[tile.scala 178:15]
  assign lsu_io_core_commit_arch_valids_1 = core_io_lsu_commit_arch_valids_1; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_switch = core_io_lsu_commit_uops_0_switch; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_switch_off = core_io_lsu_commit_uops_0_switch_off; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_is_unicore = core_io_lsu_commit_uops_0_is_unicore; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_shift = core_io_lsu_commit_uops_0_shift; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_lrs3_rtype = core_io_lsu_commit_uops_0_lrs3_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_rflag = core_io_lsu_commit_uops_0_rflag; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_wflag = core_io_lsu_commit_uops_0_wflag; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_prflag = core_io_lsu_commit_uops_0_prflag; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_pwflag = core_io_lsu_commit_uops_0_pwflag; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_pflag_busy = core_io_lsu_commit_uops_0_pflag_busy; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_stale_pflag = core_io_lsu_commit_uops_0_stale_pflag; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_op1_sel = core_io_lsu_commit_uops_0_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_op2_sel = core_io_lsu_commit_uops_0_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_split_num = core_io_lsu_commit_uops_0_split_num; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_self_index = core_io_lsu_commit_uops_0_self_index; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_rob_inst_idx = core_io_lsu_commit_uops_0_rob_inst_idx; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_address_num = core_io_lsu_commit_uops_0_address_num; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_uopc = core_io_lsu_commit_uops_0_uopc; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_inst = core_io_lsu_commit_uops_0_inst; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_debug_inst = core_io_lsu_commit_uops_0_debug_inst; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_is_rvc = core_io_lsu_commit_uops_0_is_rvc; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_debug_pc = core_io_lsu_commit_uops_0_debug_pc; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_iq_type = core_io_lsu_commit_uops_0_iq_type; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_fu_code = core_io_lsu_commit_uops_0_fu_code; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_ctrl_br_type = core_io_lsu_commit_uops_0_ctrl_br_type; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_ctrl_op1_sel = core_io_lsu_commit_uops_0_ctrl_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_ctrl_op2_sel = core_io_lsu_commit_uops_0_ctrl_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_ctrl_imm_sel = core_io_lsu_commit_uops_0_ctrl_imm_sel; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_ctrl_op_fcn = core_io_lsu_commit_uops_0_ctrl_op_fcn; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_ctrl_fcn_dw = core_io_lsu_commit_uops_0_ctrl_fcn_dw; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_ctrl_csr_cmd = core_io_lsu_commit_uops_0_ctrl_csr_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_ctrl_is_load = core_io_lsu_commit_uops_0_ctrl_is_load; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_ctrl_is_sta = core_io_lsu_commit_uops_0_ctrl_is_sta; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_ctrl_is_std = core_io_lsu_commit_uops_0_ctrl_is_std; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_ctrl_op3_sel = core_io_lsu_commit_uops_0_ctrl_op3_sel; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_iw_state = core_io_lsu_commit_uops_0_iw_state; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_iw_p1_poisoned = core_io_lsu_commit_uops_0_iw_p1_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_iw_p2_poisoned = core_io_lsu_commit_uops_0_iw_p2_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_is_br = core_io_lsu_commit_uops_0_is_br; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_is_jalr = core_io_lsu_commit_uops_0_is_jalr; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_is_jal = core_io_lsu_commit_uops_0_is_jal; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_is_sfb = core_io_lsu_commit_uops_0_is_sfb; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_br_mask = core_io_lsu_commit_uops_0_br_mask; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_br_tag = core_io_lsu_commit_uops_0_br_tag; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_ftq_idx = core_io_lsu_commit_uops_0_ftq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_edge_inst = core_io_lsu_commit_uops_0_edge_inst; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_pc_lob = core_io_lsu_commit_uops_0_pc_lob; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_taken = core_io_lsu_commit_uops_0_taken; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_imm_packed = core_io_lsu_commit_uops_0_imm_packed; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_csr_addr = core_io_lsu_commit_uops_0_csr_addr; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_rob_idx = core_io_lsu_commit_uops_0_rob_idx; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_ldq_idx = core_io_lsu_commit_uops_0_ldq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_stq_idx = core_io_lsu_commit_uops_0_stq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_rxq_idx = core_io_lsu_commit_uops_0_rxq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_pdst = core_io_lsu_commit_uops_0_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_prs1 = core_io_lsu_commit_uops_0_prs1; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_prs2 = core_io_lsu_commit_uops_0_prs2; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_prs3 = core_io_lsu_commit_uops_0_prs3; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_ppred = core_io_lsu_commit_uops_0_ppred; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_prs1_busy = core_io_lsu_commit_uops_0_prs1_busy; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_prs2_busy = core_io_lsu_commit_uops_0_prs2_busy; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_prs3_busy = core_io_lsu_commit_uops_0_prs3_busy; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_ppred_busy = core_io_lsu_commit_uops_0_ppred_busy; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_stale_pdst = core_io_lsu_commit_uops_0_stale_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_exception = core_io_lsu_commit_uops_0_exception; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_exc_cause = core_io_lsu_commit_uops_0_exc_cause; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_bypassable = core_io_lsu_commit_uops_0_bypassable; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_mem_cmd = core_io_lsu_commit_uops_0_mem_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_mem_size = core_io_lsu_commit_uops_0_mem_size; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_mem_signed = core_io_lsu_commit_uops_0_mem_signed; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_is_fence = core_io_lsu_commit_uops_0_is_fence; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_is_fencei = core_io_lsu_commit_uops_0_is_fencei; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_is_amo = core_io_lsu_commit_uops_0_is_amo; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_uses_ldq = core_io_lsu_commit_uops_0_uses_ldq; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_uses_stq = core_io_lsu_commit_uops_0_uses_stq; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_is_sys_pc2epc = core_io_lsu_commit_uops_0_is_sys_pc2epc; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_is_unique = core_io_lsu_commit_uops_0_is_unique; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_flush_on_commit = core_io_lsu_commit_uops_0_flush_on_commit; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_ldst_is_rs1 = core_io_lsu_commit_uops_0_ldst_is_rs1; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_ldst = core_io_lsu_commit_uops_0_ldst; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_lrs1 = core_io_lsu_commit_uops_0_lrs1; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_lrs2 = core_io_lsu_commit_uops_0_lrs2; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_lrs3 = core_io_lsu_commit_uops_0_lrs3; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_ldst_val = core_io_lsu_commit_uops_0_ldst_val; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_dst_rtype = core_io_lsu_commit_uops_0_dst_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_lrs1_rtype = core_io_lsu_commit_uops_0_lrs1_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_lrs2_rtype = core_io_lsu_commit_uops_0_lrs2_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_frs3_en = core_io_lsu_commit_uops_0_frs3_en; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_fp_val = core_io_lsu_commit_uops_0_fp_val; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_fp_single = core_io_lsu_commit_uops_0_fp_single; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_xcpt_pf_if = core_io_lsu_commit_uops_0_xcpt_pf_if; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_xcpt_ae_if = core_io_lsu_commit_uops_0_xcpt_ae_if; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_xcpt_ma_if = core_io_lsu_commit_uops_0_xcpt_ma_if; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_bp_debug_if = core_io_lsu_commit_uops_0_bp_debug_if; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_bp_xcpt_if = core_io_lsu_commit_uops_0_bp_xcpt_if; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_debug_fsrc = core_io_lsu_commit_uops_0_debug_fsrc; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_0_debug_tsrc = core_io_lsu_commit_uops_0_debug_tsrc; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_switch = core_io_lsu_commit_uops_1_switch; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_switch_off = core_io_lsu_commit_uops_1_switch_off; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_is_unicore = core_io_lsu_commit_uops_1_is_unicore; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_shift = core_io_lsu_commit_uops_1_shift; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_lrs3_rtype = core_io_lsu_commit_uops_1_lrs3_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_rflag = core_io_lsu_commit_uops_1_rflag; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_wflag = core_io_lsu_commit_uops_1_wflag; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_prflag = core_io_lsu_commit_uops_1_prflag; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_pwflag = core_io_lsu_commit_uops_1_pwflag; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_pflag_busy = core_io_lsu_commit_uops_1_pflag_busy; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_stale_pflag = core_io_lsu_commit_uops_1_stale_pflag; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_op1_sel = core_io_lsu_commit_uops_1_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_op2_sel = core_io_lsu_commit_uops_1_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_split_num = core_io_lsu_commit_uops_1_split_num; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_self_index = core_io_lsu_commit_uops_1_self_index; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_rob_inst_idx = core_io_lsu_commit_uops_1_rob_inst_idx; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_address_num = core_io_lsu_commit_uops_1_address_num; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_uopc = core_io_lsu_commit_uops_1_uopc; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_inst = core_io_lsu_commit_uops_1_inst; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_debug_inst = core_io_lsu_commit_uops_1_debug_inst; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_is_rvc = core_io_lsu_commit_uops_1_is_rvc; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_debug_pc = core_io_lsu_commit_uops_1_debug_pc; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_iq_type = core_io_lsu_commit_uops_1_iq_type; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_fu_code = core_io_lsu_commit_uops_1_fu_code; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_ctrl_br_type = core_io_lsu_commit_uops_1_ctrl_br_type; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_ctrl_op1_sel = core_io_lsu_commit_uops_1_ctrl_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_ctrl_op2_sel = core_io_lsu_commit_uops_1_ctrl_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_ctrl_imm_sel = core_io_lsu_commit_uops_1_ctrl_imm_sel; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_ctrl_op_fcn = core_io_lsu_commit_uops_1_ctrl_op_fcn; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_ctrl_fcn_dw = core_io_lsu_commit_uops_1_ctrl_fcn_dw; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_ctrl_csr_cmd = core_io_lsu_commit_uops_1_ctrl_csr_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_ctrl_is_load = core_io_lsu_commit_uops_1_ctrl_is_load; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_ctrl_is_sta = core_io_lsu_commit_uops_1_ctrl_is_sta; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_ctrl_is_std = core_io_lsu_commit_uops_1_ctrl_is_std; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_ctrl_op3_sel = core_io_lsu_commit_uops_1_ctrl_op3_sel; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_iw_state = core_io_lsu_commit_uops_1_iw_state; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_iw_p1_poisoned = core_io_lsu_commit_uops_1_iw_p1_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_iw_p2_poisoned = core_io_lsu_commit_uops_1_iw_p2_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_is_br = core_io_lsu_commit_uops_1_is_br; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_is_jalr = core_io_lsu_commit_uops_1_is_jalr; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_is_jal = core_io_lsu_commit_uops_1_is_jal; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_is_sfb = core_io_lsu_commit_uops_1_is_sfb; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_br_mask = core_io_lsu_commit_uops_1_br_mask; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_br_tag = core_io_lsu_commit_uops_1_br_tag; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_ftq_idx = core_io_lsu_commit_uops_1_ftq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_edge_inst = core_io_lsu_commit_uops_1_edge_inst; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_pc_lob = core_io_lsu_commit_uops_1_pc_lob; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_taken = core_io_lsu_commit_uops_1_taken; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_imm_packed = core_io_lsu_commit_uops_1_imm_packed; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_csr_addr = core_io_lsu_commit_uops_1_csr_addr; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_rob_idx = core_io_lsu_commit_uops_1_rob_idx; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_ldq_idx = core_io_lsu_commit_uops_1_ldq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_stq_idx = core_io_lsu_commit_uops_1_stq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_rxq_idx = core_io_lsu_commit_uops_1_rxq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_pdst = core_io_lsu_commit_uops_1_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_prs1 = core_io_lsu_commit_uops_1_prs1; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_prs2 = core_io_lsu_commit_uops_1_prs2; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_prs3 = core_io_lsu_commit_uops_1_prs3; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_ppred = core_io_lsu_commit_uops_1_ppred; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_prs1_busy = core_io_lsu_commit_uops_1_prs1_busy; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_prs2_busy = core_io_lsu_commit_uops_1_prs2_busy; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_prs3_busy = core_io_lsu_commit_uops_1_prs3_busy; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_ppred_busy = core_io_lsu_commit_uops_1_ppred_busy; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_stale_pdst = core_io_lsu_commit_uops_1_stale_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_exception = core_io_lsu_commit_uops_1_exception; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_exc_cause = core_io_lsu_commit_uops_1_exc_cause; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_bypassable = core_io_lsu_commit_uops_1_bypassable; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_mem_cmd = core_io_lsu_commit_uops_1_mem_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_mem_size = core_io_lsu_commit_uops_1_mem_size; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_mem_signed = core_io_lsu_commit_uops_1_mem_signed; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_is_fence = core_io_lsu_commit_uops_1_is_fence; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_is_fencei = core_io_lsu_commit_uops_1_is_fencei; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_is_amo = core_io_lsu_commit_uops_1_is_amo; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_uses_ldq = core_io_lsu_commit_uops_1_uses_ldq; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_uses_stq = core_io_lsu_commit_uops_1_uses_stq; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_is_sys_pc2epc = core_io_lsu_commit_uops_1_is_sys_pc2epc; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_is_unique = core_io_lsu_commit_uops_1_is_unique; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_flush_on_commit = core_io_lsu_commit_uops_1_flush_on_commit; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_ldst_is_rs1 = core_io_lsu_commit_uops_1_ldst_is_rs1; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_ldst = core_io_lsu_commit_uops_1_ldst; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_lrs1 = core_io_lsu_commit_uops_1_lrs1; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_lrs2 = core_io_lsu_commit_uops_1_lrs2; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_lrs3 = core_io_lsu_commit_uops_1_lrs3; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_ldst_val = core_io_lsu_commit_uops_1_ldst_val; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_dst_rtype = core_io_lsu_commit_uops_1_dst_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_lrs1_rtype = core_io_lsu_commit_uops_1_lrs1_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_lrs2_rtype = core_io_lsu_commit_uops_1_lrs2_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_frs3_en = core_io_lsu_commit_uops_1_frs3_en; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_fp_val = core_io_lsu_commit_uops_1_fp_val; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_fp_single = core_io_lsu_commit_uops_1_fp_single; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_xcpt_pf_if = core_io_lsu_commit_uops_1_xcpt_pf_if; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_xcpt_ae_if = core_io_lsu_commit_uops_1_xcpt_ae_if; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_xcpt_ma_if = core_io_lsu_commit_uops_1_xcpt_ma_if; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_bp_debug_if = core_io_lsu_commit_uops_1_bp_debug_if; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_bp_xcpt_if = core_io_lsu_commit_uops_1_bp_xcpt_if; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_debug_fsrc = core_io_lsu_commit_uops_1_debug_fsrc; // @[tile.scala 178:15]
  assign lsu_io_core_commit_uops_1_debug_tsrc = core_io_lsu_commit_uops_1_debug_tsrc; // @[tile.scala 178:15]
  assign lsu_io_core_commit_fflags_valid = core_io_lsu_commit_fflags_valid; // @[tile.scala 178:15]
  assign lsu_io_core_commit_fflags_bits = core_io_lsu_commit_fflags_bits; // @[tile.scala 178:15]
  assign lsu_io_core_commit_fflag_exception_valid = core_io_lsu_commit_fflag_exception_valid; // @[tile.scala 178:15]
  assign lsu_io_core_commit_fflag_exception_bits = core_io_lsu_commit_fflag_exception_bits; // @[tile.scala 178:15]
  assign lsu_io_core_commit_debug_insts_0 = core_io_lsu_commit_debug_insts_0; // @[tile.scala 178:15]
  assign lsu_io_core_commit_debug_insts_1 = core_io_lsu_commit_debug_insts_1; // @[tile.scala 178:15]
  assign lsu_io_core_commit_rbk_valids_0 = core_io_lsu_commit_rbk_valids_0; // @[tile.scala 178:15]
  assign lsu_io_core_commit_rbk_valids_1 = core_io_lsu_commit_rbk_valids_1; // @[tile.scala 178:15]
  assign lsu_io_core_commit_rollback = core_io_lsu_commit_rollback; // @[tile.scala 178:15]
  assign lsu_io_core_commit_debug_wdata_0 = core_io_lsu_commit_debug_wdata_0; // @[tile.scala 178:15]
  assign lsu_io_core_commit_debug_wdata_1 = core_io_lsu_commit_debug_wdata_1; // @[tile.scala 178:15]
  assign lsu_io_core_commit_debug_wflagdata_0 = core_io_lsu_commit_debug_wflagdata_0; // @[tile.scala 178:15]
  assign lsu_io_core_commit_debug_wflagdata_1 = core_io_lsu_commit_debug_wflagdata_1; // @[tile.scala 178:15]
  assign lsu_io_core_commit_load_at_rob_head = core_io_lsu_commit_load_at_rob_head; // @[tile.scala 178:15]
  assign lsu_io_core_fence_dmem = core_io_lsu_fence_dmem; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b1_resolve_mask = core_io_lsu_brupdate_b1_resolve_mask; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b1_mispredict_mask = core_io_lsu_brupdate_b1_mispredict_mask; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_switch = core_io_lsu_brupdate_b2_uop_switch; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_switch_off = core_io_lsu_brupdate_b2_uop_switch_off; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_is_unicore = core_io_lsu_brupdate_b2_uop_is_unicore; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_shift = core_io_lsu_brupdate_b2_uop_shift; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_lrs3_rtype = core_io_lsu_brupdate_b2_uop_lrs3_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_rflag = core_io_lsu_brupdate_b2_uop_rflag; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_wflag = core_io_lsu_brupdate_b2_uop_wflag; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_prflag = core_io_lsu_brupdate_b2_uop_prflag; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_pwflag = core_io_lsu_brupdate_b2_uop_pwflag; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_pflag_busy = core_io_lsu_brupdate_b2_uop_pflag_busy; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_stale_pflag = core_io_lsu_brupdate_b2_uop_stale_pflag; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_op1_sel = core_io_lsu_brupdate_b2_uop_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_op2_sel = core_io_lsu_brupdate_b2_uop_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_split_num = core_io_lsu_brupdate_b2_uop_split_num; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_self_index = core_io_lsu_brupdate_b2_uop_self_index; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_rob_inst_idx = core_io_lsu_brupdate_b2_uop_rob_inst_idx; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_address_num = core_io_lsu_brupdate_b2_uop_address_num; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_uopc = core_io_lsu_brupdate_b2_uop_uopc; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_inst = core_io_lsu_brupdate_b2_uop_inst; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_debug_inst = core_io_lsu_brupdate_b2_uop_debug_inst; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_is_rvc = core_io_lsu_brupdate_b2_uop_is_rvc; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_debug_pc = core_io_lsu_brupdate_b2_uop_debug_pc; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_iq_type = core_io_lsu_brupdate_b2_uop_iq_type; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_fu_code = core_io_lsu_brupdate_b2_uop_fu_code; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_ctrl_br_type = core_io_lsu_brupdate_b2_uop_ctrl_br_type; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_ctrl_op1_sel = core_io_lsu_brupdate_b2_uop_ctrl_op1_sel; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_ctrl_op2_sel = core_io_lsu_brupdate_b2_uop_ctrl_op2_sel; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_ctrl_imm_sel = core_io_lsu_brupdate_b2_uop_ctrl_imm_sel; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_ctrl_op_fcn = core_io_lsu_brupdate_b2_uop_ctrl_op_fcn; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_ctrl_fcn_dw = core_io_lsu_brupdate_b2_uop_ctrl_fcn_dw; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_ctrl_csr_cmd = core_io_lsu_brupdate_b2_uop_ctrl_csr_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_ctrl_is_load = core_io_lsu_brupdate_b2_uop_ctrl_is_load; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_ctrl_is_sta = core_io_lsu_brupdate_b2_uop_ctrl_is_sta; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_ctrl_is_std = core_io_lsu_brupdate_b2_uop_ctrl_is_std; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_ctrl_op3_sel = core_io_lsu_brupdate_b2_uop_ctrl_op3_sel; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_iw_state = core_io_lsu_brupdate_b2_uop_iw_state; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_iw_p1_poisoned = core_io_lsu_brupdate_b2_uop_iw_p1_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_iw_p2_poisoned = core_io_lsu_brupdate_b2_uop_iw_p2_poisoned; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_is_br = core_io_lsu_brupdate_b2_uop_is_br; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_is_jalr = core_io_lsu_brupdate_b2_uop_is_jalr; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_is_jal = core_io_lsu_brupdate_b2_uop_is_jal; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_is_sfb = core_io_lsu_brupdate_b2_uop_is_sfb; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_br_mask = core_io_lsu_brupdate_b2_uop_br_mask; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_br_tag = core_io_lsu_brupdate_b2_uop_br_tag; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_ftq_idx = core_io_lsu_brupdate_b2_uop_ftq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_edge_inst = core_io_lsu_brupdate_b2_uop_edge_inst; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_pc_lob = core_io_lsu_brupdate_b2_uop_pc_lob; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_taken = core_io_lsu_brupdate_b2_uop_taken; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_imm_packed = core_io_lsu_brupdate_b2_uop_imm_packed; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_csr_addr = core_io_lsu_brupdate_b2_uop_csr_addr; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_rob_idx = core_io_lsu_brupdate_b2_uop_rob_idx; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_ldq_idx = core_io_lsu_brupdate_b2_uop_ldq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_stq_idx = core_io_lsu_brupdate_b2_uop_stq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_rxq_idx = core_io_lsu_brupdate_b2_uop_rxq_idx; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_pdst = core_io_lsu_brupdate_b2_uop_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_prs1 = core_io_lsu_brupdate_b2_uop_prs1; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_prs2 = core_io_lsu_brupdate_b2_uop_prs2; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_prs3 = core_io_lsu_brupdate_b2_uop_prs3; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_ppred = core_io_lsu_brupdate_b2_uop_ppred; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_prs1_busy = core_io_lsu_brupdate_b2_uop_prs1_busy; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_prs2_busy = core_io_lsu_brupdate_b2_uop_prs2_busy; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_prs3_busy = core_io_lsu_brupdate_b2_uop_prs3_busy; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_ppred_busy = core_io_lsu_brupdate_b2_uop_ppred_busy; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_stale_pdst = core_io_lsu_brupdate_b2_uop_stale_pdst; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_exception = core_io_lsu_brupdate_b2_uop_exception; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_exc_cause = core_io_lsu_brupdate_b2_uop_exc_cause; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_bypassable = core_io_lsu_brupdate_b2_uop_bypassable; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_mem_cmd = core_io_lsu_brupdate_b2_uop_mem_cmd; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_mem_size = core_io_lsu_brupdate_b2_uop_mem_size; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_mem_signed = core_io_lsu_brupdate_b2_uop_mem_signed; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_is_fence = core_io_lsu_brupdate_b2_uop_is_fence; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_is_fencei = core_io_lsu_brupdate_b2_uop_is_fencei; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_is_amo = core_io_lsu_brupdate_b2_uop_is_amo; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_uses_ldq = core_io_lsu_brupdate_b2_uop_uses_ldq; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_uses_stq = core_io_lsu_brupdate_b2_uop_uses_stq; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_is_sys_pc2epc = core_io_lsu_brupdate_b2_uop_is_sys_pc2epc; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_is_unique = core_io_lsu_brupdate_b2_uop_is_unique; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_flush_on_commit = core_io_lsu_brupdate_b2_uop_flush_on_commit; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_ldst_is_rs1 = core_io_lsu_brupdate_b2_uop_ldst_is_rs1; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_ldst = core_io_lsu_brupdate_b2_uop_ldst; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_lrs1 = core_io_lsu_brupdate_b2_uop_lrs1; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_lrs2 = core_io_lsu_brupdate_b2_uop_lrs2; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_lrs3 = core_io_lsu_brupdate_b2_uop_lrs3; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_ldst_val = core_io_lsu_brupdate_b2_uop_ldst_val; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_dst_rtype = core_io_lsu_brupdate_b2_uop_dst_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_lrs1_rtype = core_io_lsu_brupdate_b2_uop_lrs1_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_lrs2_rtype = core_io_lsu_brupdate_b2_uop_lrs2_rtype; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_frs3_en = core_io_lsu_brupdate_b2_uop_frs3_en; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_fp_val = core_io_lsu_brupdate_b2_uop_fp_val; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_fp_single = core_io_lsu_brupdate_b2_uop_fp_single; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_xcpt_pf_if = core_io_lsu_brupdate_b2_uop_xcpt_pf_if; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_xcpt_ae_if = core_io_lsu_brupdate_b2_uop_xcpt_ae_if; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_xcpt_ma_if = core_io_lsu_brupdate_b2_uop_xcpt_ma_if; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_bp_debug_if = core_io_lsu_brupdate_b2_uop_bp_debug_if; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_bp_xcpt_if = core_io_lsu_brupdate_b2_uop_bp_xcpt_if; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_debug_fsrc = core_io_lsu_brupdate_b2_uop_debug_fsrc; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_uop_debug_tsrc = core_io_lsu_brupdate_b2_uop_debug_tsrc; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_valid = core_io_lsu_brupdate_b2_valid; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_mispredict = core_io_lsu_brupdate_b2_mispredict; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_taken = core_io_lsu_brupdate_b2_taken; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_cfi_type = core_io_lsu_brupdate_b2_cfi_type; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_pc_sel = core_io_lsu_brupdate_b2_pc_sel; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_jalr_target = core_io_lsu_brupdate_b2_jalr_target; // @[tile.scala 178:15]
  assign lsu_io_core_brupdate_b2_target_offset = core_io_lsu_brupdate_b2_target_offset; // @[tile.scala 178:15]
  assign lsu_io_core_rob_pnr_idx = core_io_lsu_rob_pnr_idx; // @[tile.scala 178:15]
  assign lsu_io_core_rob_head_idx = core_io_lsu_rob_head_idx; // @[tile.scala 178:15]
  assign lsu_io_core_exception = core_io_lsu_exception; // @[tile.scala 178:15]
  assign lsu_io_core_tsc_reg = core_io_lsu_tsc_reg; // @[tile.scala 178:15]
  assign lsu_io_dmem_req_ready = dcache_io_lsu_req_ready; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_valid = dcache_io_lsu_resp_0_valid; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_switch = dcache_io_lsu_resp_0_bits_uop_switch; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_switch_off = dcache_io_lsu_resp_0_bits_uop_switch_off; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_is_unicore = dcache_io_lsu_resp_0_bits_uop_is_unicore; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_shift = dcache_io_lsu_resp_0_bits_uop_shift; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_lrs3_rtype = dcache_io_lsu_resp_0_bits_uop_lrs3_rtype; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_rflag = dcache_io_lsu_resp_0_bits_uop_rflag; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_wflag = dcache_io_lsu_resp_0_bits_uop_wflag; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_prflag = dcache_io_lsu_resp_0_bits_uop_prflag; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_pwflag = dcache_io_lsu_resp_0_bits_uop_pwflag; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_pflag_busy = dcache_io_lsu_resp_0_bits_uop_pflag_busy; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_stale_pflag = dcache_io_lsu_resp_0_bits_uop_stale_pflag; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_op1_sel = dcache_io_lsu_resp_0_bits_uop_op1_sel; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_op2_sel = dcache_io_lsu_resp_0_bits_uop_op2_sel; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_split_num = dcache_io_lsu_resp_0_bits_uop_split_num; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_self_index = dcache_io_lsu_resp_0_bits_uop_self_index; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_rob_inst_idx = dcache_io_lsu_resp_0_bits_uop_rob_inst_idx; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_address_num = dcache_io_lsu_resp_0_bits_uop_address_num; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_uopc = dcache_io_lsu_resp_0_bits_uop_uopc; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_inst = dcache_io_lsu_resp_0_bits_uop_inst; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_debug_inst = dcache_io_lsu_resp_0_bits_uop_debug_inst; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_is_rvc = dcache_io_lsu_resp_0_bits_uop_is_rvc; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_debug_pc = dcache_io_lsu_resp_0_bits_uop_debug_pc; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_iq_type = dcache_io_lsu_resp_0_bits_uop_iq_type; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_fu_code = dcache_io_lsu_resp_0_bits_uop_fu_code; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_ctrl_br_type = dcache_io_lsu_resp_0_bits_uop_ctrl_br_type; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_ctrl_op1_sel = dcache_io_lsu_resp_0_bits_uop_ctrl_op1_sel; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_ctrl_op2_sel = dcache_io_lsu_resp_0_bits_uop_ctrl_op2_sel; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_ctrl_imm_sel = dcache_io_lsu_resp_0_bits_uop_ctrl_imm_sel; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_ctrl_op_fcn = dcache_io_lsu_resp_0_bits_uop_ctrl_op_fcn; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_ctrl_fcn_dw = dcache_io_lsu_resp_0_bits_uop_ctrl_fcn_dw; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_ctrl_csr_cmd = dcache_io_lsu_resp_0_bits_uop_ctrl_csr_cmd; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_ctrl_is_load = dcache_io_lsu_resp_0_bits_uop_ctrl_is_load; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_ctrl_is_sta = dcache_io_lsu_resp_0_bits_uop_ctrl_is_sta; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_ctrl_is_std = dcache_io_lsu_resp_0_bits_uop_ctrl_is_std; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_ctrl_op3_sel = dcache_io_lsu_resp_0_bits_uop_ctrl_op3_sel; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_iw_state = dcache_io_lsu_resp_0_bits_uop_iw_state; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_iw_p1_poisoned = dcache_io_lsu_resp_0_bits_uop_iw_p1_poisoned; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_iw_p2_poisoned = dcache_io_lsu_resp_0_bits_uop_iw_p2_poisoned; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_is_br = dcache_io_lsu_resp_0_bits_uop_is_br; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_is_jalr = dcache_io_lsu_resp_0_bits_uop_is_jalr; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_is_jal = dcache_io_lsu_resp_0_bits_uop_is_jal; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_is_sfb = dcache_io_lsu_resp_0_bits_uop_is_sfb; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_br_mask = dcache_io_lsu_resp_0_bits_uop_br_mask; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_br_tag = dcache_io_lsu_resp_0_bits_uop_br_tag; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_ftq_idx = dcache_io_lsu_resp_0_bits_uop_ftq_idx; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_edge_inst = dcache_io_lsu_resp_0_bits_uop_edge_inst; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_pc_lob = dcache_io_lsu_resp_0_bits_uop_pc_lob; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_taken = dcache_io_lsu_resp_0_bits_uop_taken; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_imm_packed = dcache_io_lsu_resp_0_bits_uop_imm_packed; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_csr_addr = dcache_io_lsu_resp_0_bits_uop_csr_addr; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_rob_idx = dcache_io_lsu_resp_0_bits_uop_rob_idx; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_ldq_idx = dcache_io_lsu_resp_0_bits_uop_ldq_idx; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_stq_idx = dcache_io_lsu_resp_0_bits_uop_stq_idx; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_rxq_idx = dcache_io_lsu_resp_0_bits_uop_rxq_idx; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_pdst = dcache_io_lsu_resp_0_bits_uop_pdst; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_prs1 = dcache_io_lsu_resp_0_bits_uop_prs1; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_prs2 = dcache_io_lsu_resp_0_bits_uop_prs2; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_prs3 = dcache_io_lsu_resp_0_bits_uop_prs3; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_ppred = dcache_io_lsu_resp_0_bits_uop_ppred; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_prs1_busy = dcache_io_lsu_resp_0_bits_uop_prs1_busy; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_prs2_busy = dcache_io_lsu_resp_0_bits_uop_prs2_busy; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_prs3_busy = dcache_io_lsu_resp_0_bits_uop_prs3_busy; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_ppred_busy = dcache_io_lsu_resp_0_bits_uop_ppred_busy; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_stale_pdst = dcache_io_lsu_resp_0_bits_uop_stale_pdst; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_exception = dcache_io_lsu_resp_0_bits_uop_exception; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_exc_cause = dcache_io_lsu_resp_0_bits_uop_exc_cause; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_bypassable = dcache_io_lsu_resp_0_bits_uop_bypassable; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_mem_cmd = dcache_io_lsu_resp_0_bits_uop_mem_cmd; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_mem_size = dcache_io_lsu_resp_0_bits_uop_mem_size; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_mem_signed = dcache_io_lsu_resp_0_bits_uop_mem_signed; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_is_fence = dcache_io_lsu_resp_0_bits_uop_is_fence; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_is_fencei = dcache_io_lsu_resp_0_bits_uop_is_fencei; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_is_amo = dcache_io_lsu_resp_0_bits_uop_is_amo; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_uses_ldq = dcache_io_lsu_resp_0_bits_uop_uses_ldq; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_uses_stq = dcache_io_lsu_resp_0_bits_uop_uses_stq; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_is_sys_pc2epc = dcache_io_lsu_resp_0_bits_uop_is_sys_pc2epc; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_is_unique = dcache_io_lsu_resp_0_bits_uop_is_unique; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_flush_on_commit = dcache_io_lsu_resp_0_bits_uop_flush_on_commit; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_ldst_is_rs1 = dcache_io_lsu_resp_0_bits_uop_ldst_is_rs1; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_ldst = dcache_io_lsu_resp_0_bits_uop_ldst; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_lrs1 = dcache_io_lsu_resp_0_bits_uop_lrs1; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_lrs2 = dcache_io_lsu_resp_0_bits_uop_lrs2; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_lrs3 = dcache_io_lsu_resp_0_bits_uop_lrs3; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_ldst_val = dcache_io_lsu_resp_0_bits_uop_ldst_val; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_dst_rtype = dcache_io_lsu_resp_0_bits_uop_dst_rtype; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_lrs1_rtype = dcache_io_lsu_resp_0_bits_uop_lrs1_rtype; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_lrs2_rtype = dcache_io_lsu_resp_0_bits_uop_lrs2_rtype; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_frs3_en = dcache_io_lsu_resp_0_bits_uop_frs3_en; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_fp_val = dcache_io_lsu_resp_0_bits_uop_fp_val; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_fp_single = dcache_io_lsu_resp_0_bits_uop_fp_single; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_xcpt_pf_if = dcache_io_lsu_resp_0_bits_uop_xcpt_pf_if; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_xcpt_ae_if = dcache_io_lsu_resp_0_bits_uop_xcpt_ae_if; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_xcpt_ma_if = dcache_io_lsu_resp_0_bits_uop_xcpt_ma_if; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_bp_debug_if = dcache_io_lsu_resp_0_bits_uop_bp_debug_if; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_bp_xcpt_if = dcache_io_lsu_resp_0_bits_uop_bp_xcpt_if; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_debug_fsrc = dcache_io_lsu_resp_0_bits_uop_debug_fsrc; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_uop_debug_tsrc = dcache_io_lsu_resp_0_bits_uop_debug_tsrc; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_data = dcache_io_lsu_resp_0_bits_data; // @[tile.scala 239:30]
  assign lsu_io_dmem_resp_0_bits_is_hella = dcache_io_lsu_resp_0_bits_is_hella; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_valid = dcache_io_lsu_nack_0_valid; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_switch = dcache_io_lsu_nack_0_bits_uop_switch; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_switch_off = dcache_io_lsu_nack_0_bits_uop_switch_off; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_is_unicore = dcache_io_lsu_nack_0_bits_uop_is_unicore; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_shift = dcache_io_lsu_nack_0_bits_uop_shift; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_lrs3_rtype = dcache_io_lsu_nack_0_bits_uop_lrs3_rtype; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_rflag = dcache_io_lsu_nack_0_bits_uop_rflag; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_wflag = dcache_io_lsu_nack_0_bits_uop_wflag; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_prflag = dcache_io_lsu_nack_0_bits_uop_prflag; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_pwflag = dcache_io_lsu_nack_0_bits_uop_pwflag; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_pflag_busy = dcache_io_lsu_nack_0_bits_uop_pflag_busy; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_stale_pflag = dcache_io_lsu_nack_0_bits_uop_stale_pflag; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_op1_sel = dcache_io_lsu_nack_0_bits_uop_op1_sel; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_op2_sel = dcache_io_lsu_nack_0_bits_uop_op2_sel; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_split_num = dcache_io_lsu_nack_0_bits_uop_split_num; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_self_index = dcache_io_lsu_nack_0_bits_uop_self_index; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_rob_inst_idx = dcache_io_lsu_nack_0_bits_uop_rob_inst_idx; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_address_num = dcache_io_lsu_nack_0_bits_uop_address_num; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_uopc = dcache_io_lsu_nack_0_bits_uop_uopc; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_inst = dcache_io_lsu_nack_0_bits_uop_inst; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_debug_inst = dcache_io_lsu_nack_0_bits_uop_debug_inst; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_is_rvc = dcache_io_lsu_nack_0_bits_uop_is_rvc; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_debug_pc = dcache_io_lsu_nack_0_bits_uop_debug_pc; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_iq_type = dcache_io_lsu_nack_0_bits_uop_iq_type; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_fu_code = dcache_io_lsu_nack_0_bits_uop_fu_code; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_ctrl_br_type = dcache_io_lsu_nack_0_bits_uop_ctrl_br_type; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_ctrl_op1_sel = dcache_io_lsu_nack_0_bits_uop_ctrl_op1_sel; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_ctrl_op2_sel = dcache_io_lsu_nack_0_bits_uop_ctrl_op2_sel; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_ctrl_imm_sel = dcache_io_lsu_nack_0_bits_uop_ctrl_imm_sel; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_ctrl_op_fcn = dcache_io_lsu_nack_0_bits_uop_ctrl_op_fcn; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_ctrl_fcn_dw = dcache_io_lsu_nack_0_bits_uop_ctrl_fcn_dw; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_ctrl_csr_cmd = dcache_io_lsu_nack_0_bits_uop_ctrl_csr_cmd; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_ctrl_is_load = dcache_io_lsu_nack_0_bits_uop_ctrl_is_load; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_ctrl_is_sta = dcache_io_lsu_nack_0_bits_uop_ctrl_is_sta; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_ctrl_is_std = dcache_io_lsu_nack_0_bits_uop_ctrl_is_std; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_ctrl_op3_sel = dcache_io_lsu_nack_0_bits_uop_ctrl_op3_sel; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_iw_state = dcache_io_lsu_nack_0_bits_uop_iw_state; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_iw_p1_poisoned = dcache_io_lsu_nack_0_bits_uop_iw_p1_poisoned; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_iw_p2_poisoned = dcache_io_lsu_nack_0_bits_uop_iw_p2_poisoned; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_is_br = dcache_io_lsu_nack_0_bits_uop_is_br; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_is_jalr = dcache_io_lsu_nack_0_bits_uop_is_jalr; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_is_jal = dcache_io_lsu_nack_0_bits_uop_is_jal; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_is_sfb = dcache_io_lsu_nack_0_bits_uop_is_sfb; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_br_mask = dcache_io_lsu_nack_0_bits_uop_br_mask; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_br_tag = dcache_io_lsu_nack_0_bits_uop_br_tag; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_ftq_idx = dcache_io_lsu_nack_0_bits_uop_ftq_idx; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_edge_inst = dcache_io_lsu_nack_0_bits_uop_edge_inst; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_pc_lob = dcache_io_lsu_nack_0_bits_uop_pc_lob; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_taken = dcache_io_lsu_nack_0_bits_uop_taken; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_imm_packed = dcache_io_lsu_nack_0_bits_uop_imm_packed; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_csr_addr = dcache_io_lsu_nack_0_bits_uop_csr_addr; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_rob_idx = dcache_io_lsu_nack_0_bits_uop_rob_idx; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_ldq_idx = dcache_io_lsu_nack_0_bits_uop_ldq_idx; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_stq_idx = dcache_io_lsu_nack_0_bits_uop_stq_idx; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_rxq_idx = dcache_io_lsu_nack_0_bits_uop_rxq_idx; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_pdst = dcache_io_lsu_nack_0_bits_uop_pdst; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_prs1 = dcache_io_lsu_nack_0_bits_uop_prs1; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_prs2 = dcache_io_lsu_nack_0_bits_uop_prs2; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_prs3 = dcache_io_lsu_nack_0_bits_uop_prs3; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_ppred = dcache_io_lsu_nack_0_bits_uop_ppred; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_prs1_busy = dcache_io_lsu_nack_0_bits_uop_prs1_busy; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_prs2_busy = dcache_io_lsu_nack_0_bits_uop_prs2_busy; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_prs3_busy = dcache_io_lsu_nack_0_bits_uop_prs3_busy; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_ppred_busy = dcache_io_lsu_nack_0_bits_uop_ppred_busy; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_stale_pdst = dcache_io_lsu_nack_0_bits_uop_stale_pdst; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_exception = dcache_io_lsu_nack_0_bits_uop_exception; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_exc_cause = dcache_io_lsu_nack_0_bits_uop_exc_cause; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_bypassable = dcache_io_lsu_nack_0_bits_uop_bypassable; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_mem_cmd = dcache_io_lsu_nack_0_bits_uop_mem_cmd; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_mem_size = dcache_io_lsu_nack_0_bits_uop_mem_size; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_mem_signed = dcache_io_lsu_nack_0_bits_uop_mem_signed; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_is_fence = dcache_io_lsu_nack_0_bits_uop_is_fence; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_is_fencei = dcache_io_lsu_nack_0_bits_uop_is_fencei; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_is_amo = dcache_io_lsu_nack_0_bits_uop_is_amo; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_uses_ldq = dcache_io_lsu_nack_0_bits_uop_uses_ldq; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_uses_stq = dcache_io_lsu_nack_0_bits_uop_uses_stq; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_is_sys_pc2epc = dcache_io_lsu_nack_0_bits_uop_is_sys_pc2epc; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_is_unique = dcache_io_lsu_nack_0_bits_uop_is_unique; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_flush_on_commit = dcache_io_lsu_nack_0_bits_uop_flush_on_commit; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_ldst_is_rs1 = dcache_io_lsu_nack_0_bits_uop_ldst_is_rs1; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_ldst = dcache_io_lsu_nack_0_bits_uop_ldst; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_lrs1 = dcache_io_lsu_nack_0_bits_uop_lrs1; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_lrs2 = dcache_io_lsu_nack_0_bits_uop_lrs2; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_lrs3 = dcache_io_lsu_nack_0_bits_uop_lrs3; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_ldst_val = dcache_io_lsu_nack_0_bits_uop_ldst_val; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_dst_rtype = dcache_io_lsu_nack_0_bits_uop_dst_rtype; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_lrs1_rtype = dcache_io_lsu_nack_0_bits_uop_lrs1_rtype; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_lrs2_rtype = dcache_io_lsu_nack_0_bits_uop_lrs2_rtype; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_frs3_en = dcache_io_lsu_nack_0_bits_uop_frs3_en; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_fp_val = dcache_io_lsu_nack_0_bits_uop_fp_val; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_fp_single = dcache_io_lsu_nack_0_bits_uop_fp_single; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_xcpt_pf_if = dcache_io_lsu_nack_0_bits_uop_xcpt_pf_if; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_xcpt_ae_if = dcache_io_lsu_nack_0_bits_uop_xcpt_ae_if; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_xcpt_ma_if = dcache_io_lsu_nack_0_bits_uop_xcpt_ma_if; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_bp_debug_if = dcache_io_lsu_nack_0_bits_uop_bp_debug_if; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_bp_xcpt_if = dcache_io_lsu_nack_0_bits_uop_bp_xcpt_if; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_debug_fsrc = dcache_io_lsu_nack_0_bits_uop_debug_fsrc; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_uop_debug_tsrc = dcache_io_lsu_nack_0_bits_uop_debug_tsrc; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_addr = dcache_io_lsu_nack_0_bits_addr; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_data = dcache_io_lsu_nack_0_bits_data; // @[tile.scala 239:30]
  assign lsu_io_dmem_nack_0_bits_is_hella = dcache_io_lsu_nack_0_bits_is_hella; // @[tile.scala 239:30]
  assign lsu_io_dmem_release_valid = dcache_io_lsu_release_valid; // @[tile.scala 239:30]
  assign lsu_io_dmem_release_bits_opcode = dcache_io_lsu_release_bits_opcode; // @[tile.scala 239:30]
  assign lsu_io_dmem_release_bits_param = dcache_io_lsu_release_bits_param; // @[tile.scala 239:30]
  assign lsu_io_dmem_release_bits_size = dcache_io_lsu_release_bits_size; // @[tile.scala 239:30]
  assign lsu_io_dmem_release_bits_source = dcache_io_lsu_release_bits_source; // @[tile.scala 239:30]
  assign lsu_io_dmem_release_bits_address = dcache_io_lsu_release_bits_address; // @[tile.scala 239:30]
  assign lsu_io_dmem_release_bits_data = dcache_io_lsu_release_bits_data; // @[tile.scala 239:30]
  assign lsu_io_dmem_release_bits_corrupt = dcache_io_lsu_release_bits_corrupt; // @[tile.scala 239:30]
  assign lsu_io_dmem_ordered = dcache_io_lsu_ordered; // @[tile.scala 239:30]
  assign lsu_io_dmem_perf_acquire = dcache_io_lsu_perf_acquire; // @[tile.scala 239:30]
  assign lsu_io_dmem_perf_release = dcache_io_lsu_perf_release; // @[tile.scala 239:30]
  assign lsu_io_hellacache_req_valid = hellaCacheArb_io_mem_req_valid; // @[tile.scala 238:21]
  assign lsu_io_hellacache_req_bits_addr = hellaCacheArb_io_mem_req_bits_addr; // @[tile.scala 238:21]
  assign lsu_io_hellacache_req_bits_tag = hellaCacheArb_io_mem_req_bits_tag; // @[tile.scala 238:21]
  assign lsu_io_hellacache_req_bits_cmd = hellaCacheArb_io_mem_req_bits_cmd; // @[tile.scala 238:21]
  assign lsu_io_hellacache_req_bits_size = hellaCacheArb_io_mem_req_bits_size; // @[tile.scala 238:21]
  assign lsu_io_hellacache_req_bits_signed = hellaCacheArb_io_mem_req_bits_signed; // @[tile.scala 238:21]
  assign lsu_io_hellacache_req_bits_dprv = hellaCacheArb_io_mem_req_bits_dprv; // @[tile.scala 238:21]
  assign lsu_io_hellacache_req_bits_phys = hellaCacheArb_io_mem_req_bits_phys; // @[tile.scala 238:21]
  assign lsu_io_hellacache_req_bits_no_alloc = hellaCacheArb_io_mem_req_bits_no_alloc; // @[tile.scala 238:21]
  assign lsu_io_hellacache_req_bits_no_xcpt = hellaCacheArb_io_mem_req_bits_no_xcpt; // @[tile.scala 238:21]
  assign lsu_io_hellacache_req_bits_data = hellaCacheArb_io_mem_req_bits_data; // @[tile.scala 238:21]
  assign lsu_io_hellacache_req_bits_mask = hellaCacheArb_io_mem_req_bits_mask; // @[tile.scala 238:21]
  assign lsu_io_hellacache_s1_kill = hellaCacheArb_io_mem_s1_kill; // @[tile.scala 238:21]
  assign lsu_io_hellacache_s1_data_data = hellaCacheArb_io_mem_s1_data_data; // @[tile.scala 238:21]
  assign lsu_io_hellacache_s1_data_mask = hellaCacheArb_io_mem_s1_data_mask; // @[tile.scala 238:21]
  assign lsu_io_hellacache_s2_kill = hellaCacheArb_io_mem_s2_kill; // @[tile.scala 238:21]
  assign lsu_io_hellacache_keep_clock_enabled = hellaCacheArb_io_mem_keep_clock_enabled; // @[tile.scala 238:21]
  assign ptw_clock = clock;
  assign ptw_reset = reset;
  assign ptw_io_requestor_0_req_valid = lsu_io_ptw_req_valid; // @[tile.scala 232:20]
  assign ptw_io_requestor_0_req_bits_valid = lsu_io_ptw_req_bits_valid; // @[tile.scala 232:20]
  assign ptw_io_requestor_0_req_bits_bits_addr = lsu_io_ptw_req_bits_bits_addr; // @[tile.scala 232:20]
  assign ptw_io_requestor_1_req_valid = frontend_io_ptw_req_valid; // @[tile.scala 232:20]
  assign ptw_io_requestor_1_req_bits_valid = frontend_io_ptw_req_bits_valid; // @[tile.scala 232:20]
  assign ptw_io_requestor_1_req_bits_bits_addr = frontend_io_ptw_req_bits_bits_addr; // @[tile.scala 232:20]
  assign ptw_io_requestor_2_req_valid = core_io_ptw_tlb_req_valid; // @[tile.scala 232:20]
  assign ptw_io_requestor_2_req_bits_valid = core_io_ptw_tlb_req_bits_valid; // @[tile.scala 232:20]
  assign ptw_io_requestor_2_req_bits_bits_addr = core_io_ptw_tlb_req_bits_bits_addr; // @[tile.scala 232:20]
  assign ptw_io_mem_req_ready = hellaCacheArb_io_requestor_0_req_ready; // @[tile.scala 237:30]
  assign ptw_io_mem_s2_nack = hellaCacheArb_io_requestor_0_s2_nack; // @[tile.scala 237:30]
  assign ptw_io_mem_s2_nack_cause_raw = hellaCacheArb_io_requestor_0_s2_nack_cause_raw; // @[tile.scala 237:30]
  assign ptw_io_mem_s2_uncached = hellaCacheArb_io_requestor_0_s2_uncached; // @[tile.scala 237:30]
  assign ptw_io_mem_s2_paddr = hellaCacheArb_io_requestor_0_s2_paddr; // @[tile.scala 237:30]
  assign ptw_io_mem_resp_valid = hellaCacheArb_io_requestor_0_resp_valid; // @[tile.scala 237:30]
  assign ptw_io_mem_resp_bits_addr = hellaCacheArb_io_requestor_0_resp_bits_addr; // @[tile.scala 237:30]
  assign ptw_io_mem_resp_bits_tag = hellaCacheArb_io_requestor_0_resp_bits_tag; // @[tile.scala 237:30]
  assign ptw_io_mem_resp_bits_cmd = hellaCacheArb_io_requestor_0_resp_bits_cmd; // @[tile.scala 237:30]
  assign ptw_io_mem_resp_bits_size = hellaCacheArb_io_requestor_0_resp_bits_size; // @[tile.scala 237:30]
  assign ptw_io_mem_resp_bits_signed = hellaCacheArb_io_requestor_0_resp_bits_signed; // @[tile.scala 237:30]
  assign ptw_io_mem_resp_bits_dprv = hellaCacheArb_io_requestor_0_resp_bits_dprv; // @[tile.scala 237:30]
  assign ptw_io_mem_resp_bits_data = hellaCacheArb_io_requestor_0_resp_bits_data; // @[tile.scala 237:30]
  assign ptw_io_mem_resp_bits_mask = hellaCacheArb_io_requestor_0_resp_bits_mask; // @[tile.scala 237:30]
  assign ptw_io_mem_resp_bits_replay = hellaCacheArb_io_requestor_0_resp_bits_replay; // @[tile.scala 237:30]
  assign ptw_io_mem_resp_bits_has_data = hellaCacheArb_io_requestor_0_resp_bits_has_data; // @[tile.scala 237:30]
  assign ptw_io_mem_resp_bits_data_word_bypass = hellaCacheArb_io_requestor_0_resp_bits_data_word_bypass; // @[tile.scala 237:30]
  assign ptw_io_mem_resp_bits_data_raw = hellaCacheArb_io_requestor_0_resp_bits_data_raw; // @[tile.scala 237:30]
  assign ptw_io_mem_resp_bits_store_data = hellaCacheArb_io_requestor_0_resp_bits_store_data; // @[tile.scala 237:30]
  assign ptw_io_mem_replay_next = hellaCacheArb_io_requestor_0_replay_next; // @[tile.scala 237:30]
  assign ptw_io_mem_s2_xcpt_ma_ld = hellaCacheArb_io_requestor_0_s2_xcpt_ma_ld; // @[tile.scala 237:30]
  assign ptw_io_mem_s2_xcpt_ma_st = hellaCacheArb_io_requestor_0_s2_xcpt_ma_st; // @[tile.scala 237:30]
  assign ptw_io_mem_s2_xcpt_pf_ld = hellaCacheArb_io_requestor_0_s2_xcpt_pf_ld; // @[tile.scala 237:30]
  assign ptw_io_mem_s2_xcpt_pf_st = hellaCacheArb_io_requestor_0_s2_xcpt_pf_st; // @[tile.scala 237:30]
  assign ptw_io_mem_s2_xcpt_ae_ld = hellaCacheArb_io_requestor_0_s2_xcpt_ae_ld; // @[tile.scala 237:30]
  assign ptw_io_mem_s2_xcpt_ae_st = hellaCacheArb_io_requestor_0_s2_xcpt_ae_st; // @[tile.scala 237:30]
  assign ptw_io_mem_ordered = hellaCacheArb_io_requestor_0_ordered; // @[tile.scala 237:30]
  assign ptw_io_mem_perf_acquire = hellaCacheArb_io_requestor_0_perf_acquire; // @[tile.scala 237:30]
  assign ptw_io_mem_perf_release = hellaCacheArb_io_requestor_0_perf_release; // @[tile.scala 237:30]
  assign ptw_io_mem_perf_grant = hellaCacheArb_io_requestor_0_perf_grant; // @[tile.scala 237:30]
  assign ptw_io_mem_perf_tlbMiss = hellaCacheArb_io_requestor_0_perf_tlbMiss; // @[tile.scala 237:30]
  assign ptw_io_mem_perf_blocked = hellaCacheArb_io_requestor_0_perf_blocked; // @[tile.scala 237:30]
  assign ptw_io_mem_perf_canAcceptStoreThenLoad = hellaCacheArb_io_requestor_0_perf_canAcceptStoreThenLoad; // @[tile.scala 237:30]
  assign ptw_io_mem_perf_canAcceptStoreThenRMW = hellaCacheArb_io_requestor_0_perf_canAcceptStoreThenRMW; // @[tile.scala 237:30]
  assign ptw_io_mem_perf_canAcceptLoadThenLoad = hellaCacheArb_io_requestor_0_perf_canAcceptLoadThenLoad; // @[tile.scala 237:30]
  assign ptw_io_mem_perf_storeBufferEmptyAfterLoad = hellaCacheArb_io_requestor_0_perf_storeBufferEmptyAfterLoad; // @[tile.scala 237:30]
  assign ptw_io_mem_perf_storeBufferEmptyAfterStore = hellaCacheArb_io_requestor_0_perf_storeBufferEmptyAfterStore; // @[tile.scala 237:30]
  assign ptw_io_mem_clock_enabled = hellaCacheArb_io_requestor_0_clock_enabled; // @[tile.scala 237:30]
  assign ptw_io_dpath_ptbr_mode = core_io_ptw_ptbr_mode; // @[tile.scala 231:15]
  assign ptw_io_dpath_ptbr_asid = core_io_ptw_ptbr_asid; // @[tile.scala 231:15]
  assign ptw_io_dpath_ptbr_ppn = core_io_ptw_ptbr_ppn; // @[tile.scala 231:15]
  assign ptw_io_dpath_sfence_valid = core_io_ptw_sfence_valid; // @[tile.scala 231:15]
  assign ptw_io_dpath_sfence_bits_rs1 = core_io_ptw_sfence_bits_rs1; // @[tile.scala 231:15]
  assign ptw_io_dpath_sfence_bits_rs2 = core_io_ptw_sfence_bits_rs2; // @[tile.scala 231:15]
  assign ptw_io_dpath_sfence_bits_addr = core_io_ptw_sfence_bits_addr; // @[tile.scala 231:15]
  assign ptw_io_dpath_sfence_bits_asid = core_io_ptw_sfence_bits_asid; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_debug = core_io_ptw_status_debug; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_cease = core_io_ptw_status_cease; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_wfi = core_io_ptw_status_wfi; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_isa = core_io_ptw_status_isa; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_dprv = core_io_ptw_status_dprv; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_prv = core_io_ptw_status_prv; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_sd = core_io_ptw_status_sd; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_zero2 = core_io_ptw_status_zero2; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_sxl = core_io_ptw_status_sxl; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_uxl = core_io_ptw_status_uxl; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_sd_rv32 = core_io_ptw_status_sd_rv32; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_zero1 = core_io_ptw_status_zero1; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_tsr = core_io_ptw_status_tsr; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_tw = core_io_ptw_status_tw; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_tvm = core_io_ptw_status_tvm; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_mxr = core_io_ptw_status_mxr; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_sum = core_io_ptw_status_sum; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_mprv = core_io_ptw_status_mprv; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_xs = core_io_ptw_status_xs; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_fs = core_io_ptw_status_fs; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_mpp = core_io_ptw_status_mpp; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_vs = core_io_ptw_status_vs; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_spp = core_io_ptw_status_spp; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_mpie = core_io_ptw_status_mpie; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_hpie = core_io_ptw_status_hpie; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_spie = core_io_ptw_status_spie; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_upie = core_io_ptw_status_upie; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_mie = core_io_ptw_status_mie; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_hie = core_io_ptw_status_hie; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_sie = core_io_ptw_status_sie; // @[tile.scala 231:15]
  assign ptw_io_dpath_status_uie = core_io_ptw_status_uie; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_0_cfg_l = core_io_ptw_pmp_0_cfg_l; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_0_cfg_res = core_io_ptw_pmp_0_cfg_res; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_0_cfg_a = core_io_ptw_pmp_0_cfg_a; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_0_cfg_x = core_io_ptw_pmp_0_cfg_x; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_0_cfg_w = core_io_ptw_pmp_0_cfg_w; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_0_cfg_r = core_io_ptw_pmp_0_cfg_r; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_0_addr = core_io_ptw_pmp_0_addr; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_0_mask = core_io_ptw_pmp_0_mask; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_1_cfg_l = core_io_ptw_pmp_1_cfg_l; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_1_cfg_res = core_io_ptw_pmp_1_cfg_res; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_1_cfg_a = core_io_ptw_pmp_1_cfg_a; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_1_cfg_x = core_io_ptw_pmp_1_cfg_x; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_1_cfg_w = core_io_ptw_pmp_1_cfg_w; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_1_cfg_r = core_io_ptw_pmp_1_cfg_r; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_1_addr = core_io_ptw_pmp_1_addr; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_1_mask = core_io_ptw_pmp_1_mask; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_2_cfg_l = core_io_ptw_pmp_2_cfg_l; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_2_cfg_res = core_io_ptw_pmp_2_cfg_res; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_2_cfg_a = core_io_ptw_pmp_2_cfg_a; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_2_cfg_x = core_io_ptw_pmp_2_cfg_x; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_2_cfg_w = core_io_ptw_pmp_2_cfg_w; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_2_cfg_r = core_io_ptw_pmp_2_cfg_r; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_2_addr = core_io_ptw_pmp_2_addr; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_2_mask = core_io_ptw_pmp_2_mask; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_3_cfg_l = core_io_ptw_pmp_3_cfg_l; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_3_cfg_res = core_io_ptw_pmp_3_cfg_res; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_3_cfg_a = core_io_ptw_pmp_3_cfg_a; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_3_cfg_x = core_io_ptw_pmp_3_cfg_x; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_3_cfg_w = core_io_ptw_pmp_3_cfg_w; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_3_cfg_r = core_io_ptw_pmp_3_cfg_r; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_3_addr = core_io_ptw_pmp_3_addr; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_3_mask = core_io_ptw_pmp_3_mask; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_4_cfg_l = core_io_ptw_pmp_4_cfg_l; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_4_cfg_res = core_io_ptw_pmp_4_cfg_res; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_4_cfg_a = core_io_ptw_pmp_4_cfg_a; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_4_cfg_x = core_io_ptw_pmp_4_cfg_x; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_4_cfg_w = core_io_ptw_pmp_4_cfg_w; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_4_cfg_r = core_io_ptw_pmp_4_cfg_r; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_4_addr = core_io_ptw_pmp_4_addr; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_4_mask = core_io_ptw_pmp_4_mask; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_5_cfg_l = core_io_ptw_pmp_5_cfg_l; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_5_cfg_res = core_io_ptw_pmp_5_cfg_res; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_5_cfg_a = core_io_ptw_pmp_5_cfg_a; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_5_cfg_x = core_io_ptw_pmp_5_cfg_x; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_5_cfg_w = core_io_ptw_pmp_5_cfg_w; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_5_cfg_r = core_io_ptw_pmp_5_cfg_r; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_5_addr = core_io_ptw_pmp_5_addr; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_5_mask = core_io_ptw_pmp_5_mask; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_6_cfg_l = core_io_ptw_pmp_6_cfg_l; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_6_cfg_res = core_io_ptw_pmp_6_cfg_res; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_6_cfg_a = core_io_ptw_pmp_6_cfg_a; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_6_cfg_x = core_io_ptw_pmp_6_cfg_x; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_6_cfg_w = core_io_ptw_pmp_6_cfg_w; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_6_cfg_r = core_io_ptw_pmp_6_cfg_r; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_6_addr = core_io_ptw_pmp_6_addr; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_6_mask = core_io_ptw_pmp_6_mask; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_7_cfg_l = core_io_ptw_pmp_7_cfg_l; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_7_cfg_res = core_io_ptw_pmp_7_cfg_res; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_7_cfg_a = core_io_ptw_pmp_7_cfg_a; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_7_cfg_x = core_io_ptw_pmp_7_cfg_x; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_7_cfg_w = core_io_ptw_pmp_7_cfg_w; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_7_cfg_r = core_io_ptw_pmp_7_cfg_r; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_7_addr = core_io_ptw_pmp_7_addr; // @[tile.scala 231:15]
  assign ptw_io_dpath_pmp_7_mask = core_io_ptw_pmp_7_mask; // @[tile.scala 231:15]
  assign ptw_io_dpath_customCSRs_csrs_0_wen = core_io_ptw_customCSRs_csrs_0_wen; // @[tile.scala 231:15]
  assign ptw_io_dpath_customCSRs_csrs_0_wdata = core_io_ptw_customCSRs_csrs_0_wdata; // @[tile.scala 231:15]
  assign ptw_io_dpath_customCSRs_csrs_0_value = core_io_ptw_customCSRs_csrs_0_value; // @[tile.scala 231:15]
  assign hellaCacheArb_clock = clock;
  assign hellaCacheArb_reset = reset;
  assign hellaCacheArb_io_requestor_0_req_valid = ptw_io_mem_req_valid; // @[tile.scala 237:30]
  assign hellaCacheArb_io_requestor_0_req_bits_addr = ptw_io_mem_req_bits_addr; // @[tile.scala 237:30]
  assign hellaCacheArb_io_requestor_0_req_bits_tag = ptw_io_mem_req_bits_tag; // @[tile.scala 237:30]
  assign hellaCacheArb_io_requestor_0_req_bits_cmd = ptw_io_mem_req_bits_cmd; // @[tile.scala 237:30]
  assign hellaCacheArb_io_requestor_0_req_bits_size = ptw_io_mem_req_bits_size; // @[tile.scala 237:30]
  assign hellaCacheArb_io_requestor_0_req_bits_signed = ptw_io_mem_req_bits_signed; // @[tile.scala 237:30]
  assign hellaCacheArb_io_requestor_0_req_bits_dprv = ptw_io_mem_req_bits_dprv; // @[tile.scala 237:30]
  assign hellaCacheArb_io_requestor_0_req_bits_phys = ptw_io_mem_req_bits_phys; // @[tile.scala 237:30]
  assign hellaCacheArb_io_requestor_0_req_bits_no_alloc = ptw_io_mem_req_bits_no_alloc; // @[tile.scala 237:30]
  assign hellaCacheArb_io_requestor_0_req_bits_no_xcpt = ptw_io_mem_req_bits_no_xcpt; // @[tile.scala 237:30]
  assign hellaCacheArb_io_requestor_0_req_bits_data = ptw_io_mem_req_bits_data; // @[tile.scala 237:30]
  assign hellaCacheArb_io_requestor_0_req_bits_mask = ptw_io_mem_req_bits_mask; // @[tile.scala 237:30]
  assign hellaCacheArb_io_requestor_0_s1_kill = ptw_io_mem_s1_kill; // @[tile.scala 237:30]
  assign hellaCacheArb_io_requestor_0_s1_data_data = ptw_io_mem_s1_data_data; // @[tile.scala 237:30]
  assign hellaCacheArb_io_requestor_0_s1_data_mask = ptw_io_mem_s1_data_mask; // @[tile.scala 237:30]
  assign hellaCacheArb_io_requestor_0_s2_kill = ptw_io_mem_s2_kill; // @[tile.scala 237:30]
  assign hellaCacheArb_io_requestor_0_keep_clock_enabled = ptw_io_mem_keep_clock_enabled; // @[tile.scala 237:30]
  assign hellaCacheArb_io_mem_req_ready = lsu_io_hellacache_req_ready; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_s2_nack = lsu_io_hellacache_s2_nack; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_s2_nack_cause_raw = lsu_io_hellacache_s2_nack_cause_raw; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_s2_uncached = lsu_io_hellacache_s2_uncached; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_s2_paddr = lsu_io_hellacache_s2_paddr; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_resp_valid = lsu_io_hellacache_resp_valid; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_resp_bits_addr = lsu_io_hellacache_resp_bits_addr; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_resp_bits_tag = lsu_io_hellacache_resp_bits_tag; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_resp_bits_cmd = lsu_io_hellacache_resp_bits_cmd; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_resp_bits_size = lsu_io_hellacache_resp_bits_size; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_resp_bits_signed = lsu_io_hellacache_resp_bits_signed; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_resp_bits_dprv = lsu_io_hellacache_resp_bits_dprv; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_resp_bits_data = lsu_io_hellacache_resp_bits_data; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_resp_bits_mask = lsu_io_hellacache_resp_bits_mask; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_resp_bits_replay = lsu_io_hellacache_resp_bits_replay; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_resp_bits_has_data = lsu_io_hellacache_resp_bits_has_data; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_resp_bits_data_word_bypass = lsu_io_hellacache_resp_bits_data_word_bypass; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_resp_bits_data_raw = lsu_io_hellacache_resp_bits_data_raw; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_resp_bits_store_data = lsu_io_hellacache_resp_bits_store_data; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_replay_next = lsu_io_hellacache_replay_next; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_s2_xcpt_ma_ld = lsu_io_hellacache_s2_xcpt_ma_ld; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_s2_xcpt_ma_st = lsu_io_hellacache_s2_xcpt_ma_st; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_s2_xcpt_pf_ld = lsu_io_hellacache_s2_xcpt_pf_ld; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_s2_xcpt_pf_st = lsu_io_hellacache_s2_xcpt_pf_st; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_s2_xcpt_ae_ld = lsu_io_hellacache_s2_xcpt_ae_ld; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_s2_xcpt_ae_st = lsu_io_hellacache_s2_xcpt_ae_st; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_ordered = lsu_io_hellacache_ordered; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_perf_acquire = lsu_io_hellacache_perf_acquire; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_perf_release = lsu_io_hellacache_perf_release; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_perf_grant = lsu_io_hellacache_perf_grant; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_perf_tlbMiss = lsu_io_hellacache_perf_tlbMiss; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_perf_blocked = lsu_io_hellacache_perf_blocked; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_perf_canAcceptStoreThenLoad = lsu_io_hellacache_perf_canAcceptStoreThenLoad; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_perf_canAcceptStoreThenRMW = lsu_io_hellacache_perf_canAcceptStoreThenRMW; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_perf_canAcceptLoadThenLoad = lsu_io_hellacache_perf_canAcceptLoadThenLoad; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_perf_storeBufferEmptyAfterLoad = lsu_io_hellacache_perf_storeBufferEmptyAfterLoad; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_perf_storeBufferEmptyAfterStore = lsu_io_hellacache_perf_storeBufferEmptyAfterStore; // @[tile.scala 238:21]
  assign hellaCacheArb_io_mem_clock_enabled = lsu_io_hellacache_clock_enabled; // @[tile.scala 238:21]
endmodule
