module RegisterRead(
  input         clock,
  input         reset,
  input         io_iss_valids_0,
  input         io_iss_valids_1,
  input         io_iss_valids_2,
  input         io_iss_uops_0_switch,
  input         io_iss_uops_0_switch_off,
  input         io_iss_uops_0_is_unicore,
  input  [2:0]  io_iss_uops_0_shift,
  input  [1:0]  io_iss_uops_0_lrs3_rtype,
  input         io_iss_uops_0_rflag,
  input         io_iss_uops_0_wflag,
  input  [3:0]  io_iss_uops_0_prflag,
  input  [3:0]  io_iss_uops_0_pwflag,
  input         io_iss_uops_0_pflag_busy,
  input  [3:0]  io_iss_uops_0_stale_pflag,
  input  [3:0]  io_iss_uops_0_op1_sel,
  input  [3:0]  io_iss_uops_0_op2_sel,
  input  [5:0]  io_iss_uops_0_split_num,
  input  [5:0]  io_iss_uops_0_self_index,
  input  [5:0]  io_iss_uops_0_rob_inst_idx,
  input  [5:0]  io_iss_uops_0_address_num,
  input  [6:0]  io_iss_uops_0_uopc,
  input  [31:0] io_iss_uops_0_inst,
  input  [31:0] io_iss_uops_0_debug_inst,
  input         io_iss_uops_0_is_rvc,
  input  [39:0] io_iss_uops_0_debug_pc,
  input  [2:0]  io_iss_uops_0_iq_type,
  input  [9:0]  io_iss_uops_0_fu_code,
  input  [3:0]  io_iss_uops_0_ctrl_br_type,
  input  [1:0]  io_iss_uops_0_ctrl_op1_sel,
  input  [2:0]  io_iss_uops_0_ctrl_op2_sel,
  input  [2:0]  io_iss_uops_0_ctrl_imm_sel,
  input  [3:0]  io_iss_uops_0_ctrl_op_fcn,
  input         io_iss_uops_0_ctrl_fcn_dw,
  input  [2:0]  io_iss_uops_0_ctrl_csr_cmd,
  input         io_iss_uops_0_ctrl_is_load,
  input         io_iss_uops_0_ctrl_is_sta,
  input         io_iss_uops_0_ctrl_is_std,
  input  [1:0]  io_iss_uops_0_ctrl_op3_sel,
  input  [1:0]  io_iss_uops_0_iw_state,
  input         io_iss_uops_0_iw_p1_poisoned,
  input         io_iss_uops_0_iw_p2_poisoned,
  input         io_iss_uops_0_is_br,
  input         io_iss_uops_0_is_jalr,
  input         io_iss_uops_0_is_jal,
  input         io_iss_uops_0_is_sfb,
  input  [11:0] io_iss_uops_0_br_mask,
  input  [3:0]  io_iss_uops_0_br_tag,
  input  [4:0]  io_iss_uops_0_ftq_idx,
  input         io_iss_uops_0_edge_inst,
  input  [5:0]  io_iss_uops_0_pc_lob,
  input         io_iss_uops_0_taken,
  input  [19:0] io_iss_uops_0_imm_packed,
  input  [11:0] io_iss_uops_0_csr_addr,
  input  [5:0]  io_iss_uops_0_rob_idx,
  input  [4:0]  io_iss_uops_0_ldq_idx,
  input  [4:0]  io_iss_uops_0_stq_idx,
  input  [1:0]  io_iss_uops_0_rxq_idx,
  input  [6:0]  io_iss_uops_0_pdst,
  input  [6:0]  io_iss_uops_0_prs1,
  input  [6:0]  io_iss_uops_0_prs2,
  input  [6:0]  io_iss_uops_0_prs3,
  input  [4:0]  io_iss_uops_0_ppred,
  input         io_iss_uops_0_prs1_busy,
  input         io_iss_uops_0_prs2_busy,
  input         io_iss_uops_0_prs3_busy,
  input         io_iss_uops_0_ppred_busy,
  input  [6:0]  io_iss_uops_0_stale_pdst,
  input         io_iss_uops_0_exception,
  input  [63:0] io_iss_uops_0_exc_cause,
  input         io_iss_uops_0_bypassable,
  input  [4:0]  io_iss_uops_0_mem_cmd,
  input  [1:0]  io_iss_uops_0_mem_size,
  input         io_iss_uops_0_mem_signed,
  input         io_iss_uops_0_is_fence,
  input         io_iss_uops_0_is_fencei,
  input         io_iss_uops_0_is_amo,
  input         io_iss_uops_0_uses_ldq,
  input         io_iss_uops_0_uses_stq,
  input         io_iss_uops_0_is_sys_pc2epc,
  input         io_iss_uops_0_is_unique,
  input         io_iss_uops_0_flush_on_commit,
  input         io_iss_uops_0_ldst_is_rs1,
  input  [5:0]  io_iss_uops_0_ldst,
  input  [5:0]  io_iss_uops_0_lrs1,
  input  [5:0]  io_iss_uops_0_lrs2,
  input  [5:0]  io_iss_uops_0_lrs3,
  input         io_iss_uops_0_ldst_val,
  input  [1:0]  io_iss_uops_0_dst_rtype,
  input  [1:0]  io_iss_uops_0_lrs1_rtype,
  input  [1:0]  io_iss_uops_0_lrs2_rtype,
  input         io_iss_uops_0_frs3_en,
  input         io_iss_uops_0_fp_val,
  input         io_iss_uops_0_fp_single,
  input         io_iss_uops_0_xcpt_pf_if,
  input         io_iss_uops_0_xcpt_ae_if,
  input         io_iss_uops_0_xcpt_ma_if,
  input         io_iss_uops_0_bp_debug_if,
  input         io_iss_uops_0_bp_xcpt_if,
  input  [1:0]  io_iss_uops_0_debug_fsrc,
  input  [1:0]  io_iss_uops_0_debug_tsrc,
  input         io_iss_uops_1_switch,
  input         io_iss_uops_1_switch_off,
  input         io_iss_uops_1_is_unicore,
  input  [2:0]  io_iss_uops_1_shift,
  input  [1:0]  io_iss_uops_1_lrs3_rtype,
  input         io_iss_uops_1_rflag,
  input         io_iss_uops_1_wflag,
  input  [3:0]  io_iss_uops_1_prflag,
  input  [3:0]  io_iss_uops_1_pwflag,
  input         io_iss_uops_1_pflag_busy,
  input  [3:0]  io_iss_uops_1_stale_pflag,
  input  [3:0]  io_iss_uops_1_op1_sel,
  input  [3:0]  io_iss_uops_1_op2_sel,
  input  [5:0]  io_iss_uops_1_split_num,
  input  [5:0]  io_iss_uops_1_self_index,
  input  [5:0]  io_iss_uops_1_rob_inst_idx,
  input  [5:0]  io_iss_uops_1_address_num,
  input  [6:0]  io_iss_uops_1_uopc,
  input  [31:0] io_iss_uops_1_inst,
  input  [31:0] io_iss_uops_1_debug_inst,
  input         io_iss_uops_1_is_rvc,
  input  [39:0] io_iss_uops_1_debug_pc,
  input  [2:0]  io_iss_uops_1_iq_type,
  input  [9:0]  io_iss_uops_1_fu_code,
  input  [3:0]  io_iss_uops_1_ctrl_br_type,
  input  [1:0]  io_iss_uops_1_ctrl_op1_sel,
  input  [2:0]  io_iss_uops_1_ctrl_op2_sel,
  input  [2:0]  io_iss_uops_1_ctrl_imm_sel,
  input  [3:0]  io_iss_uops_1_ctrl_op_fcn,
  input         io_iss_uops_1_ctrl_fcn_dw,
  input  [2:0]  io_iss_uops_1_ctrl_csr_cmd,
  input         io_iss_uops_1_ctrl_is_load,
  input         io_iss_uops_1_ctrl_is_sta,
  input         io_iss_uops_1_ctrl_is_std,
  input  [1:0]  io_iss_uops_1_ctrl_op3_sel,
  input  [1:0]  io_iss_uops_1_iw_state,
  input         io_iss_uops_1_iw_p1_poisoned,
  input         io_iss_uops_1_iw_p2_poisoned,
  input         io_iss_uops_1_is_br,
  input         io_iss_uops_1_is_jalr,
  input         io_iss_uops_1_is_jal,
  input         io_iss_uops_1_is_sfb,
  input  [11:0] io_iss_uops_1_br_mask,
  input  [3:0]  io_iss_uops_1_br_tag,
  input  [4:0]  io_iss_uops_1_ftq_idx,
  input         io_iss_uops_1_edge_inst,
  input  [5:0]  io_iss_uops_1_pc_lob,
  input         io_iss_uops_1_taken,
  input  [19:0] io_iss_uops_1_imm_packed,
  input  [11:0] io_iss_uops_1_csr_addr,
  input  [5:0]  io_iss_uops_1_rob_idx,
  input  [4:0]  io_iss_uops_1_ldq_idx,
  input  [4:0]  io_iss_uops_1_stq_idx,
  input  [1:0]  io_iss_uops_1_rxq_idx,
  input  [6:0]  io_iss_uops_1_pdst,
  input  [6:0]  io_iss_uops_1_prs1,
  input  [6:0]  io_iss_uops_1_prs2,
  input  [6:0]  io_iss_uops_1_prs3,
  input  [4:0]  io_iss_uops_1_ppred,
  input         io_iss_uops_1_prs1_busy,
  input         io_iss_uops_1_prs2_busy,
  input         io_iss_uops_1_prs3_busy,
  input         io_iss_uops_1_ppred_busy,
  input  [6:0]  io_iss_uops_1_stale_pdst,
  input         io_iss_uops_1_exception,
  input  [63:0] io_iss_uops_1_exc_cause,
  input         io_iss_uops_1_bypassable,
  input  [4:0]  io_iss_uops_1_mem_cmd,
  input  [1:0]  io_iss_uops_1_mem_size,
  input         io_iss_uops_1_mem_signed,
  input         io_iss_uops_1_is_fence,
  input         io_iss_uops_1_is_fencei,
  input         io_iss_uops_1_is_amo,
  input         io_iss_uops_1_uses_ldq,
  input         io_iss_uops_1_uses_stq,
  input         io_iss_uops_1_is_sys_pc2epc,
  input         io_iss_uops_1_is_unique,
  input         io_iss_uops_1_flush_on_commit,
  input         io_iss_uops_1_ldst_is_rs1,
  input  [5:0]  io_iss_uops_1_ldst,
  input  [5:0]  io_iss_uops_1_lrs1,
  input  [5:0]  io_iss_uops_1_lrs2,
  input  [5:0]  io_iss_uops_1_lrs3,
  input         io_iss_uops_1_ldst_val,
  input  [1:0]  io_iss_uops_1_dst_rtype,
  input  [1:0]  io_iss_uops_1_lrs1_rtype,
  input  [1:0]  io_iss_uops_1_lrs2_rtype,
  input         io_iss_uops_1_frs3_en,
  input         io_iss_uops_1_fp_val,
  input         io_iss_uops_1_fp_single,
  input         io_iss_uops_1_xcpt_pf_if,
  input         io_iss_uops_1_xcpt_ae_if,
  input         io_iss_uops_1_xcpt_ma_if,
  input         io_iss_uops_1_bp_debug_if,
  input         io_iss_uops_1_bp_xcpt_if,
  input  [1:0]  io_iss_uops_1_debug_fsrc,
  input  [1:0]  io_iss_uops_1_debug_tsrc,
  input         io_iss_uops_2_switch,
  input         io_iss_uops_2_switch_off,
  input         io_iss_uops_2_is_unicore,
  input  [2:0]  io_iss_uops_2_shift,
  input  [1:0]  io_iss_uops_2_lrs3_rtype,
  input         io_iss_uops_2_rflag,
  input         io_iss_uops_2_wflag,
  input  [3:0]  io_iss_uops_2_prflag,
  input  [3:0]  io_iss_uops_2_pwflag,
  input         io_iss_uops_2_pflag_busy,
  input  [3:0]  io_iss_uops_2_stale_pflag,
  input  [3:0]  io_iss_uops_2_op1_sel,
  input  [3:0]  io_iss_uops_2_op2_sel,
  input  [5:0]  io_iss_uops_2_split_num,
  input  [5:0]  io_iss_uops_2_self_index,
  input  [5:0]  io_iss_uops_2_rob_inst_idx,
  input  [5:0]  io_iss_uops_2_address_num,
  input  [6:0]  io_iss_uops_2_uopc,
  input  [31:0] io_iss_uops_2_inst,
  input  [31:0] io_iss_uops_2_debug_inst,
  input         io_iss_uops_2_is_rvc,
  input  [39:0] io_iss_uops_2_debug_pc,
  input  [2:0]  io_iss_uops_2_iq_type,
  input  [9:0]  io_iss_uops_2_fu_code,
  input  [3:0]  io_iss_uops_2_ctrl_br_type,
  input  [1:0]  io_iss_uops_2_ctrl_op1_sel,
  input  [2:0]  io_iss_uops_2_ctrl_op2_sel,
  input  [2:0]  io_iss_uops_2_ctrl_imm_sel,
  input  [3:0]  io_iss_uops_2_ctrl_op_fcn,
  input         io_iss_uops_2_ctrl_fcn_dw,
  input  [2:0]  io_iss_uops_2_ctrl_csr_cmd,
  input         io_iss_uops_2_ctrl_is_load,
  input         io_iss_uops_2_ctrl_is_sta,
  input         io_iss_uops_2_ctrl_is_std,
  input  [1:0]  io_iss_uops_2_ctrl_op3_sel,
  input  [1:0]  io_iss_uops_2_iw_state,
  input         io_iss_uops_2_iw_p1_poisoned,
  input         io_iss_uops_2_iw_p2_poisoned,
  input         io_iss_uops_2_is_br,
  input         io_iss_uops_2_is_jalr,
  input         io_iss_uops_2_is_jal,
  input         io_iss_uops_2_is_sfb,
  input  [11:0] io_iss_uops_2_br_mask,
  input  [3:0]  io_iss_uops_2_br_tag,
  input  [4:0]  io_iss_uops_2_ftq_idx,
  input         io_iss_uops_2_edge_inst,
  input  [5:0]  io_iss_uops_2_pc_lob,
  input         io_iss_uops_2_taken,
  input  [19:0] io_iss_uops_2_imm_packed,
  input  [11:0] io_iss_uops_2_csr_addr,
  input  [5:0]  io_iss_uops_2_rob_idx,
  input  [4:0]  io_iss_uops_2_ldq_idx,
  input  [4:0]  io_iss_uops_2_stq_idx,
  input  [1:0]  io_iss_uops_2_rxq_idx,
  input  [6:0]  io_iss_uops_2_pdst,
  input  [6:0]  io_iss_uops_2_prs1,
  input  [6:0]  io_iss_uops_2_prs2,
  input  [6:0]  io_iss_uops_2_prs3,
  input  [4:0]  io_iss_uops_2_ppred,
  input         io_iss_uops_2_prs1_busy,
  input         io_iss_uops_2_prs2_busy,
  input         io_iss_uops_2_prs3_busy,
  input         io_iss_uops_2_ppred_busy,
  input  [6:0]  io_iss_uops_2_stale_pdst,
  input         io_iss_uops_2_exception,
  input  [63:0] io_iss_uops_2_exc_cause,
  input         io_iss_uops_2_bypassable,
  input  [4:0]  io_iss_uops_2_mem_cmd,
  input  [1:0]  io_iss_uops_2_mem_size,
  input         io_iss_uops_2_mem_signed,
  input         io_iss_uops_2_is_fence,
  input         io_iss_uops_2_is_fencei,
  input         io_iss_uops_2_is_amo,
  input         io_iss_uops_2_uses_ldq,
  input         io_iss_uops_2_uses_stq,
  input         io_iss_uops_2_is_sys_pc2epc,
  input         io_iss_uops_2_is_unique,
  input         io_iss_uops_2_flush_on_commit,
  input         io_iss_uops_2_ldst_is_rs1,
  input  [5:0]  io_iss_uops_2_ldst,
  input  [5:0]  io_iss_uops_2_lrs1,
  input  [5:0]  io_iss_uops_2_lrs2,
  input  [5:0]  io_iss_uops_2_lrs3,
  input         io_iss_uops_2_ldst_val,
  input  [1:0]  io_iss_uops_2_dst_rtype,
  input  [1:0]  io_iss_uops_2_lrs1_rtype,
  input  [1:0]  io_iss_uops_2_lrs2_rtype,
  input         io_iss_uops_2_frs3_en,
  input         io_iss_uops_2_fp_val,
  input         io_iss_uops_2_fp_single,
  input         io_iss_uops_2_xcpt_pf_if,
  input         io_iss_uops_2_xcpt_ae_if,
  input         io_iss_uops_2_xcpt_ma_if,
  input         io_iss_uops_2_bp_debug_if,
  input         io_iss_uops_2_bp_xcpt_if,
  input  [1:0]  io_iss_uops_2_debug_fsrc,
  input  [1:0]  io_iss_uops_2_debug_tsrc,
  output [6:0]  io_rf_read_ports_0_addr,
  input  [63:0] io_rf_read_ports_0_data,
  output [6:0]  io_rf_read_ports_1_addr,
  input  [63:0] io_rf_read_ports_1_data,
  output [6:0]  io_rf_read_ports_2_addr,
  input  [63:0] io_rf_read_ports_2_data,
  output [6:0]  io_rf_read_ports_3_addr,
  input  [63:0] io_rf_read_ports_3_data,
  output [6:0]  io_rf_read_ports_4_addr,
  input  [63:0] io_rf_read_ports_4_data,
  output [6:0]  io_rf_read_ports_5_addr,
  input  [63:0] io_rf_read_ports_5_data,
  output [6:0]  io_rf_read_ports_6_addr,
  input  [63:0] io_rf_read_ports_6_data,
  output [6:0]  io_rf_read_ports_7_addr,
  input  [63:0] io_rf_read_ports_7_data,
  output [6:0]  io_rf_read_ports_8_addr,
  input  [63:0] io_rf_read_ports_8_data,
  output [4:0]  io_prf_read_ports_0_addr,
  input         io_prf_read_ports_0_data,
  output [4:0]  io_prf_read_ports_1_addr,
  input         io_prf_read_ports_1_data,
  output [4:0]  io_prf_read_ports_2_addr,
  input         io_prf_read_ports_2_data,
  output [6:0]  io_flag_rf_read_ports_0_addr,
  input  [3:0]  io_flag_rf_read_ports_0_data,
  output [6:0]  io_flag_rf_read_ports_1_addr,
  input  [3:0]  io_flag_rf_read_ports_1_data,
  output [6:0]  io_flag_rf_read_ports_2_addr,
  input  [3:0]  io_flag_rf_read_ports_2_data,
  input         io_bypass_0_valid,
  input         io_bypass_0_bits_uop_switch,
  input         io_bypass_0_bits_uop_switch_off,
  input         io_bypass_0_bits_uop_is_unicore,
  input  [2:0]  io_bypass_0_bits_uop_shift,
  input  [1:0]  io_bypass_0_bits_uop_lrs3_rtype,
  input         io_bypass_0_bits_uop_rflag,
  input         io_bypass_0_bits_uop_wflag,
  input  [3:0]  io_bypass_0_bits_uop_prflag,
  input  [3:0]  io_bypass_0_bits_uop_pwflag,
  input         io_bypass_0_bits_uop_pflag_busy,
  input  [3:0]  io_bypass_0_bits_uop_stale_pflag,
  input  [3:0]  io_bypass_0_bits_uop_op1_sel,
  input  [3:0]  io_bypass_0_bits_uop_op2_sel,
  input  [5:0]  io_bypass_0_bits_uop_split_num,
  input  [5:0]  io_bypass_0_bits_uop_self_index,
  input  [5:0]  io_bypass_0_bits_uop_rob_inst_idx,
  input  [5:0]  io_bypass_0_bits_uop_address_num,
  input  [6:0]  io_bypass_0_bits_uop_uopc,
  input  [31:0] io_bypass_0_bits_uop_inst,
  input  [31:0] io_bypass_0_bits_uop_debug_inst,
  input         io_bypass_0_bits_uop_is_rvc,
  input  [39:0] io_bypass_0_bits_uop_debug_pc,
  input  [2:0]  io_bypass_0_bits_uop_iq_type,
  input  [9:0]  io_bypass_0_bits_uop_fu_code,
  input  [3:0]  io_bypass_0_bits_uop_ctrl_br_type,
  input  [1:0]  io_bypass_0_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_bypass_0_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_bypass_0_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_bypass_0_bits_uop_ctrl_op_fcn,
  input         io_bypass_0_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_bypass_0_bits_uop_ctrl_csr_cmd,
  input         io_bypass_0_bits_uop_ctrl_is_load,
  input         io_bypass_0_bits_uop_ctrl_is_sta,
  input         io_bypass_0_bits_uop_ctrl_is_std,
  input  [1:0]  io_bypass_0_bits_uop_ctrl_op3_sel,
  input  [1:0]  io_bypass_0_bits_uop_iw_state,
  input         io_bypass_0_bits_uop_iw_p1_poisoned,
  input         io_bypass_0_bits_uop_iw_p2_poisoned,
  input         io_bypass_0_bits_uop_is_br,
  input         io_bypass_0_bits_uop_is_jalr,
  input         io_bypass_0_bits_uop_is_jal,
  input         io_bypass_0_bits_uop_is_sfb,
  input  [11:0] io_bypass_0_bits_uop_br_mask,
  input  [3:0]  io_bypass_0_bits_uop_br_tag,
  input  [4:0]  io_bypass_0_bits_uop_ftq_idx,
  input         io_bypass_0_bits_uop_edge_inst,
  input  [5:0]  io_bypass_0_bits_uop_pc_lob,
  input         io_bypass_0_bits_uop_taken,
  input  [19:0] io_bypass_0_bits_uop_imm_packed,
  input  [11:0] io_bypass_0_bits_uop_csr_addr,
  input  [5:0]  io_bypass_0_bits_uop_rob_idx,
  input  [4:0]  io_bypass_0_bits_uop_ldq_idx,
  input  [4:0]  io_bypass_0_bits_uop_stq_idx,
  input  [1:0]  io_bypass_0_bits_uop_rxq_idx,
  input  [6:0]  io_bypass_0_bits_uop_pdst,
  input  [6:0]  io_bypass_0_bits_uop_prs1,
  input  [6:0]  io_bypass_0_bits_uop_prs2,
  input  [6:0]  io_bypass_0_bits_uop_prs3,
  input  [4:0]  io_bypass_0_bits_uop_ppred,
  input         io_bypass_0_bits_uop_prs1_busy,
  input         io_bypass_0_bits_uop_prs2_busy,
  input         io_bypass_0_bits_uop_prs3_busy,
  input         io_bypass_0_bits_uop_ppred_busy,
  input  [6:0]  io_bypass_0_bits_uop_stale_pdst,
  input         io_bypass_0_bits_uop_exception,
  input  [63:0] io_bypass_0_bits_uop_exc_cause,
  input         io_bypass_0_bits_uop_bypassable,
  input  [4:0]  io_bypass_0_bits_uop_mem_cmd,
  input  [1:0]  io_bypass_0_bits_uop_mem_size,
  input         io_bypass_0_bits_uop_mem_signed,
  input         io_bypass_0_bits_uop_is_fence,
  input         io_bypass_0_bits_uop_is_fencei,
  input         io_bypass_0_bits_uop_is_amo,
  input         io_bypass_0_bits_uop_uses_ldq,
  input         io_bypass_0_bits_uop_uses_stq,
  input         io_bypass_0_bits_uop_is_sys_pc2epc,
  input         io_bypass_0_bits_uop_is_unique,
  input         io_bypass_0_bits_uop_flush_on_commit,
  input         io_bypass_0_bits_uop_ldst_is_rs1,
  input  [5:0]  io_bypass_0_bits_uop_ldst,
  input  [5:0]  io_bypass_0_bits_uop_lrs1,
  input  [5:0]  io_bypass_0_bits_uop_lrs2,
  input  [5:0]  io_bypass_0_bits_uop_lrs3,
  input         io_bypass_0_bits_uop_ldst_val,
  input  [1:0]  io_bypass_0_bits_uop_dst_rtype,
  input  [1:0]  io_bypass_0_bits_uop_lrs1_rtype,
  input  [1:0]  io_bypass_0_bits_uop_lrs2_rtype,
  input         io_bypass_0_bits_uop_frs3_en,
  input         io_bypass_0_bits_uop_fp_val,
  input         io_bypass_0_bits_uop_fp_single,
  input         io_bypass_0_bits_uop_xcpt_pf_if,
  input         io_bypass_0_bits_uop_xcpt_ae_if,
  input         io_bypass_0_bits_uop_xcpt_ma_if,
  input         io_bypass_0_bits_uop_bp_debug_if,
  input         io_bypass_0_bits_uop_bp_xcpt_if,
  input  [1:0]  io_bypass_0_bits_uop_debug_fsrc,
  input  [1:0]  io_bypass_0_bits_uop_debug_tsrc,
  input  [63:0] io_bypass_0_bits_data,
  input         io_bypass_0_bits_predicated,
  input         io_bypass_0_bits_fflags_valid,
  input         io_bypass_0_bits_fflags_bits_uop_switch,
  input         io_bypass_0_bits_fflags_bits_uop_switch_off,
  input         io_bypass_0_bits_fflags_bits_uop_is_unicore,
  input  [2:0]  io_bypass_0_bits_fflags_bits_uop_shift,
  input  [1:0]  io_bypass_0_bits_fflags_bits_uop_lrs3_rtype,
  input         io_bypass_0_bits_fflags_bits_uop_rflag,
  input         io_bypass_0_bits_fflags_bits_uop_wflag,
  input  [3:0]  io_bypass_0_bits_fflags_bits_uop_prflag,
  input  [3:0]  io_bypass_0_bits_fflags_bits_uop_pwflag,
  input         io_bypass_0_bits_fflags_bits_uop_pflag_busy,
  input  [3:0]  io_bypass_0_bits_fflags_bits_uop_stale_pflag,
  input  [3:0]  io_bypass_0_bits_fflags_bits_uop_op1_sel,
  input  [3:0]  io_bypass_0_bits_fflags_bits_uop_op2_sel,
  input  [5:0]  io_bypass_0_bits_fflags_bits_uop_split_num,
  input  [5:0]  io_bypass_0_bits_fflags_bits_uop_self_index,
  input  [5:0]  io_bypass_0_bits_fflags_bits_uop_rob_inst_idx,
  input  [5:0]  io_bypass_0_bits_fflags_bits_uop_address_num,
  input  [6:0]  io_bypass_0_bits_fflags_bits_uop_uopc,
  input  [31:0] io_bypass_0_bits_fflags_bits_uop_inst,
  input  [31:0] io_bypass_0_bits_fflags_bits_uop_debug_inst,
  input         io_bypass_0_bits_fflags_bits_uop_is_rvc,
  input  [39:0] io_bypass_0_bits_fflags_bits_uop_debug_pc,
  input  [2:0]  io_bypass_0_bits_fflags_bits_uop_iq_type,
  input  [9:0]  io_bypass_0_bits_fflags_bits_uop_fu_code,
  input  [3:0]  io_bypass_0_bits_fflags_bits_uop_ctrl_br_type,
  input  [1:0]  io_bypass_0_bits_fflags_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_bypass_0_bits_fflags_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_bypass_0_bits_fflags_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_bypass_0_bits_fflags_bits_uop_ctrl_op_fcn,
  input         io_bypass_0_bits_fflags_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_bypass_0_bits_fflags_bits_uop_ctrl_csr_cmd,
  input         io_bypass_0_bits_fflags_bits_uop_ctrl_is_load,
  input         io_bypass_0_bits_fflags_bits_uop_ctrl_is_sta,
  input         io_bypass_0_bits_fflags_bits_uop_ctrl_is_std,
  input  [1:0]  io_bypass_0_bits_fflags_bits_uop_ctrl_op3_sel,
  input  [1:0]  io_bypass_0_bits_fflags_bits_uop_iw_state,
  input         io_bypass_0_bits_fflags_bits_uop_iw_p1_poisoned,
  input         io_bypass_0_bits_fflags_bits_uop_iw_p2_poisoned,
  input         io_bypass_0_bits_fflags_bits_uop_is_br,
  input         io_bypass_0_bits_fflags_bits_uop_is_jalr,
  input         io_bypass_0_bits_fflags_bits_uop_is_jal,
  input         io_bypass_0_bits_fflags_bits_uop_is_sfb,
  input  [11:0] io_bypass_0_bits_fflags_bits_uop_br_mask,
  input  [3:0]  io_bypass_0_bits_fflags_bits_uop_br_tag,
  input  [4:0]  io_bypass_0_bits_fflags_bits_uop_ftq_idx,
  input         io_bypass_0_bits_fflags_bits_uop_edge_inst,
  input  [5:0]  io_bypass_0_bits_fflags_bits_uop_pc_lob,
  input         io_bypass_0_bits_fflags_bits_uop_taken,
  input  [19:0] io_bypass_0_bits_fflags_bits_uop_imm_packed,
  input  [11:0] io_bypass_0_bits_fflags_bits_uop_csr_addr,
  input  [5:0]  io_bypass_0_bits_fflags_bits_uop_rob_idx,
  input  [4:0]  io_bypass_0_bits_fflags_bits_uop_ldq_idx,
  input  [4:0]  io_bypass_0_bits_fflags_bits_uop_stq_idx,
  input  [1:0]  io_bypass_0_bits_fflags_bits_uop_rxq_idx,
  input  [6:0]  io_bypass_0_bits_fflags_bits_uop_pdst,
  input  [6:0]  io_bypass_0_bits_fflags_bits_uop_prs1,
  input  [6:0]  io_bypass_0_bits_fflags_bits_uop_prs2,
  input  [6:0]  io_bypass_0_bits_fflags_bits_uop_prs3,
  input  [4:0]  io_bypass_0_bits_fflags_bits_uop_ppred,
  input         io_bypass_0_bits_fflags_bits_uop_prs1_busy,
  input         io_bypass_0_bits_fflags_bits_uop_prs2_busy,
  input         io_bypass_0_bits_fflags_bits_uop_prs3_busy,
  input         io_bypass_0_bits_fflags_bits_uop_ppred_busy,
  input  [6:0]  io_bypass_0_bits_fflags_bits_uop_stale_pdst,
  input         io_bypass_0_bits_fflags_bits_uop_exception,
  input  [63:0] io_bypass_0_bits_fflags_bits_uop_exc_cause,
  input         io_bypass_0_bits_fflags_bits_uop_bypassable,
  input  [4:0]  io_bypass_0_bits_fflags_bits_uop_mem_cmd,
  input  [1:0]  io_bypass_0_bits_fflags_bits_uop_mem_size,
  input         io_bypass_0_bits_fflags_bits_uop_mem_signed,
  input         io_bypass_0_bits_fflags_bits_uop_is_fence,
  input         io_bypass_0_bits_fflags_bits_uop_is_fencei,
  input         io_bypass_0_bits_fflags_bits_uop_is_amo,
  input         io_bypass_0_bits_fflags_bits_uop_uses_ldq,
  input         io_bypass_0_bits_fflags_bits_uop_uses_stq,
  input         io_bypass_0_bits_fflags_bits_uop_is_sys_pc2epc,
  input         io_bypass_0_bits_fflags_bits_uop_is_unique,
  input         io_bypass_0_bits_fflags_bits_uop_flush_on_commit,
  input         io_bypass_0_bits_fflags_bits_uop_ldst_is_rs1,
  input  [5:0]  io_bypass_0_bits_fflags_bits_uop_ldst,
  input  [5:0]  io_bypass_0_bits_fflags_bits_uop_lrs1,
  input  [5:0]  io_bypass_0_bits_fflags_bits_uop_lrs2,
  input  [5:0]  io_bypass_0_bits_fflags_bits_uop_lrs3,
  input         io_bypass_0_bits_fflags_bits_uop_ldst_val,
  input  [1:0]  io_bypass_0_bits_fflags_bits_uop_dst_rtype,
  input  [1:0]  io_bypass_0_bits_fflags_bits_uop_lrs1_rtype,
  input  [1:0]  io_bypass_0_bits_fflags_bits_uop_lrs2_rtype,
  input         io_bypass_0_bits_fflags_bits_uop_frs3_en,
  input         io_bypass_0_bits_fflags_bits_uop_fp_val,
  input         io_bypass_0_bits_fflags_bits_uop_fp_single,
  input         io_bypass_0_bits_fflags_bits_uop_xcpt_pf_if,
  input         io_bypass_0_bits_fflags_bits_uop_xcpt_ae_if,
  input         io_bypass_0_bits_fflags_bits_uop_xcpt_ma_if,
  input         io_bypass_0_bits_fflags_bits_uop_bp_debug_if,
  input         io_bypass_0_bits_fflags_bits_uop_bp_xcpt_if,
  input  [1:0]  io_bypass_0_bits_fflags_bits_uop_debug_fsrc,
  input  [1:0]  io_bypass_0_bits_fflags_bits_uop_debug_tsrc,
  input  [4:0]  io_bypass_0_bits_fflags_bits_flags,
  input  [3:0]  io_bypass_0_bits_flagdata,
  input         io_bypass_0_bits_fflagdata_valid,
  input         io_bypass_0_bits_fflagdata_bits_uop_switch,
  input         io_bypass_0_bits_fflagdata_bits_uop_switch_off,
  input         io_bypass_0_bits_fflagdata_bits_uop_is_unicore,
  input  [2:0]  io_bypass_0_bits_fflagdata_bits_uop_shift,
  input  [1:0]  io_bypass_0_bits_fflagdata_bits_uop_lrs3_rtype,
  input         io_bypass_0_bits_fflagdata_bits_uop_rflag,
  input         io_bypass_0_bits_fflagdata_bits_uop_wflag,
  input  [3:0]  io_bypass_0_bits_fflagdata_bits_uop_prflag,
  input  [3:0]  io_bypass_0_bits_fflagdata_bits_uop_pwflag,
  input         io_bypass_0_bits_fflagdata_bits_uop_pflag_busy,
  input  [3:0]  io_bypass_0_bits_fflagdata_bits_uop_stale_pflag,
  input  [3:0]  io_bypass_0_bits_fflagdata_bits_uop_op1_sel,
  input  [3:0]  io_bypass_0_bits_fflagdata_bits_uop_op2_sel,
  input  [5:0]  io_bypass_0_bits_fflagdata_bits_uop_split_num,
  input  [5:0]  io_bypass_0_bits_fflagdata_bits_uop_self_index,
  input  [5:0]  io_bypass_0_bits_fflagdata_bits_uop_rob_inst_idx,
  input  [5:0]  io_bypass_0_bits_fflagdata_bits_uop_address_num,
  input  [6:0]  io_bypass_0_bits_fflagdata_bits_uop_uopc,
  input  [31:0] io_bypass_0_bits_fflagdata_bits_uop_inst,
  input  [31:0] io_bypass_0_bits_fflagdata_bits_uop_debug_inst,
  input         io_bypass_0_bits_fflagdata_bits_uop_is_rvc,
  input  [39:0] io_bypass_0_bits_fflagdata_bits_uop_debug_pc,
  input  [2:0]  io_bypass_0_bits_fflagdata_bits_uop_iq_type,
  input  [9:0]  io_bypass_0_bits_fflagdata_bits_uop_fu_code,
  input  [3:0]  io_bypass_0_bits_fflagdata_bits_uop_ctrl_br_type,
  input  [1:0]  io_bypass_0_bits_fflagdata_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_bypass_0_bits_fflagdata_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_bypass_0_bits_fflagdata_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_bypass_0_bits_fflagdata_bits_uop_ctrl_op_fcn,
  input         io_bypass_0_bits_fflagdata_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_bypass_0_bits_fflagdata_bits_uop_ctrl_csr_cmd,
  input         io_bypass_0_bits_fflagdata_bits_uop_ctrl_is_load,
  input         io_bypass_0_bits_fflagdata_bits_uop_ctrl_is_sta,
  input         io_bypass_0_bits_fflagdata_bits_uop_ctrl_is_std,
  input  [1:0]  io_bypass_0_bits_fflagdata_bits_uop_ctrl_op3_sel,
  input  [1:0]  io_bypass_0_bits_fflagdata_bits_uop_iw_state,
  input         io_bypass_0_bits_fflagdata_bits_uop_iw_p1_poisoned,
  input         io_bypass_0_bits_fflagdata_bits_uop_iw_p2_poisoned,
  input         io_bypass_0_bits_fflagdata_bits_uop_is_br,
  input         io_bypass_0_bits_fflagdata_bits_uop_is_jalr,
  input         io_bypass_0_bits_fflagdata_bits_uop_is_jal,
  input         io_bypass_0_bits_fflagdata_bits_uop_is_sfb,
  input  [11:0] io_bypass_0_bits_fflagdata_bits_uop_br_mask,
  input  [3:0]  io_bypass_0_bits_fflagdata_bits_uop_br_tag,
  input  [4:0]  io_bypass_0_bits_fflagdata_bits_uop_ftq_idx,
  input         io_bypass_0_bits_fflagdata_bits_uop_edge_inst,
  input  [5:0]  io_bypass_0_bits_fflagdata_bits_uop_pc_lob,
  input         io_bypass_0_bits_fflagdata_bits_uop_taken,
  input  [19:0] io_bypass_0_bits_fflagdata_bits_uop_imm_packed,
  input  [11:0] io_bypass_0_bits_fflagdata_bits_uop_csr_addr,
  input  [5:0]  io_bypass_0_bits_fflagdata_bits_uop_rob_idx,
  input  [4:0]  io_bypass_0_bits_fflagdata_bits_uop_ldq_idx,
  input  [4:0]  io_bypass_0_bits_fflagdata_bits_uop_stq_idx,
  input  [1:0]  io_bypass_0_bits_fflagdata_bits_uop_rxq_idx,
  input  [6:0]  io_bypass_0_bits_fflagdata_bits_uop_pdst,
  input  [6:0]  io_bypass_0_bits_fflagdata_bits_uop_prs1,
  input  [6:0]  io_bypass_0_bits_fflagdata_bits_uop_prs2,
  input  [6:0]  io_bypass_0_bits_fflagdata_bits_uop_prs3,
  input  [4:0]  io_bypass_0_bits_fflagdata_bits_uop_ppred,
  input         io_bypass_0_bits_fflagdata_bits_uop_prs1_busy,
  input         io_bypass_0_bits_fflagdata_bits_uop_prs2_busy,
  input         io_bypass_0_bits_fflagdata_bits_uop_prs3_busy,
  input         io_bypass_0_bits_fflagdata_bits_uop_ppred_busy,
  input  [6:0]  io_bypass_0_bits_fflagdata_bits_uop_stale_pdst,
  input         io_bypass_0_bits_fflagdata_bits_uop_exception,
  input  [63:0] io_bypass_0_bits_fflagdata_bits_uop_exc_cause,
  input         io_bypass_0_bits_fflagdata_bits_uop_bypassable,
  input  [4:0]  io_bypass_0_bits_fflagdata_bits_uop_mem_cmd,
  input  [1:0]  io_bypass_0_bits_fflagdata_bits_uop_mem_size,
  input         io_bypass_0_bits_fflagdata_bits_uop_mem_signed,
  input         io_bypass_0_bits_fflagdata_bits_uop_is_fence,
  input         io_bypass_0_bits_fflagdata_bits_uop_is_fencei,
  input         io_bypass_0_bits_fflagdata_bits_uop_is_amo,
  input         io_bypass_0_bits_fflagdata_bits_uop_uses_ldq,
  input         io_bypass_0_bits_fflagdata_bits_uop_uses_stq,
  input         io_bypass_0_bits_fflagdata_bits_uop_is_sys_pc2epc,
  input         io_bypass_0_bits_fflagdata_bits_uop_is_unique,
  input         io_bypass_0_bits_fflagdata_bits_uop_flush_on_commit,
  input         io_bypass_0_bits_fflagdata_bits_uop_ldst_is_rs1,
  input  [5:0]  io_bypass_0_bits_fflagdata_bits_uop_ldst,
  input  [5:0]  io_bypass_0_bits_fflagdata_bits_uop_lrs1,
  input  [5:0]  io_bypass_0_bits_fflagdata_bits_uop_lrs2,
  input  [5:0]  io_bypass_0_bits_fflagdata_bits_uop_lrs3,
  input         io_bypass_0_bits_fflagdata_bits_uop_ldst_val,
  input  [1:0]  io_bypass_0_bits_fflagdata_bits_uop_dst_rtype,
  input  [1:0]  io_bypass_0_bits_fflagdata_bits_uop_lrs1_rtype,
  input  [1:0]  io_bypass_0_bits_fflagdata_bits_uop_lrs2_rtype,
  input         io_bypass_0_bits_fflagdata_bits_uop_frs3_en,
  input         io_bypass_0_bits_fflagdata_bits_uop_fp_val,
  input         io_bypass_0_bits_fflagdata_bits_uop_fp_single,
  input         io_bypass_0_bits_fflagdata_bits_uop_xcpt_pf_if,
  input         io_bypass_0_bits_fflagdata_bits_uop_xcpt_ae_if,
  input         io_bypass_0_bits_fflagdata_bits_uop_xcpt_ma_if,
  input         io_bypass_0_bits_fflagdata_bits_uop_bp_debug_if,
  input         io_bypass_0_bits_fflagdata_bits_uop_bp_xcpt_if,
  input  [1:0]  io_bypass_0_bits_fflagdata_bits_uop_debug_fsrc,
  input  [1:0]  io_bypass_0_bits_fflagdata_bits_uop_debug_tsrc,
  input  [31:0] io_bypass_0_bits_fflagdata_bits_fflag,
  input         io_bypass_1_valid,
  input         io_bypass_1_bits_uop_switch,
  input         io_bypass_1_bits_uop_switch_off,
  input         io_bypass_1_bits_uop_is_unicore,
  input  [2:0]  io_bypass_1_bits_uop_shift,
  input  [1:0]  io_bypass_1_bits_uop_lrs3_rtype,
  input         io_bypass_1_bits_uop_rflag,
  input         io_bypass_1_bits_uop_wflag,
  input  [3:0]  io_bypass_1_bits_uop_prflag,
  input  [3:0]  io_bypass_1_bits_uop_pwflag,
  input         io_bypass_1_bits_uop_pflag_busy,
  input  [3:0]  io_bypass_1_bits_uop_stale_pflag,
  input  [3:0]  io_bypass_1_bits_uop_op1_sel,
  input  [3:0]  io_bypass_1_bits_uop_op2_sel,
  input  [5:0]  io_bypass_1_bits_uop_split_num,
  input  [5:0]  io_bypass_1_bits_uop_self_index,
  input  [5:0]  io_bypass_1_bits_uop_rob_inst_idx,
  input  [5:0]  io_bypass_1_bits_uop_address_num,
  input  [6:0]  io_bypass_1_bits_uop_uopc,
  input  [31:0] io_bypass_1_bits_uop_inst,
  input  [31:0] io_bypass_1_bits_uop_debug_inst,
  input         io_bypass_1_bits_uop_is_rvc,
  input  [39:0] io_bypass_1_bits_uop_debug_pc,
  input  [2:0]  io_bypass_1_bits_uop_iq_type,
  input  [9:0]  io_bypass_1_bits_uop_fu_code,
  input  [3:0]  io_bypass_1_bits_uop_ctrl_br_type,
  input  [1:0]  io_bypass_1_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_bypass_1_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_bypass_1_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_bypass_1_bits_uop_ctrl_op_fcn,
  input         io_bypass_1_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_bypass_1_bits_uop_ctrl_csr_cmd,
  input         io_bypass_1_bits_uop_ctrl_is_load,
  input         io_bypass_1_bits_uop_ctrl_is_sta,
  input         io_bypass_1_bits_uop_ctrl_is_std,
  input  [1:0]  io_bypass_1_bits_uop_ctrl_op3_sel,
  input  [1:0]  io_bypass_1_bits_uop_iw_state,
  input         io_bypass_1_bits_uop_iw_p1_poisoned,
  input         io_bypass_1_bits_uop_iw_p2_poisoned,
  input         io_bypass_1_bits_uop_is_br,
  input         io_bypass_1_bits_uop_is_jalr,
  input         io_bypass_1_bits_uop_is_jal,
  input         io_bypass_1_bits_uop_is_sfb,
  input  [11:0] io_bypass_1_bits_uop_br_mask,
  input  [3:0]  io_bypass_1_bits_uop_br_tag,
  input  [4:0]  io_bypass_1_bits_uop_ftq_idx,
  input         io_bypass_1_bits_uop_edge_inst,
  input  [5:0]  io_bypass_1_bits_uop_pc_lob,
  input         io_bypass_1_bits_uop_taken,
  input  [19:0] io_bypass_1_bits_uop_imm_packed,
  input  [11:0] io_bypass_1_bits_uop_csr_addr,
  input  [5:0]  io_bypass_1_bits_uop_rob_idx,
  input  [4:0]  io_bypass_1_bits_uop_ldq_idx,
  input  [4:0]  io_bypass_1_bits_uop_stq_idx,
  input  [1:0]  io_bypass_1_bits_uop_rxq_idx,
  input  [6:0]  io_bypass_1_bits_uop_pdst,
  input  [6:0]  io_bypass_1_bits_uop_prs1,
  input  [6:0]  io_bypass_1_bits_uop_prs2,
  input  [6:0]  io_bypass_1_bits_uop_prs3,
  input  [4:0]  io_bypass_1_bits_uop_ppred,
  input         io_bypass_1_bits_uop_prs1_busy,
  input         io_bypass_1_bits_uop_prs2_busy,
  input         io_bypass_1_bits_uop_prs3_busy,
  input         io_bypass_1_bits_uop_ppred_busy,
  input  [6:0]  io_bypass_1_bits_uop_stale_pdst,
  input         io_bypass_1_bits_uop_exception,
  input  [63:0] io_bypass_1_bits_uop_exc_cause,
  input         io_bypass_1_bits_uop_bypassable,
  input  [4:0]  io_bypass_1_bits_uop_mem_cmd,
  input  [1:0]  io_bypass_1_bits_uop_mem_size,
  input         io_bypass_1_bits_uop_mem_signed,
  input         io_bypass_1_bits_uop_is_fence,
  input         io_bypass_1_bits_uop_is_fencei,
  input         io_bypass_1_bits_uop_is_amo,
  input         io_bypass_1_bits_uop_uses_ldq,
  input         io_bypass_1_bits_uop_uses_stq,
  input         io_bypass_1_bits_uop_is_sys_pc2epc,
  input         io_bypass_1_bits_uop_is_unique,
  input         io_bypass_1_bits_uop_flush_on_commit,
  input         io_bypass_1_bits_uop_ldst_is_rs1,
  input  [5:0]  io_bypass_1_bits_uop_ldst,
  input  [5:0]  io_bypass_1_bits_uop_lrs1,
  input  [5:0]  io_bypass_1_bits_uop_lrs2,
  input  [5:0]  io_bypass_1_bits_uop_lrs3,
  input         io_bypass_1_bits_uop_ldst_val,
  input  [1:0]  io_bypass_1_bits_uop_dst_rtype,
  input  [1:0]  io_bypass_1_bits_uop_lrs1_rtype,
  input  [1:0]  io_bypass_1_bits_uop_lrs2_rtype,
  input         io_bypass_1_bits_uop_frs3_en,
  input         io_bypass_1_bits_uop_fp_val,
  input         io_bypass_1_bits_uop_fp_single,
  input         io_bypass_1_bits_uop_xcpt_pf_if,
  input         io_bypass_1_bits_uop_xcpt_ae_if,
  input         io_bypass_1_bits_uop_xcpt_ma_if,
  input         io_bypass_1_bits_uop_bp_debug_if,
  input         io_bypass_1_bits_uop_bp_xcpt_if,
  input  [1:0]  io_bypass_1_bits_uop_debug_fsrc,
  input  [1:0]  io_bypass_1_bits_uop_debug_tsrc,
  input  [63:0] io_bypass_1_bits_data,
  input         io_bypass_1_bits_predicated,
  input         io_bypass_1_bits_fflags_valid,
  input         io_bypass_1_bits_fflags_bits_uop_switch,
  input         io_bypass_1_bits_fflags_bits_uop_switch_off,
  input         io_bypass_1_bits_fflags_bits_uop_is_unicore,
  input  [2:0]  io_bypass_1_bits_fflags_bits_uop_shift,
  input  [1:0]  io_bypass_1_bits_fflags_bits_uop_lrs3_rtype,
  input         io_bypass_1_bits_fflags_bits_uop_rflag,
  input         io_bypass_1_bits_fflags_bits_uop_wflag,
  input  [3:0]  io_bypass_1_bits_fflags_bits_uop_prflag,
  input  [3:0]  io_bypass_1_bits_fflags_bits_uop_pwflag,
  input         io_bypass_1_bits_fflags_bits_uop_pflag_busy,
  input  [3:0]  io_bypass_1_bits_fflags_bits_uop_stale_pflag,
  input  [3:0]  io_bypass_1_bits_fflags_bits_uop_op1_sel,
  input  [3:0]  io_bypass_1_bits_fflags_bits_uop_op2_sel,
  input  [5:0]  io_bypass_1_bits_fflags_bits_uop_split_num,
  input  [5:0]  io_bypass_1_bits_fflags_bits_uop_self_index,
  input  [5:0]  io_bypass_1_bits_fflags_bits_uop_rob_inst_idx,
  input  [5:0]  io_bypass_1_bits_fflags_bits_uop_address_num,
  input  [6:0]  io_bypass_1_bits_fflags_bits_uop_uopc,
  input  [31:0] io_bypass_1_bits_fflags_bits_uop_inst,
  input  [31:0] io_bypass_1_bits_fflags_bits_uop_debug_inst,
  input         io_bypass_1_bits_fflags_bits_uop_is_rvc,
  input  [39:0] io_bypass_1_bits_fflags_bits_uop_debug_pc,
  input  [2:0]  io_bypass_1_bits_fflags_bits_uop_iq_type,
  input  [9:0]  io_bypass_1_bits_fflags_bits_uop_fu_code,
  input  [3:0]  io_bypass_1_bits_fflags_bits_uop_ctrl_br_type,
  input  [1:0]  io_bypass_1_bits_fflags_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_bypass_1_bits_fflags_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_bypass_1_bits_fflags_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_bypass_1_bits_fflags_bits_uop_ctrl_op_fcn,
  input         io_bypass_1_bits_fflags_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_bypass_1_bits_fflags_bits_uop_ctrl_csr_cmd,
  input         io_bypass_1_bits_fflags_bits_uop_ctrl_is_load,
  input         io_bypass_1_bits_fflags_bits_uop_ctrl_is_sta,
  input         io_bypass_1_bits_fflags_bits_uop_ctrl_is_std,
  input  [1:0]  io_bypass_1_bits_fflags_bits_uop_ctrl_op3_sel,
  input  [1:0]  io_bypass_1_bits_fflags_bits_uop_iw_state,
  input         io_bypass_1_bits_fflags_bits_uop_iw_p1_poisoned,
  input         io_bypass_1_bits_fflags_bits_uop_iw_p2_poisoned,
  input         io_bypass_1_bits_fflags_bits_uop_is_br,
  input         io_bypass_1_bits_fflags_bits_uop_is_jalr,
  input         io_bypass_1_bits_fflags_bits_uop_is_jal,
  input         io_bypass_1_bits_fflags_bits_uop_is_sfb,
  input  [11:0] io_bypass_1_bits_fflags_bits_uop_br_mask,
  input  [3:0]  io_bypass_1_bits_fflags_bits_uop_br_tag,
  input  [4:0]  io_bypass_1_bits_fflags_bits_uop_ftq_idx,
  input         io_bypass_1_bits_fflags_bits_uop_edge_inst,
  input  [5:0]  io_bypass_1_bits_fflags_bits_uop_pc_lob,
  input         io_bypass_1_bits_fflags_bits_uop_taken,
  input  [19:0] io_bypass_1_bits_fflags_bits_uop_imm_packed,
  input  [11:0] io_bypass_1_bits_fflags_bits_uop_csr_addr,
  input  [5:0]  io_bypass_1_bits_fflags_bits_uop_rob_idx,
  input  [4:0]  io_bypass_1_bits_fflags_bits_uop_ldq_idx,
  input  [4:0]  io_bypass_1_bits_fflags_bits_uop_stq_idx,
  input  [1:0]  io_bypass_1_bits_fflags_bits_uop_rxq_idx,
  input  [6:0]  io_bypass_1_bits_fflags_bits_uop_pdst,
  input  [6:0]  io_bypass_1_bits_fflags_bits_uop_prs1,
  input  [6:0]  io_bypass_1_bits_fflags_bits_uop_prs2,
  input  [6:0]  io_bypass_1_bits_fflags_bits_uop_prs3,
  input  [4:0]  io_bypass_1_bits_fflags_bits_uop_ppred,
  input         io_bypass_1_bits_fflags_bits_uop_prs1_busy,
  input         io_bypass_1_bits_fflags_bits_uop_prs2_busy,
  input         io_bypass_1_bits_fflags_bits_uop_prs3_busy,
  input         io_bypass_1_bits_fflags_bits_uop_ppred_busy,
  input  [6:0]  io_bypass_1_bits_fflags_bits_uop_stale_pdst,
  input         io_bypass_1_bits_fflags_bits_uop_exception,
  input  [63:0] io_bypass_1_bits_fflags_bits_uop_exc_cause,
  input         io_bypass_1_bits_fflags_bits_uop_bypassable,
  input  [4:0]  io_bypass_1_bits_fflags_bits_uop_mem_cmd,
  input  [1:0]  io_bypass_1_bits_fflags_bits_uop_mem_size,
  input         io_bypass_1_bits_fflags_bits_uop_mem_signed,
  input         io_bypass_1_bits_fflags_bits_uop_is_fence,
  input         io_bypass_1_bits_fflags_bits_uop_is_fencei,
  input         io_bypass_1_bits_fflags_bits_uop_is_amo,
  input         io_bypass_1_bits_fflags_bits_uop_uses_ldq,
  input         io_bypass_1_bits_fflags_bits_uop_uses_stq,
  input         io_bypass_1_bits_fflags_bits_uop_is_sys_pc2epc,
  input         io_bypass_1_bits_fflags_bits_uop_is_unique,
  input         io_bypass_1_bits_fflags_bits_uop_flush_on_commit,
  input         io_bypass_1_bits_fflags_bits_uop_ldst_is_rs1,
  input  [5:0]  io_bypass_1_bits_fflags_bits_uop_ldst,
  input  [5:0]  io_bypass_1_bits_fflags_bits_uop_lrs1,
  input  [5:0]  io_bypass_1_bits_fflags_bits_uop_lrs2,
  input  [5:0]  io_bypass_1_bits_fflags_bits_uop_lrs3,
  input         io_bypass_1_bits_fflags_bits_uop_ldst_val,
  input  [1:0]  io_bypass_1_bits_fflags_bits_uop_dst_rtype,
  input  [1:0]  io_bypass_1_bits_fflags_bits_uop_lrs1_rtype,
  input  [1:0]  io_bypass_1_bits_fflags_bits_uop_lrs2_rtype,
  input         io_bypass_1_bits_fflags_bits_uop_frs3_en,
  input         io_bypass_1_bits_fflags_bits_uop_fp_val,
  input         io_bypass_1_bits_fflags_bits_uop_fp_single,
  input         io_bypass_1_bits_fflags_bits_uop_xcpt_pf_if,
  input         io_bypass_1_bits_fflags_bits_uop_xcpt_ae_if,
  input         io_bypass_1_bits_fflags_bits_uop_xcpt_ma_if,
  input         io_bypass_1_bits_fflags_bits_uop_bp_debug_if,
  input         io_bypass_1_bits_fflags_bits_uop_bp_xcpt_if,
  input  [1:0]  io_bypass_1_bits_fflags_bits_uop_debug_fsrc,
  input  [1:0]  io_bypass_1_bits_fflags_bits_uop_debug_tsrc,
  input  [4:0]  io_bypass_1_bits_fflags_bits_flags,
  input  [3:0]  io_bypass_1_bits_flagdata,
  input         io_bypass_1_bits_fflagdata_valid,
  input         io_bypass_1_bits_fflagdata_bits_uop_switch,
  input         io_bypass_1_bits_fflagdata_bits_uop_switch_off,
  input         io_bypass_1_bits_fflagdata_bits_uop_is_unicore,
  input  [2:0]  io_bypass_1_bits_fflagdata_bits_uop_shift,
  input  [1:0]  io_bypass_1_bits_fflagdata_bits_uop_lrs3_rtype,
  input         io_bypass_1_bits_fflagdata_bits_uop_rflag,
  input         io_bypass_1_bits_fflagdata_bits_uop_wflag,
  input  [3:0]  io_bypass_1_bits_fflagdata_bits_uop_prflag,
  input  [3:0]  io_bypass_1_bits_fflagdata_bits_uop_pwflag,
  input         io_bypass_1_bits_fflagdata_bits_uop_pflag_busy,
  input  [3:0]  io_bypass_1_bits_fflagdata_bits_uop_stale_pflag,
  input  [3:0]  io_bypass_1_bits_fflagdata_bits_uop_op1_sel,
  input  [3:0]  io_bypass_1_bits_fflagdata_bits_uop_op2_sel,
  input  [5:0]  io_bypass_1_bits_fflagdata_bits_uop_split_num,
  input  [5:0]  io_bypass_1_bits_fflagdata_bits_uop_self_index,
  input  [5:0]  io_bypass_1_bits_fflagdata_bits_uop_rob_inst_idx,
  input  [5:0]  io_bypass_1_bits_fflagdata_bits_uop_address_num,
  input  [6:0]  io_bypass_1_bits_fflagdata_bits_uop_uopc,
  input  [31:0] io_bypass_1_bits_fflagdata_bits_uop_inst,
  input  [31:0] io_bypass_1_bits_fflagdata_bits_uop_debug_inst,
  input         io_bypass_1_bits_fflagdata_bits_uop_is_rvc,
  input  [39:0] io_bypass_1_bits_fflagdata_bits_uop_debug_pc,
  input  [2:0]  io_bypass_1_bits_fflagdata_bits_uop_iq_type,
  input  [9:0]  io_bypass_1_bits_fflagdata_bits_uop_fu_code,
  input  [3:0]  io_bypass_1_bits_fflagdata_bits_uop_ctrl_br_type,
  input  [1:0]  io_bypass_1_bits_fflagdata_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_bypass_1_bits_fflagdata_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_bypass_1_bits_fflagdata_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_bypass_1_bits_fflagdata_bits_uop_ctrl_op_fcn,
  input         io_bypass_1_bits_fflagdata_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_bypass_1_bits_fflagdata_bits_uop_ctrl_csr_cmd,
  input         io_bypass_1_bits_fflagdata_bits_uop_ctrl_is_load,
  input         io_bypass_1_bits_fflagdata_bits_uop_ctrl_is_sta,
  input         io_bypass_1_bits_fflagdata_bits_uop_ctrl_is_std,
  input  [1:0]  io_bypass_1_bits_fflagdata_bits_uop_ctrl_op3_sel,
  input  [1:0]  io_bypass_1_bits_fflagdata_bits_uop_iw_state,
  input         io_bypass_1_bits_fflagdata_bits_uop_iw_p1_poisoned,
  input         io_bypass_1_bits_fflagdata_bits_uop_iw_p2_poisoned,
  input         io_bypass_1_bits_fflagdata_bits_uop_is_br,
  input         io_bypass_1_bits_fflagdata_bits_uop_is_jalr,
  input         io_bypass_1_bits_fflagdata_bits_uop_is_jal,
  input         io_bypass_1_bits_fflagdata_bits_uop_is_sfb,
  input  [11:0] io_bypass_1_bits_fflagdata_bits_uop_br_mask,
  input  [3:0]  io_bypass_1_bits_fflagdata_bits_uop_br_tag,
  input  [4:0]  io_bypass_1_bits_fflagdata_bits_uop_ftq_idx,
  input         io_bypass_1_bits_fflagdata_bits_uop_edge_inst,
  input  [5:0]  io_bypass_1_bits_fflagdata_bits_uop_pc_lob,
  input         io_bypass_1_bits_fflagdata_bits_uop_taken,
  input  [19:0] io_bypass_1_bits_fflagdata_bits_uop_imm_packed,
  input  [11:0] io_bypass_1_bits_fflagdata_bits_uop_csr_addr,
  input  [5:0]  io_bypass_1_bits_fflagdata_bits_uop_rob_idx,
  input  [4:0]  io_bypass_1_bits_fflagdata_bits_uop_ldq_idx,
  input  [4:0]  io_bypass_1_bits_fflagdata_bits_uop_stq_idx,
  input  [1:0]  io_bypass_1_bits_fflagdata_bits_uop_rxq_idx,
  input  [6:0]  io_bypass_1_bits_fflagdata_bits_uop_pdst,
  input  [6:0]  io_bypass_1_bits_fflagdata_bits_uop_prs1,
  input  [6:0]  io_bypass_1_bits_fflagdata_bits_uop_prs2,
  input  [6:0]  io_bypass_1_bits_fflagdata_bits_uop_prs3,
  input  [4:0]  io_bypass_1_bits_fflagdata_bits_uop_ppred,
  input         io_bypass_1_bits_fflagdata_bits_uop_prs1_busy,
  input         io_bypass_1_bits_fflagdata_bits_uop_prs2_busy,
  input         io_bypass_1_bits_fflagdata_bits_uop_prs3_busy,
  input         io_bypass_1_bits_fflagdata_bits_uop_ppred_busy,
  input  [6:0]  io_bypass_1_bits_fflagdata_bits_uop_stale_pdst,
  input         io_bypass_1_bits_fflagdata_bits_uop_exception,
  input  [63:0] io_bypass_1_bits_fflagdata_bits_uop_exc_cause,
  input         io_bypass_1_bits_fflagdata_bits_uop_bypassable,
  input  [4:0]  io_bypass_1_bits_fflagdata_bits_uop_mem_cmd,
  input  [1:0]  io_bypass_1_bits_fflagdata_bits_uop_mem_size,
  input         io_bypass_1_bits_fflagdata_bits_uop_mem_signed,
  input         io_bypass_1_bits_fflagdata_bits_uop_is_fence,
  input         io_bypass_1_bits_fflagdata_bits_uop_is_fencei,
  input         io_bypass_1_bits_fflagdata_bits_uop_is_amo,
  input         io_bypass_1_bits_fflagdata_bits_uop_uses_ldq,
  input         io_bypass_1_bits_fflagdata_bits_uop_uses_stq,
  input         io_bypass_1_bits_fflagdata_bits_uop_is_sys_pc2epc,
  input         io_bypass_1_bits_fflagdata_bits_uop_is_unique,
  input         io_bypass_1_bits_fflagdata_bits_uop_flush_on_commit,
  input         io_bypass_1_bits_fflagdata_bits_uop_ldst_is_rs1,
  input  [5:0]  io_bypass_1_bits_fflagdata_bits_uop_ldst,
  input  [5:0]  io_bypass_1_bits_fflagdata_bits_uop_lrs1,
  input  [5:0]  io_bypass_1_bits_fflagdata_bits_uop_lrs2,
  input  [5:0]  io_bypass_1_bits_fflagdata_bits_uop_lrs3,
  input         io_bypass_1_bits_fflagdata_bits_uop_ldst_val,
  input  [1:0]  io_bypass_1_bits_fflagdata_bits_uop_dst_rtype,
  input  [1:0]  io_bypass_1_bits_fflagdata_bits_uop_lrs1_rtype,
  input  [1:0]  io_bypass_1_bits_fflagdata_bits_uop_lrs2_rtype,
  input         io_bypass_1_bits_fflagdata_bits_uop_frs3_en,
  input         io_bypass_1_bits_fflagdata_bits_uop_fp_val,
  input         io_bypass_1_bits_fflagdata_bits_uop_fp_single,
  input         io_bypass_1_bits_fflagdata_bits_uop_xcpt_pf_if,
  input         io_bypass_1_bits_fflagdata_bits_uop_xcpt_ae_if,
  input         io_bypass_1_bits_fflagdata_bits_uop_xcpt_ma_if,
  input         io_bypass_1_bits_fflagdata_bits_uop_bp_debug_if,
  input         io_bypass_1_bits_fflagdata_bits_uop_bp_xcpt_if,
  input  [1:0]  io_bypass_1_bits_fflagdata_bits_uop_debug_fsrc,
  input  [1:0]  io_bypass_1_bits_fflagdata_bits_uop_debug_tsrc,
  input  [31:0] io_bypass_1_bits_fflagdata_bits_fflag,
  input         io_bypass_2_valid,
  input         io_bypass_2_bits_uop_switch,
  input         io_bypass_2_bits_uop_switch_off,
  input         io_bypass_2_bits_uop_is_unicore,
  input  [2:0]  io_bypass_2_bits_uop_shift,
  input  [1:0]  io_bypass_2_bits_uop_lrs3_rtype,
  input         io_bypass_2_bits_uop_rflag,
  input         io_bypass_2_bits_uop_wflag,
  input  [3:0]  io_bypass_2_bits_uop_prflag,
  input  [3:0]  io_bypass_2_bits_uop_pwflag,
  input         io_bypass_2_bits_uop_pflag_busy,
  input  [3:0]  io_bypass_2_bits_uop_stale_pflag,
  input  [3:0]  io_bypass_2_bits_uop_op1_sel,
  input  [3:0]  io_bypass_2_bits_uop_op2_sel,
  input  [5:0]  io_bypass_2_bits_uop_split_num,
  input  [5:0]  io_bypass_2_bits_uop_self_index,
  input  [5:0]  io_bypass_2_bits_uop_rob_inst_idx,
  input  [5:0]  io_bypass_2_bits_uop_address_num,
  input  [6:0]  io_bypass_2_bits_uop_uopc,
  input  [31:0] io_bypass_2_bits_uop_inst,
  input  [31:0] io_bypass_2_bits_uop_debug_inst,
  input         io_bypass_2_bits_uop_is_rvc,
  input  [39:0] io_bypass_2_bits_uop_debug_pc,
  input  [2:0]  io_bypass_2_bits_uop_iq_type,
  input  [9:0]  io_bypass_2_bits_uop_fu_code,
  input  [3:0]  io_bypass_2_bits_uop_ctrl_br_type,
  input  [1:0]  io_bypass_2_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_bypass_2_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_bypass_2_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_bypass_2_bits_uop_ctrl_op_fcn,
  input         io_bypass_2_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_bypass_2_bits_uop_ctrl_csr_cmd,
  input         io_bypass_2_bits_uop_ctrl_is_load,
  input         io_bypass_2_bits_uop_ctrl_is_sta,
  input         io_bypass_2_bits_uop_ctrl_is_std,
  input  [1:0]  io_bypass_2_bits_uop_ctrl_op3_sel,
  input  [1:0]  io_bypass_2_bits_uop_iw_state,
  input         io_bypass_2_bits_uop_iw_p1_poisoned,
  input         io_bypass_2_bits_uop_iw_p2_poisoned,
  input         io_bypass_2_bits_uop_is_br,
  input         io_bypass_2_bits_uop_is_jalr,
  input         io_bypass_2_bits_uop_is_jal,
  input         io_bypass_2_bits_uop_is_sfb,
  input  [11:0] io_bypass_2_bits_uop_br_mask,
  input  [3:0]  io_bypass_2_bits_uop_br_tag,
  input  [4:0]  io_bypass_2_bits_uop_ftq_idx,
  input         io_bypass_2_bits_uop_edge_inst,
  input  [5:0]  io_bypass_2_bits_uop_pc_lob,
  input         io_bypass_2_bits_uop_taken,
  input  [19:0] io_bypass_2_bits_uop_imm_packed,
  input  [11:0] io_bypass_2_bits_uop_csr_addr,
  input  [5:0]  io_bypass_2_bits_uop_rob_idx,
  input  [4:0]  io_bypass_2_bits_uop_ldq_idx,
  input  [4:0]  io_bypass_2_bits_uop_stq_idx,
  input  [1:0]  io_bypass_2_bits_uop_rxq_idx,
  input  [6:0]  io_bypass_2_bits_uop_pdst,
  input  [6:0]  io_bypass_2_bits_uop_prs1,
  input  [6:0]  io_bypass_2_bits_uop_prs2,
  input  [6:0]  io_bypass_2_bits_uop_prs3,
  input  [4:0]  io_bypass_2_bits_uop_ppred,
  input         io_bypass_2_bits_uop_prs1_busy,
  input         io_bypass_2_bits_uop_prs2_busy,
  input         io_bypass_2_bits_uop_prs3_busy,
  input         io_bypass_2_bits_uop_ppred_busy,
  input  [6:0]  io_bypass_2_bits_uop_stale_pdst,
  input         io_bypass_2_bits_uop_exception,
  input  [63:0] io_bypass_2_bits_uop_exc_cause,
  input         io_bypass_2_bits_uop_bypassable,
  input  [4:0]  io_bypass_2_bits_uop_mem_cmd,
  input  [1:0]  io_bypass_2_bits_uop_mem_size,
  input         io_bypass_2_bits_uop_mem_signed,
  input         io_bypass_2_bits_uop_is_fence,
  input         io_bypass_2_bits_uop_is_fencei,
  input         io_bypass_2_bits_uop_is_amo,
  input         io_bypass_2_bits_uop_uses_ldq,
  input         io_bypass_2_bits_uop_uses_stq,
  input         io_bypass_2_bits_uop_is_sys_pc2epc,
  input         io_bypass_2_bits_uop_is_unique,
  input         io_bypass_2_bits_uop_flush_on_commit,
  input         io_bypass_2_bits_uop_ldst_is_rs1,
  input  [5:0]  io_bypass_2_bits_uop_ldst,
  input  [5:0]  io_bypass_2_bits_uop_lrs1,
  input  [5:0]  io_bypass_2_bits_uop_lrs2,
  input  [5:0]  io_bypass_2_bits_uop_lrs3,
  input         io_bypass_2_bits_uop_ldst_val,
  input  [1:0]  io_bypass_2_bits_uop_dst_rtype,
  input  [1:0]  io_bypass_2_bits_uop_lrs1_rtype,
  input  [1:0]  io_bypass_2_bits_uop_lrs2_rtype,
  input         io_bypass_2_bits_uop_frs3_en,
  input         io_bypass_2_bits_uop_fp_val,
  input         io_bypass_2_bits_uop_fp_single,
  input         io_bypass_2_bits_uop_xcpt_pf_if,
  input         io_bypass_2_bits_uop_xcpt_ae_if,
  input         io_bypass_2_bits_uop_xcpt_ma_if,
  input         io_bypass_2_bits_uop_bp_debug_if,
  input         io_bypass_2_bits_uop_bp_xcpt_if,
  input  [1:0]  io_bypass_2_bits_uop_debug_fsrc,
  input  [1:0]  io_bypass_2_bits_uop_debug_tsrc,
  input  [63:0] io_bypass_2_bits_data,
  input         io_bypass_2_bits_predicated,
  input         io_bypass_2_bits_fflags_valid,
  input         io_bypass_2_bits_fflags_bits_uop_switch,
  input         io_bypass_2_bits_fflags_bits_uop_switch_off,
  input         io_bypass_2_bits_fflags_bits_uop_is_unicore,
  input  [2:0]  io_bypass_2_bits_fflags_bits_uop_shift,
  input  [1:0]  io_bypass_2_bits_fflags_bits_uop_lrs3_rtype,
  input         io_bypass_2_bits_fflags_bits_uop_rflag,
  input         io_bypass_2_bits_fflags_bits_uop_wflag,
  input  [3:0]  io_bypass_2_bits_fflags_bits_uop_prflag,
  input  [3:0]  io_bypass_2_bits_fflags_bits_uop_pwflag,
  input         io_bypass_2_bits_fflags_bits_uop_pflag_busy,
  input  [3:0]  io_bypass_2_bits_fflags_bits_uop_stale_pflag,
  input  [3:0]  io_bypass_2_bits_fflags_bits_uop_op1_sel,
  input  [3:0]  io_bypass_2_bits_fflags_bits_uop_op2_sel,
  input  [5:0]  io_bypass_2_bits_fflags_bits_uop_split_num,
  input  [5:0]  io_bypass_2_bits_fflags_bits_uop_self_index,
  input  [5:0]  io_bypass_2_bits_fflags_bits_uop_rob_inst_idx,
  input  [5:0]  io_bypass_2_bits_fflags_bits_uop_address_num,
  input  [6:0]  io_bypass_2_bits_fflags_bits_uop_uopc,
  input  [31:0] io_bypass_2_bits_fflags_bits_uop_inst,
  input  [31:0] io_bypass_2_bits_fflags_bits_uop_debug_inst,
  input         io_bypass_2_bits_fflags_bits_uop_is_rvc,
  input  [39:0] io_bypass_2_bits_fflags_bits_uop_debug_pc,
  input  [2:0]  io_bypass_2_bits_fflags_bits_uop_iq_type,
  input  [9:0]  io_bypass_2_bits_fflags_bits_uop_fu_code,
  input  [3:0]  io_bypass_2_bits_fflags_bits_uop_ctrl_br_type,
  input  [1:0]  io_bypass_2_bits_fflags_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_bypass_2_bits_fflags_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_bypass_2_bits_fflags_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_bypass_2_bits_fflags_bits_uop_ctrl_op_fcn,
  input         io_bypass_2_bits_fflags_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_bypass_2_bits_fflags_bits_uop_ctrl_csr_cmd,
  input         io_bypass_2_bits_fflags_bits_uop_ctrl_is_load,
  input         io_bypass_2_bits_fflags_bits_uop_ctrl_is_sta,
  input         io_bypass_2_bits_fflags_bits_uop_ctrl_is_std,
  input  [1:0]  io_bypass_2_bits_fflags_bits_uop_ctrl_op3_sel,
  input  [1:0]  io_bypass_2_bits_fflags_bits_uop_iw_state,
  input         io_bypass_2_bits_fflags_bits_uop_iw_p1_poisoned,
  input         io_bypass_2_bits_fflags_bits_uop_iw_p2_poisoned,
  input         io_bypass_2_bits_fflags_bits_uop_is_br,
  input         io_bypass_2_bits_fflags_bits_uop_is_jalr,
  input         io_bypass_2_bits_fflags_bits_uop_is_jal,
  input         io_bypass_2_bits_fflags_bits_uop_is_sfb,
  input  [11:0] io_bypass_2_bits_fflags_bits_uop_br_mask,
  input  [3:0]  io_bypass_2_bits_fflags_bits_uop_br_tag,
  input  [4:0]  io_bypass_2_bits_fflags_bits_uop_ftq_idx,
  input         io_bypass_2_bits_fflags_bits_uop_edge_inst,
  input  [5:0]  io_bypass_2_bits_fflags_bits_uop_pc_lob,
  input         io_bypass_2_bits_fflags_bits_uop_taken,
  input  [19:0] io_bypass_2_bits_fflags_bits_uop_imm_packed,
  input  [11:0] io_bypass_2_bits_fflags_bits_uop_csr_addr,
  input  [5:0]  io_bypass_2_bits_fflags_bits_uop_rob_idx,
  input  [4:0]  io_bypass_2_bits_fflags_bits_uop_ldq_idx,
  input  [4:0]  io_bypass_2_bits_fflags_bits_uop_stq_idx,
  input  [1:0]  io_bypass_2_bits_fflags_bits_uop_rxq_idx,
  input  [6:0]  io_bypass_2_bits_fflags_bits_uop_pdst,
  input  [6:0]  io_bypass_2_bits_fflags_bits_uop_prs1,
  input  [6:0]  io_bypass_2_bits_fflags_bits_uop_prs2,
  input  [6:0]  io_bypass_2_bits_fflags_bits_uop_prs3,
  input  [4:0]  io_bypass_2_bits_fflags_bits_uop_ppred,
  input         io_bypass_2_bits_fflags_bits_uop_prs1_busy,
  input         io_bypass_2_bits_fflags_bits_uop_prs2_busy,
  input         io_bypass_2_bits_fflags_bits_uop_prs3_busy,
  input         io_bypass_2_bits_fflags_bits_uop_ppred_busy,
  input  [6:0]  io_bypass_2_bits_fflags_bits_uop_stale_pdst,
  input         io_bypass_2_bits_fflags_bits_uop_exception,
  input  [63:0] io_bypass_2_bits_fflags_bits_uop_exc_cause,
  input         io_bypass_2_bits_fflags_bits_uop_bypassable,
  input  [4:0]  io_bypass_2_bits_fflags_bits_uop_mem_cmd,
  input  [1:0]  io_bypass_2_bits_fflags_bits_uop_mem_size,
  input         io_bypass_2_bits_fflags_bits_uop_mem_signed,
  input         io_bypass_2_bits_fflags_bits_uop_is_fence,
  input         io_bypass_2_bits_fflags_bits_uop_is_fencei,
  input         io_bypass_2_bits_fflags_bits_uop_is_amo,
  input         io_bypass_2_bits_fflags_bits_uop_uses_ldq,
  input         io_bypass_2_bits_fflags_bits_uop_uses_stq,
  input         io_bypass_2_bits_fflags_bits_uop_is_sys_pc2epc,
  input         io_bypass_2_bits_fflags_bits_uop_is_unique,
  input         io_bypass_2_bits_fflags_bits_uop_flush_on_commit,
  input         io_bypass_2_bits_fflags_bits_uop_ldst_is_rs1,
  input  [5:0]  io_bypass_2_bits_fflags_bits_uop_ldst,
  input  [5:0]  io_bypass_2_bits_fflags_bits_uop_lrs1,
  input  [5:0]  io_bypass_2_bits_fflags_bits_uop_lrs2,
  input  [5:0]  io_bypass_2_bits_fflags_bits_uop_lrs3,
  input         io_bypass_2_bits_fflags_bits_uop_ldst_val,
  input  [1:0]  io_bypass_2_bits_fflags_bits_uop_dst_rtype,
  input  [1:0]  io_bypass_2_bits_fflags_bits_uop_lrs1_rtype,
  input  [1:0]  io_bypass_2_bits_fflags_bits_uop_lrs2_rtype,
  input         io_bypass_2_bits_fflags_bits_uop_frs3_en,
  input         io_bypass_2_bits_fflags_bits_uop_fp_val,
  input         io_bypass_2_bits_fflags_bits_uop_fp_single,
  input         io_bypass_2_bits_fflags_bits_uop_xcpt_pf_if,
  input         io_bypass_2_bits_fflags_bits_uop_xcpt_ae_if,
  input         io_bypass_2_bits_fflags_bits_uop_xcpt_ma_if,
  input         io_bypass_2_bits_fflags_bits_uop_bp_debug_if,
  input         io_bypass_2_bits_fflags_bits_uop_bp_xcpt_if,
  input  [1:0]  io_bypass_2_bits_fflags_bits_uop_debug_fsrc,
  input  [1:0]  io_bypass_2_bits_fflags_bits_uop_debug_tsrc,
  input  [4:0]  io_bypass_2_bits_fflags_bits_flags,
  input  [3:0]  io_bypass_2_bits_flagdata,
  input         io_bypass_2_bits_fflagdata_valid,
  input         io_bypass_2_bits_fflagdata_bits_uop_switch,
  input         io_bypass_2_bits_fflagdata_bits_uop_switch_off,
  input         io_bypass_2_bits_fflagdata_bits_uop_is_unicore,
  input  [2:0]  io_bypass_2_bits_fflagdata_bits_uop_shift,
  input  [1:0]  io_bypass_2_bits_fflagdata_bits_uop_lrs3_rtype,
  input         io_bypass_2_bits_fflagdata_bits_uop_rflag,
  input         io_bypass_2_bits_fflagdata_bits_uop_wflag,
  input  [3:0]  io_bypass_2_bits_fflagdata_bits_uop_prflag,
  input  [3:0]  io_bypass_2_bits_fflagdata_bits_uop_pwflag,
  input         io_bypass_2_bits_fflagdata_bits_uop_pflag_busy,
  input  [3:0]  io_bypass_2_bits_fflagdata_bits_uop_stale_pflag,
  input  [3:0]  io_bypass_2_bits_fflagdata_bits_uop_op1_sel,
  input  [3:0]  io_bypass_2_bits_fflagdata_bits_uop_op2_sel,
  input  [5:0]  io_bypass_2_bits_fflagdata_bits_uop_split_num,
  input  [5:0]  io_bypass_2_bits_fflagdata_bits_uop_self_index,
  input  [5:0]  io_bypass_2_bits_fflagdata_bits_uop_rob_inst_idx,
  input  [5:0]  io_bypass_2_bits_fflagdata_bits_uop_address_num,
  input  [6:0]  io_bypass_2_bits_fflagdata_bits_uop_uopc,
  input  [31:0] io_bypass_2_bits_fflagdata_bits_uop_inst,
  input  [31:0] io_bypass_2_bits_fflagdata_bits_uop_debug_inst,
  input         io_bypass_2_bits_fflagdata_bits_uop_is_rvc,
  input  [39:0] io_bypass_2_bits_fflagdata_bits_uop_debug_pc,
  input  [2:0]  io_bypass_2_bits_fflagdata_bits_uop_iq_type,
  input  [9:0]  io_bypass_2_bits_fflagdata_bits_uop_fu_code,
  input  [3:0]  io_bypass_2_bits_fflagdata_bits_uop_ctrl_br_type,
  input  [1:0]  io_bypass_2_bits_fflagdata_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_bypass_2_bits_fflagdata_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_bypass_2_bits_fflagdata_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_bypass_2_bits_fflagdata_bits_uop_ctrl_op_fcn,
  input         io_bypass_2_bits_fflagdata_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_bypass_2_bits_fflagdata_bits_uop_ctrl_csr_cmd,
  input         io_bypass_2_bits_fflagdata_bits_uop_ctrl_is_load,
  input         io_bypass_2_bits_fflagdata_bits_uop_ctrl_is_sta,
  input         io_bypass_2_bits_fflagdata_bits_uop_ctrl_is_std,
  input  [1:0]  io_bypass_2_bits_fflagdata_bits_uop_ctrl_op3_sel,
  input  [1:0]  io_bypass_2_bits_fflagdata_bits_uop_iw_state,
  input         io_bypass_2_bits_fflagdata_bits_uop_iw_p1_poisoned,
  input         io_bypass_2_bits_fflagdata_bits_uop_iw_p2_poisoned,
  input         io_bypass_2_bits_fflagdata_bits_uop_is_br,
  input         io_bypass_2_bits_fflagdata_bits_uop_is_jalr,
  input         io_bypass_2_bits_fflagdata_bits_uop_is_jal,
  input         io_bypass_2_bits_fflagdata_bits_uop_is_sfb,
  input  [11:0] io_bypass_2_bits_fflagdata_bits_uop_br_mask,
  input  [3:0]  io_bypass_2_bits_fflagdata_bits_uop_br_tag,
  input  [4:0]  io_bypass_2_bits_fflagdata_bits_uop_ftq_idx,
  input         io_bypass_2_bits_fflagdata_bits_uop_edge_inst,
  input  [5:0]  io_bypass_2_bits_fflagdata_bits_uop_pc_lob,
  input         io_bypass_2_bits_fflagdata_bits_uop_taken,
  input  [19:0] io_bypass_2_bits_fflagdata_bits_uop_imm_packed,
  input  [11:0] io_bypass_2_bits_fflagdata_bits_uop_csr_addr,
  input  [5:0]  io_bypass_2_bits_fflagdata_bits_uop_rob_idx,
  input  [4:0]  io_bypass_2_bits_fflagdata_bits_uop_ldq_idx,
  input  [4:0]  io_bypass_2_bits_fflagdata_bits_uop_stq_idx,
  input  [1:0]  io_bypass_2_bits_fflagdata_bits_uop_rxq_idx,
  input  [6:0]  io_bypass_2_bits_fflagdata_bits_uop_pdst,
  input  [6:0]  io_bypass_2_bits_fflagdata_bits_uop_prs1,
  input  [6:0]  io_bypass_2_bits_fflagdata_bits_uop_prs2,
  input  [6:0]  io_bypass_2_bits_fflagdata_bits_uop_prs3,
  input  [4:0]  io_bypass_2_bits_fflagdata_bits_uop_ppred,
  input         io_bypass_2_bits_fflagdata_bits_uop_prs1_busy,
  input         io_bypass_2_bits_fflagdata_bits_uop_prs2_busy,
  input         io_bypass_2_bits_fflagdata_bits_uop_prs3_busy,
  input         io_bypass_2_bits_fflagdata_bits_uop_ppred_busy,
  input  [6:0]  io_bypass_2_bits_fflagdata_bits_uop_stale_pdst,
  input         io_bypass_2_bits_fflagdata_bits_uop_exception,
  input  [63:0] io_bypass_2_bits_fflagdata_bits_uop_exc_cause,
  input         io_bypass_2_bits_fflagdata_bits_uop_bypassable,
  input  [4:0]  io_bypass_2_bits_fflagdata_bits_uop_mem_cmd,
  input  [1:0]  io_bypass_2_bits_fflagdata_bits_uop_mem_size,
  input         io_bypass_2_bits_fflagdata_bits_uop_mem_signed,
  input         io_bypass_2_bits_fflagdata_bits_uop_is_fence,
  input         io_bypass_2_bits_fflagdata_bits_uop_is_fencei,
  input         io_bypass_2_bits_fflagdata_bits_uop_is_amo,
  input         io_bypass_2_bits_fflagdata_bits_uop_uses_ldq,
  input         io_bypass_2_bits_fflagdata_bits_uop_uses_stq,
  input         io_bypass_2_bits_fflagdata_bits_uop_is_sys_pc2epc,
  input         io_bypass_2_bits_fflagdata_bits_uop_is_unique,
  input         io_bypass_2_bits_fflagdata_bits_uop_flush_on_commit,
  input         io_bypass_2_bits_fflagdata_bits_uop_ldst_is_rs1,
  input  [5:0]  io_bypass_2_bits_fflagdata_bits_uop_ldst,
  input  [5:0]  io_bypass_2_bits_fflagdata_bits_uop_lrs1,
  input  [5:0]  io_bypass_2_bits_fflagdata_bits_uop_lrs2,
  input  [5:0]  io_bypass_2_bits_fflagdata_bits_uop_lrs3,
  input         io_bypass_2_bits_fflagdata_bits_uop_ldst_val,
  input  [1:0]  io_bypass_2_bits_fflagdata_bits_uop_dst_rtype,
  input  [1:0]  io_bypass_2_bits_fflagdata_bits_uop_lrs1_rtype,
  input  [1:0]  io_bypass_2_bits_fflagdata_bits_uop_lrs2_rtype,
  input         io_bypass_2_bits_fflagdata_bits_uop_frs3_en,
  input         io_bypass_2_bits_fflagdata_bits_uop_fp_val,
  input         io_bypass_2_bits_fflagdata_bits_uop_fp_single,
  input         io_bypass_2_bits_fflagdata_bits_uop_xcpt_pf_if,
  input         io_bypass_2_bits_fflagdata_bits_uop_xcpt_ae_if,
  input         io_bypass_2_bits_fflagdata_bits_uop_xcpt_ma_if,
  input         io_bypass_2_bits_fflagdata_bits_uop_bp_debug_if,
  input         io_bypass_2_bits_fflagdata_bits_uop_bp_xcpt_if,
  input  [1:0]  io_bypass_2_bits_fflagdata_bits_uop_debug_fsrc,
  input  [1:0]  io_bypass_2_bits_fflagdata_bits_uop_debug_tsrc,
  input  [31:0] io_bypass_2_bits_fflagdata_bits_fflag,
  input         io_bypass_3_valid,
  input         io_bypass_3_bits_uop_switch,
  input         io_bypass_3_bits_uop_switch_off,
  input         io_bypass_3_bits_uop_is_unicore,
  input  [2:0]  io_bypass_3_bits_uop_shift,
  input  [1:0]  io_bypass_3_bits_uop_lrs3_rtype,
  input         io_bypass_3_bits_uop_rflag,
  input         io_bypass_3_bits_uop_wflag,
  input  [3:0]  io_bypass_3_bits_uop_prflag,
  input  [3:0]  io_bypass_3_bits_uop_pwflag,
  input         io_bypass_3_bits_uop_pflag_busy,
  input  [3:0]  io_bypass_3_bits_uop_stale_pflag,
  input  [3:0]  io_bypass_3_bits_uop_op1_sel,
  input  [3:0]  io_bypass_3_bits_uop_op2_sel,
  input  [5:0]  io_bypass_3_bits_uop_split_num,
  input  [5:0]  io_bypass_3_bits_uop_self_index,
  input  [5:0]  io_bypass_3_bits_uop_rob_inst_idx,
  input  [5:0]  io_bypass_3_bits_uop_address_num,
  input  [6:0]  io_bypass_3_bits_uop_uopc,
  input  [31:0] io_bypass_3_bits_uop_inst,
  input  [31:0] io_bypass_3_bits_uop_debug_inst,
  input         io_bypass_3_bits_uop_is_rvc,
  input  [39:0] io_bypass_3_bits_uop_debug_pc,
  input  [2:0]  io_bypass_3_bits_uop_iq_type,
  input  [9:0]  io_bypass_3_bits_uop_fu_code,
  input  [3:0]  io_bypass_3_bits_uop_ctrl_br_type,
  input  [1:0]  io_bypass_3_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_bypass_3_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_bypass_3_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_bypass_3_bits_uop_ctrl_op_fcn,
  input         io_bypass_3_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_bypass_3_bits_uop_ctrl_csr_cmd,
  input         io_bypass_3_bits_uop_ctrl_is_load,
  input         io_bypass_3_bits_uop_ctrl_is_sta,
  input         io_bypass_3_bits_uop_ctrl_is_std,
  input  [1:0]  io_bypass_3_bits_uop_ctrl_op3_sel,
  input  [1:0]  io_bypass_3_bits_uop_iw_state,
  input         io_bypass_3_bits_uop_iw_p1_poisoned,
  input         io_bypass_3_bits_uop_iw_p2_poisoned,
  input         io_bypass_3_bits_uop_is_br,
  input         io_bypass_3_bits_uop_is_jalr,
  input         io_bypass_3_bits_uop_is_jal,
  input         io_bypass_3_bits_uop_is_sfb,
  input  [11:0] io_bypass_3_bits_uop_br_mask,
  input  [3:0]  io_bypass_3_bits_uop_br_tag,
  input  [4:0]  io_bypass_3_bits_uop_ftq_idx,
  input         io_bypass_3_bits_uop_edge_inst,
  input  [5:0]  io_bypass_3_bits_uop_pc_lob,
  input         io_bypass_3_bits_uop_taken,
  input  [19:0] io_bypass_3_bits_uop_imm_packed,
  input  [11:0] io_bypass_3_bits_uop_csr_addr,
  input  [5:0]  io_bypass_3_bits_uop_rob_idx,
  input  [4:0]  io_bypass_3_bits_uop_ldq_idx,
  input  [4:0]  io_bypass_3_bits_uop_stq_idx,
  input  [1:0]  io_bypass_3_bits_uop_rxq_idx,
  input  [6:0]  io_bypass_3_bits_uop_pdst,
  input  [6:0]  io_bypass_3_bits_uop_prs1,
  input  [6:0]  io_bypass_3_bits_uop_prs2,
  input  [6:0]  io_bypass_3_bits_uop_prs3,
  input  [4:0]  io_bypass_3_bits_uop_ppred,
  input         io_bypass_3_bits_uop_prs1_busy,
  input         io_bypass_3_bits_uop_prs2_busy,
  input         io_bypass_3_bits_uop_prs3_busy,
  input         io_bypass_3_bits_uop_ppred_busy,
  input  [6:0]  io_bypass_3_bits_uop_stale_pdst,
  input         io_bypass_3_bits_uop_exception,
  input  [63:0] io_bypass_3_bits_uop_exc_cause,
  input         io_bypass_3_bits_uop_bypassable,
  input  [4:0]  io_bypass_3_bits_uop_mem_cmd,
  input  [1:0]  io_bypass_3_bits_uop_mem_size,
  input         io_bypass_3_bits_uop_mem_signed,
  input         io_bypass_3_bits_uop_is_fence,
  input         io_bypass_3_bits_uop_is_fencei,
  input         io_bypass_3_bits_uop_is_amo,
  input         io_bypass_3_bits_uop_uses_ldq,
  input         io_bypass_3_bits_uop_uses_stq,
  input         io_bypass_3_bits_uop_is_sys_pc2epc,
  input         io_bypass_3_bits_uop_is_unique,
  input         io_bypass_3_bits_uop_flush_on_commit,
  input         io_bypass_3_bits_uop_ldst_is_rs1,
  input  [5:0]  io_bypass_3_bits_uop_ldst,
  input  [5:0]  io_bypass_3_bits_uop_lrs1,
  input  [5:0]  io_bypass_3_bits_uop_lrs2,
  input  [5:0]  io_bypass_3_bits_uop_lrs3,
  input         io_bypass_3_bits_uop_ldst_val,
  input  [1:0]  io_bypass_3_bits_uop_dst_rtype,
  input  [1:0]  io_bypass_3_bits_uop_lrs1_rtype,
  input  [1:0]  io_bypass_3_bits_uop_lrs2_rtype,
  input         io_bypass_3_bits_uop_frs3_en,
  input         io_bypass_3_bits_uop_fp_val,
  input         io_bypass_3_bits_uop_fp_single,
  input         io_bypass_3_bits_uop_xcpt_pf_if,
  input         io_bypass_3_bits_uop_xcpt_ae_if,
  input         io_bypass_3_bits_uop_xcpt_ma_if,
  input         io_bypass_3_bits_uop_bp_debug_if,
  input         io_bypass_3_bits_uop_bp_xcpt_if,
  input  [1:0]  io_bypass_3_bits_uop_debug_fsrc,
  input  [1:0]  io_bypass_3_bits_uop_debug_tsrc,
  input  [63:0] io_bypass_3_bits_data,
  input         io_bypass_3_bits_predicated,
  input         io_bypass_3_bits_fflags_valid,
  input         io_bypass_3_bits_fflags_bits_uop_switch,
  input         io_bypass_3_bits_fflags_bits_uop_switch_off,
  input         io_bypass_3_bits_fflags_bits_uop_is_unicore,
  input  [2:0]  io_bypass_3_bits_fflags_bits_uop_shift,
  input  [1:0]  io_bypass_3_bits_fflags_bits_uop_lrs3_rtype,
  input         io_bypass_3_bits_fflags_bits_uop_rflag,
  input         io_bypass_3_bits_fflags_bits_uop_wflag,
  input  [3:0]  io_bypass_3_bits_fflags_bits_uop_prflag,
  input  [3:0]  io_bypass_3_bits_fflags_bits_uop_pwflag,
  input         io_bypass_3_bits_fflags_bits_uop_pflag_busy,
  input  [3:0]  io_bypass_3_bits_fflags_bits_uop_stale_pflag,
  input  [3:0]  io_bypass_3_bits_fflags_bits_uop_op1_sel,
  input  [3:0]  io_bypass_3_bits_fflags_bits_uop_op2_sel,
  input  [5:0]  io_bypass_3_bits_fflags_bits_uop_split_num,
  input  [5:0]  io_bypass_3_bits_fflags_bits_uop_self_index,
  input  [5:0]  io_bypass_3_bits_fflags_bits_uop_rob_inst_idx,
  input  [5:0]  io_bypass_3_bits_fflags_bits_uop_address_num,
  input  [6:0]  io_bypass_3_bits_fflags_bits_uop_uopc,
  input  [31:0] io_bypass_3_bits_fflags_bits_uop_inst,
  input  [31:0] io_bypass_3_bits_fflags_bits_uop_debug_inst,
  input         io_bypass_3_bits_fflags_bits_uop_is_rvc,
  input  [39:0] io_bypass_3_bits_fflags_bits_uop_debug_pc,
  input  [2:0]  io_bypass_3_bits_fflags_bits_uop_iq_type,
  input  [9:0]  io_bypass_3_bits_fflags_bits_uop_fu_code,
  input  [3:0]  io_bypass_3_bits_fflags_bits_uop_ctrl_br_type,
  input  [1:0]  io_bypass_3_bits_fflags_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_bypass_3_bits_fflags_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_bypass_3_bits_fflags_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_bypass_3_bits_fflags_bits_uop_ctrl_op_fcn,
  input         io_bypass_3_bits_fflags_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_bypass_3_bits_fflags_bits_uop_ctrl_csr_cmd,
  input         io_bypass_3_bits_fflags_bits_uop_ctrl_is_load,
  input         io_bypass_3_bits_fflags_bits_uop_ctrl_is_sta,
  input         io_bypass_3_bits_fflags_bits_uop_ctrl_is_std,
  input  [1:0]  io_bypass_3_bits_fflags_bits_uop_ctrl_op3_sel,
  input  [1:0]  io_bypass_3_bits_fflags_bits_uop_iw_state,
  input         io_bypass_3_bits_fflags_bits_uop_iw_p1_poisoned,
  input         io_bypass_3_bits_fflags_bits_uop_iw_p2_poisoned,
  input         io_bypass_3_bits_fflags_bits_uop_is_br,
  input         io_bypass_3_bits_fflags_bits_uop_is_jalr,
  input         io_bypass_3_bits_fflags_bits_uop_is_jal,
  input         io_bypass_3_bits_fflags_bits_uop_is_sfb,
  input  [11:0] io_bypass_3_bits_fflags_bits_uop_br_mask,
  input  [3:0]  io_bypass_3_bits_fflags_bits_uop_br_tag,
  input  [4:0]  io_bypass_3_bits_fflags_bits_uop_ftq_idx,
  input         io_bypass_3_bits_fflags_bits_uop_edge_inst,
  input  [5:0]  io_bypass_3_bits_fflags_bits_uop_pc_lob,
  input         io_bypass_3_bits_fflags_bits_uop_taken,
  input  [19:0] io_bypass_3_bits_fflags_bits_uop_imm_packed,
  input  [11:0] io_bypass_3_bits_fflags_bits_uop_csr_addr,
  input  [5:0]  io_bypass_3_bits_fflags_bits_uop_rob_idx,
  input  [4:0]  io_bypass_3_bits_fflags_bits_uop_ldq_idx,
  input  [4:0]  io_bypass_3_bits_fflags_bits_uop_stq_idx,
  input  [1:0]  io_bypass_3_bits_fflags_bits_uop_rxq_idx,
  input  [6:0]  io_bypass_3_bits_fflags_bits_uop_pdst,
  input  [6:0]  io_bypass_3_bits_fflags_bits_uop_prs1,
  input  [6:0]  io_bypass_3_bits_fflags_bits_uop_prs2,
  input  [6:0]  io_bypass_3_bits_fflags_bits_uop_prs3,
  input  [4:0]  io_bypass_3_bits_fflags_bits_uop_ppred,
  input         io_bypass_3_bits_fflags_bits_uop_prs1_busy,
  input         io_bypass_3_bits_fflags_bits_uop_prs2_busy,
  input         io_bypass_3_bits_fflags_bits_uop_prs3_busy,
  input         io_bypass_3_bits_fflags_bits_uop_ppred_busy,
  input  [6:0]  io_bypass_3_bits_fflags_bits_uop_stale_pdst,
  input         io_bypass_3_bits_fflags_bits_uop_exception,
  input  [63:0] io_bypass_3_bits_fflags_bits_uop_exc_cause,
  input         io_bypass_3_bits_fflags_bits_uop_bypassable,
  input  [4:0]  io_bypass_3_bits_fflags_bits_uop_mem_cmd,
  input  [1:0]  io_bypass_3_bits_fflags_bits_uop_mem_size,
  input         io_bypass_3_bits_fflags_bits_uop_mem_signed,
  input         io_bypass_3_bits_fflags_bits_uop_is_fence,
  input         io_bypass_3_bits_fflags_bits_uop_is_fencei,
  input         io_bypass_3_bits_fflags_bits_uop_is_amo,
  input         io_bypass_3_bits_fflags_bits_uop_uses_ldq,
  input         io_bypass_3_bits_fflags_bits_uop_uses_stq,
  input         io_bypass_3_bits_fflags_bits_uop_is_sys_pc2epc,
  input         io_bypass_3_bits_fflags_bits_uop_is_unique,
  input         io_bypass_3_bits_fflags_bits_uop_flush_on_commit,
  input         io_bypass_3_bits_fflags_bits_uop_ldst_is_rs1,
  input  [5:0]  io_bypass_3_bits_fflags_bits_uop_ldst,
  input  [5:0]  io_bypass_3_bits_fflags_bits_uop_lrs1,
  input  [5:0]  io_bypass_3_bits_fflags_bits_uop_lrs2,
  input  [5:0]  io_bypass_3_bits_fflags_bits_uop_lrs3,
  input         io_bypass_3_bits_fflags_bits_uop_ldst_val,
  input  [1:0]  io_bypass_3_bits_fflags_bits_uop_dst_rtype,
  input  [1:0]  io_bypass_3_bits_fflags_bits_uop_lrs1_rtype,
  input  [1:0]  io_bypass_3_bits_fflags_bits_uop_lrs2_rtype,
  input         io_bypass_3_bits_fflags_bits_uop_frs3_en,
  input         io_bypass_3_bits_fflags_bits_uop_fp_val,
  input         io_bypass_3_bits_fflags_bits_uop_fp_single,
  input         io_bypass_3_bits_fflags_bits_uop_xcpt_pf_if,
  input         io_bypass_3_bits_fflags_bits_uop_xcpt_ae_if,
  input         io_bypass_3_bits_fflags_bits_uop_xcpt_ma_if,
  input         io_bypass_3_bits_fflags_bits_uop_bp_debug_if,
  input         io_bypass_3_bits_fflags_bits_uop_bp_xcpt_if,
  input  [1:0]  io_bypass_3_bits_fflags_bits_uop_debug_fsrc,
  input  [1:0]  io_bypass_3_bits_fflags_bits_uop_debug_tsrc,
  input  [4:0]  io_bypass_3_bits_fflags_bits_flags,
  input  [3:0]  io_bypass_3_bits_flagdata,
  input         io_bypass_3_bits_fflagdata_valid,
  input         io_bypass_3_bits_fflagdata_bits_uop_switch,
  input         io_bypass_3_bits_fflagdata_bits_uop_switch_off,
  input         io_bypass_3_bits_fflagdata_bits_uop_is_unicore,
  input  [2:0]  io_bypass_3_bits_fflagdata_bits_uop_shift,
  input  [1:0]  io_bypass_3_bits_fflagdata_bits_uop_lrs3_rtype,
  input         io_bypass_3_bits_fflagdata_bits_uop_rflag,
  input         io_bypass_3_bits_fflagdata_bits_uop_wflag,
  input  [3:0]  io_bypass_3_bits_fflagdata_bits_uop_prflag,
  input  [3:0]  io_bypass_3_bits_fflagdata_bits_uop_pwflag,
  input         io_bypass_3_bits_fflagdata_bits_uop_pflag_busy,
  input  [3:0]  io_bypass_3_bits_fflagdata_bits_uop_stale_pflag,
  input  [3:0]  io_bypass_3_bits_fflagdata_bits_uop_op1_sel,
  input  [3:0]  io_bypass_3_bits_fflagdata_bits_uop_op2_sel,
  input  [5:0]  io_bypass_3_bits_fflagdata_bits_uop_split_num,
  input  [5:0]  io_bypass_3_bits_fflagdata_bits_uop_self_index,
  input  [5:0]  io_bypass_3_bits_fflagdata_bits_uop_rob_inst_idx,
  input  [5:0]  io_bypass_3_bits_fflagdata_bits_uop_address_num,
  input  [6:0]  io_bypass_3_bits_fflagdata_bits_uop_uopc,
  input  [31:0] io_bypass_3_bits_fflagdata_bits_uop_inst,
  input  [31:0] io_bypass_3_bits_fflagdata_bits_uop_debug_inst,
  input         io_bypass_3_bits_fflagdata_bits_uop_is_rvc,
  input  [39:0] io_bypass_3_bits_fflagdata_bits_uop_debug_pc,
  input  [2:0]  io_bypass_3_bits_fflagdata_bits_uop_iq_type,
  input  [9:0]  io_bypass_3_bits_fflagdata_bits_uop_fu_code,
  input  [3:0]  io_bypass_3_bits_fflagdata_bits_uop_ctrl_br_type,
  input  [1:0]  io_bypass_3_bits_fflagdata_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_bypass_3_bits_fflagdata_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_bypass_3_bits_fflagdata_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_bypass_3_bits_fflagdata_bits_uop_ctrl_op_fcn,
  input         io_bypass_3_bits_fflagdata_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_bypass_3_bits_fflagdata_bits_uop_ctrl_csr_cmd,
  input         io_bypass_3_bits_fflagdata_bits_uop_ctrl_is_load,
  input         io_bypass_3_bits_fflagdata_bits_uop_ctrl_is_sta,
  input         io_bypass_3_bits_fflagdata_bits_uop_ctrl_is_std,
  input  [1:0]  io_bypass_3_bits_fflagdata_bits_uop_ctrl_op3_sel,
  input  [1:0]  io_bypass_3_bits_fflagdata_bits_uop_iw_state,
  input         io_bypass_3_bits_fflagdata_bits_uop_iw_p1_poisoned,
  input         io_bypass_3_bits_fflagdata_bits_uop_iw_p2_poisoned,
  input         io_bypass_3_bits_fflagdata_bits_uop_is_br,
  input         io_bypass_3_bits_fflagdata_bits_uop_is_jalr,
  input         io_bypass_3_bits_fflagdata_bits_uop_is_jal,
  input         io_bypass_3_bits_fflagdata_bits_uop_is_sfb,
  input  [11:0] io_bypass_3_bits_fflagdata_bits_uop_br_mask,
  input  [3:0]  io_bypass_3_bits_fflagdata_bits_uop_br_tag,
  input  [4:0]  io_bypass_3_bits_fflagdata_bits_uop_ftq_idx,
  input         io_bypass_3_bits_fflagdata_bits_uop_edge_inst,
  input  [5:0]  io_bypass_3_bits_fflagdata_bits_uop_pc_lob,
  input         io_bypass_3_bits_fflagdata_bits_uop_taken,
  input  [19:0] io_bypass_3_bits_fflagdata_bits_uop_imm_packed,
  input  [11:0] io_bypass_3_bits_fflagdata_bits_uop_csr_addr,
  input  [5:0]  io_bypass_3_bits_fflagdata_bits_uop_rob_idx,
  input  [4:0]  io_bypass_3_bits_fflagdata_bits_uop_ldq_idx,
  input  [4:0]  io_bypass_3_bits_fflagdata_bits_uop_stq_idx,
  input  [1:0]  io_bypass_3_bits_fflagdata_bits_uop_rxq_idx,
  input  [6:0]  io_bypass_3_bits_fflagdata_bits_uop_pdst,
  input  [6:0]  io_bypass_3_bits_fflagdata_bits_uop_prs1,
  input  [6:0]  io_bypass_3_bits_fflagdata_bits_uop_prs2,
  input  [6:0]  io_bypass_3_bits_fflagdata_bits_uop_prs3,
  input  [4:0]  io_bypass_3_bits_fflagdata_bits_uop_ppred,
  input         io_bypass_3_bits_fflagdata_bits_uop_prs1_busy,
  input         io_bypass_3_bits_fflagdata_bits_uop_prs2_busy,
  input         io_bypass_3_bits_fflagdata_bits_uop_prs3_busy,
  input         io_bypass_3_bits_fflagdata_bits_uop_ppred_busy,
  input  [6:0]  io_bypass_3_bits_fflagdata_bits_uop_stale_pdst,
  input         io_bypass_3_bits_fflagdata_bits_uop_exception,
  input  [63:0] io_bypass_3_bits_fflagdata_bits_uop_exc_cause,
  input         io_bypass_3_bits_fflagdata_bits_uop_bypassable,
  input  [4:0]  io_bypass_3_bits_fflagdata_bits_uop_mem_cmd,
  input  [1:0]  io_bypass_3_bits_fflagdata_bits_uop_mem_size,
  input         io_bypass_3_bits_fflagdata_bits_uop_mem_signed,
  input         io_bypass_3_bits_fflagdata_bits_uop_is_fence,
  input         io_bypass_3_bits_fflagdata_bits_uop_is_fencei,
  input         io_bypass_3_bits_fflagdata_bits_uop_is_amo,
  input         io_bypass_3_bits_fflagdata_bits_uop_uses_ldq,
  input         io_bypass_3_bits_fflagdata_bits_uop_uses_stq,
  input         io_bypass_3_bits_fflagdata_bits_uop_is_sys_pc2epc,
  input         io_bypass_3_bits_fflagdata_bits_uop_is_unique,
  input         io_bypass_3_bits_fflagdata_bits_uop_flush_on_commit,
  input         io_bypass_3_bits_fflagdata_bits_uop_ldst_is_rs1,
  input  [5:0]  io_bypass_3_bits_fflagdata_bits_uop_ldst,
  input  [5:0]  io_bypass_3_bits_fflagdata_bits_uop_lrs1,
  input  [5:0]  io_bypass_3_bits_fflagdata_bits_uop_lrs2,
  input  [5:0]  io_bypass_3_bits_fflagdata_bits_uop_lrs3,
  input         io_bypass_3_bits_fflagdata_bits_uop_ldst_val,
  input  [1:0]  io_bypass_3_bits_fflagdata_bits_uop_dst_rtype,
  input  [1:0]  io_bypass_3_bits_fflagdata_bits_uop_lrs1_rtype,
  input  [1:0]  io_bypass_3_bits_fflagdata_bits_uop_lrs2_rtype,
  input         io_bypass_3_bits_fflagdata_bits_uop_frs3_en,
  input         io_bypass_3_bits_fflagdata_bits_uop_fp_val,
  input         io_bypass_3_bits_fflagdata_bits_uop_fp_single,
  input         io_bypass_3_bits_fflagdata_bits_uop_xcpt_pf_if,
  input         io_bypass_3_bits_fflagdata_bits_uop_xcpt_ae_if,
  input         io_bypass_3_bits_fflagdata_bits_uop_xcpt_ma_if,
  input         io_bypass_3_bits_fflagdata_bits_uop_bp_debug_if,
  input         io_bypass_3_bits_fflagdata_bits_uop_bp_xcpt_if,
  input  [1:0]  io_bypass_3_bits_fflagdata_bits_uop_debug_fsrc,
  input  [1:0]  io_bypass_3_bits_fflagdata_bits_uop_debug_tsrc,
  input  [31:0] io_bypass_3_bits_fflagdata_bits_fflag,
  input         io_pred_bypass_0_valid,
  input         io_pred_bypass_0_bits_uop_switch,
  input         io_pred_bypass_0_bits_uop_switch_off,
  input         io_pred_bypass_0_bits_uop_is_unicore,
  input  [2:0]  io_pred_bypass_0_bits_uop_shift,
  input  [1:0]  io_pred_bypass_0_bits_uop_lrs3_rtype,
  input         io_pred_bypass_0_bits_uop_rflag,
  input         io_pred_bypass_0_bits_uop_wflag,
  input  [3:0]  io_pred_bypass_0_bits_uop_prflag,
  input  [3:0]  io_pred_bypass_0_bits_uop_pwflag,
  input         io_pred_bypass_0_bits_uop_pflag_busy,
  input  [3:0]  io_pred_bypass_0_bits_uop_stale_pflag,
  input  [3:0]  io_pred_bypass_0_bits_uop_op1_sel,
  input  [3:0]  io_pred_bypass_0_bits_uop_op2_sel,
  input  [5:0]  io_pred_bypass_0_bits_uop_split_num,
  input  [5:0]  io_pred_bypass_0_bits_uop_self_index,
  input  [5:0]  io_pred_bypass_0_bits_uop_rob_inst_idx,
  input  [5:0]  io_pred_bypass_0_bits_uop_address_num,
  input  [6:0]  io_pred_bypass_0_bits_uop_uopc,
  input  [31:0] io_pred_bypass_0_bits_uop_inst,
  input  [31:0] io_pred_bypass_0_bits_uop_debug_inst,
  input         io_pred_bypass_0_bits_uop_is_rvc,
  input  [39:0] io_pred_bypass_0_bits_uop_debug_pc,
  input  [2:0]  io_pred_bypass_0_bits_uop_iq_type,
  input  [9:0]  io_pred_bypass_0_bits_uop_fu_code,
  input  [3:0]  io_pred_bypass_0_bits_uop_ctrl_br_type,
  input  [1:0]  io_pred_bypass_0_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_pred_bypass_0_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_pred_bypass_0_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_pred_bypass_0_bits_uop_ctrl_op_fcn,
  input         io_pred_bypass_0_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_pred_bypass_0_bits_uop_ctrl_csr_cmd,
  input         io_pred_bypass_0_bits_uop_ctrl_is_load,
  input         io_pred_bypass_0_bits_uop_ctrl_is_sta,
  input         io_pred_bypass_0_bits_uop_ctrl_is_std,
  input  [1:0]  io_pred_bypass_0_bits_uop_ctrl_op3_sel,
  input  [1:0]  io_pred_bypass_0_bits_uop_iw_state,
  input         io_pred_bypass_0_bits_uop_iw_p1_poisoned,
  input         io_pred_bypass_0_bits_uop_iw_p2_poisoned,
  input         io_pred_bypass_0_bits_uop_is_br,
  input         io_pred_bypass_0_bits_uop_is_jalr,
  input         io_pred_bypass_0_bits_uop_is_jal,
  input         io_pred_bypass_0_bits_uop_is_sfb,
  input  [11:0] io_pred_bypass_0_bits_uop_br_mask,
  input  [3:0]  io_pred_bypass_0_bits_uop_br_tag,
  input  [4:0]  io_pred_bypass_0_bits_uop_ftq_idx,
  input         io_pred_bypass_0_bits_uop_edge_inst,
  input  [5:0]  io_pred_bypass_0_bits_uop_pc_lob,
  input         io_pred_bypass_0_bits_uop_taken,
  input  [19:0] io_pred_bypass_0_bits_uop_imm_packed,
  input  [11:0] io_pred_bypass_0_bits_uop_csr_addr,
  input  [5:0]  io_pred_bypass_0_bits_uop_rob_idx,
  input  [4:0]  io_pred_bypass_0_bits_uop_ldq_idx,
  input  [4:0]  io_pred_bypass_0_bits_uop_stq_idx,
  input  [1:0]  io_pred_bypass_0_bits_uop_rxq_idx,
  input  [6:0]  io_pred_bypass_0_bits_uop_pdst,
  input  [6:0]  io_pred_bypass_0_bits_uop_prs1,
  input  [6:0]  io_pred_bypass_0_bits_uop_prs2,
  input  [6:0]  io_pred_bypass_0_bits_uop_prs3,
  input  [4:0]  io_pred_bypass_0_bits_uop_ppred,
  input         io_pred_bypass_0_bits_uop_prs1_busy,
  input         io_pred_bypass_0_bits_uop_prs2_busy,
  input         io_pred_bypass_0_bits_uop_prs3_busy,
  input         io_pred_bypass_0_bits_uop_ppred_busy,
  input  [6:0]  io_pred_bypass_0_bits_uop_stale_pdst,
  input         io_pred_bypass_0_bits_uop_exception,
  input  [63:0] io_pred_bypass_0_bits_uop_exc_cause,
  input         io_pred_bypass_0_bits_uop_bypassable,
  input  [4:0]  io_pred_bypass_0_bits_uop_mem_cmd,
  input  [1:0]  io_pred_bypass_0_bits_uop_mem_size,
  input         io_pred_bypass_0_bits_uop_mem_signed,
  input         io_pred_bypass_0_bits_uop_is_fence,
  input         io_pred_bypass_0_bits_uop_is_fencei,
  input         io_pred_bypass_0_bits_uop_is_amo,
  input         io_pred_bypass_0_bits_uop_uses_ldq,
  input         io_pred_bypass_0_bits_uop_uses_stq,
  input         io_pred_bypass_0_bits_uop_is_sys_pc2epc,
  input         io_pred_bypass_0_bits_uop_is_unique,
  input         io_pred_bypass_0_bits_uop_flush_on_commit,
  input         io_pred_bypass_0_bits_uop_ldst_is_rs1,
  input  [5:0]  io_pred_bypass_0_bits_uop_ldst,
  input  [5:0]  io_pred_bypass_0_bits_uop_lrs1,
  input  [5:0]  io_pred_bypass_0_bits_uop_lrs2,
  input  [5:0]  io_pred_bypass_0_bits_uop_lrs3,
  input         io_pred_bypass_0_bits_uop_ldst_val,
  input  [1:0]  io_pred_bypass_0_bits_uop_dst_rtype,
  input  [1:0]  io_pred_bypass_0_bits_uop_lrs1_rtype,
  input  [1:0]  io_pred_bypass_0_bits_uop_lrs2_rtype,
  input         io_pred_bypass_0_bits_uop_frs3_en,
  input         io_pred_bypass_0_bits_uop_fp_val,
  input         io_pred_bypass_0_bits_uop_fp_single,
  input         io_pred_bypass_0_bits_uop_xcpt_pf_if,
  input         io_pred_bypass_0_bits_uop_xcpt_ae_if,
  input         io_pred_bypass_0_bits_uop_xcpt_ma_if,
  input         io_pred_bypass_0_bits_uop_bp_debug_if,
  input         io_pred_bypass_0_bits_uop_bp_xcpt_if,
  input  [1:0]  io_pred_bypass_0_bits_uop_debug_fsrc,
  input  [1:0]  io_pred_bypass_0_bits_uop_debug_tsrc,
  input         io_pred_bypass_0_bits_data,
  input         io_pred_bypass_0_bits_predicated,
  input         io_pred_bypass_0_bits_fflags_valid,
  input         io_pred_bypass_0_bits_fflags_bits_uop_switch,
  input         io_pred_bypass_0_bits_fflags_bits_uop_switch_off,
  input         io_pred_bypass_0_bits_fflags_bits_uop_is_unicore,
  input  [2:0]  io_pred_bypass_0_bits_fflags_bits_uop_shift,
  input  [1:0]  io_pred_bypass_0_bits_fflags_bits_uop_lrs3_rtype,
  input         io_pred_bypass_0_bits_fflags_bits_uop_rflag,
  input         io_pred_bypass_0_bits_fflags_bits_uop_wflag,
  input  [3:0]  io_pred_bypass_0_bits_fflags_bits_uop_prflag,
  input  [3:0]  io_pred_bypass_0_bits_fflags_bits_uop_pwflag,
  input         io_pred_bypass_0_bits_fflags_bits_uop_pflag_busy,
  input  [3:0]  io_pred_bypass_0_bits_fflags_bits_uop_stale_pflag,
  input  [3:0]  io_pred_bypass_0_bits_fflags_bits_uop_op1_sel,
  input  [3:0]  io_pred_bypass_0_bits_fflags_bits_uop_op2_sel,
  input  [5:0]  io_pred_bypass_0_bits_fflags_bits_uop_split_num,
  input  [5:0]  io_pred_bypass_0_bits_fflags_bits_uop_self_index,
  input  [5:0]  io_pred_bypass_0_bits_fflags_bits_uop_rob_inst_idx,
  input  [5:0]  io_pred_bypass_0_bits_fflags_bits_uop_address_num,
  input  [6:0]  io_pred_bypass_0_bits_fflags_bits_uop_uopc,
  input  [31:0] io_pred_bypass_0_bits_fflags_bits_uop_inst,
  input  [31:0] io_pred_bypass_0_bits_fflags_bits_uop_debug_inst,
  input         io_pred_bypass_0_bits_fflags_bits_uop_is_rvc,
  input  [39:0] io_pred_bypass_0_bits_fflags_bits_uop_debug_pc,
  input  [2:0]  io_pred_bypass_0_bits_fflags_bits_uop_iq_type,
  input  [9:0]  io_pred_bypass_0_bits_fflags_bits_uop_fu_code,
  input  [3:0]  io_pred_bypass_0_bits_fflags_bits_uop_ctrl_br_type,
  input  [1:0]  io_pred_bypass_0_bits_fflags_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_pred_bypass_0_bits_fflags_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_pred_bypass_0_bits_fflags_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_pred_bypass_0_bits_fflags_bits_uop_ctrl_op_fcn,
  input         io_pred_bypass_0_bits_fflags_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_pred_bypass_0_bits_fflags_bits_uop_ctrl_csr_cmd,
  input         io_pred_bypass_0_bits_fflags_bits_uop_ctrl_is_load,
  input         io_pred_bypass_0_bits_fflags_bits_uop_ctrl_is_sta,
  input         io_pred_bypass_0_bits_fflags_bits_uop_ctrl_is_std,
  input  [1:0]  io_pred_bypass_0_bits_fflags_bits_uop_ctrl_op3_sel,
  input  [1:0]  io_pred_bypass_0_bits_fflags_bits_uop_iw_state,
  input         io_pred_bypass_0_bits_fflags_bits_uop_iw_p1_poisoned,
  input         io_pred_bypass_0_bits_fflags_bits_uop_iw_p2_poisoned,
  input         io_pred_bypass_0_bits_fflags_bits_uop_is_br,
  input         io_pred_bypass_0_bits_fflags_bits_uop_is_jalr,
  input         io_pred_bypass_0_bits_fflags_bits_uop_is_jal,
  input         io_pred_bypass_0_bits_fflags_bits_uop_is_sfb,
  input  [11:0] io_pred_bypass_0_bits_fflags_bits_uop_br_mask,
  input  [3:0]  io_pred_bypass_0_bits_fflags_bits_uop_br_tag,
  input  [4:0]  io_pred_bypass_0_bits_fflags_bits_uop_ftq_idx,
  input         io_pred_bypass_0_bits_fflags_bits_uop_edge_inst,
  input  [5:0]  io_pred_bypass_0_bits_fflags_bits_uop_pc_lob,
  input         io_pred_bypass_0_bits_fflags_bits_uop_taken,
  input  [19:0] io_pred_bypass_0_bits_fflags_bits_uop_imm_packed,
  input  [11:0] io_pred_bypass_0_bits_fflags_bits_uop_csr_addr,
  input  [5:0]  io_pred_bypass_0_bits_fflags_bits_uop_rob_idx,
  input  [4:0]  io_pred_bypass_0_bits_fflags_bits_uop_ldq_idx,
  input  [4:0]  io_pred_bypass_0_bits_fflags_bits_uop_stq_idx,
  input  [1:0]  io_pred_bypass_0_bits_fflags_bits_uop_rxq_idx,
  input  [6:0]  io_pred_bypass_0_bits_fflags_bits_uop_pdst,
  input  [6:0]  io_pred_bypass_0_bits_fflags_bits_uop_prs1,
  input  [6:0]  io_pred_bypass_0_bits_fflags_bits_uop_prs2,
  input  [6:0]  io_pred_bypass_0_bits_fflags_bits_uop_prs3,
  input  [4:0]  io_pred_bypass_0_bits_fflags_bits_uop_ppred,
  input         io_pred_bypass_0_bits_fflags_bits_uop_prs1_busy,
  input         io_pred_bypass_0_bits_fflags_bits_uop_prs2_busy,
  input         io_pred_bypass_0_bits_fflags_bits_uop_prs3_busy,
  input         io_pred_bypass_0_bits_fflags_bits_uop_ppred_busy,
  input  [6:0]  io_pred_bypass_0_bits_fflags_bits_uop_stale_pdst,
  input         io_pred_bypass_0_bits_fflags_bits_uop_exception,
  input  [63:0] io_pred_bypass_0_bits_fflags_bits_uop_exc_cause,
  input         io_pred_bypass_0_bits_fflags_bits_uop_bypassable,
  input  [4:0]  io_pred_bypass_0_bits_fflags_bits_uop_mem_cmd,
  input  [1:0]  io_pred_bypass_0_bits_fflags_bits_uop_mem_size,
  input         io_pred_bypass_0_bits_fflags_bits_uop_mem_signed,
  input         io_pred_bypass_0_bits_fflags_bits_uop_is_fence,
  input         io_pred_bypass_0_bits_fflags_bits_uop_is_fencei,
  input         io_pred_bypass_0_bits_fflags_bits_uop_is_amo,
  input         io_pred_bypass_0_bits_fflags_bits_uop_uses_ldq,
  input         io_pred_bypass_0_bits_fflags_bits_uop_uses_stq,
  input         io_pred_bypass_0_bits_fflags_bits_uop_is_sys_pc2epc,
  input         io_pred_bypass_0_bits_fflags_bits_uop_is_unique,
  input         io_pred_bypass_0_bits_fflags_bits_uop_flush_on_commit,
  input         io_pred_bypass_0_bits_fflags_bits_uop_ldst_is_rs1,
  input  [5:0]  io_pred_bypass_0_bits_fflags_bits_uop_ldst,
  input  [5:0]  io_pred_bypass_0_bits_fflags_bits_uop_lrs1,
  input  [5:0]  io_pred_bypass_0_bits_fflags_bits_uop_lrs2,
  input  [5:0]  io_pred_bypass_0_bits_fflags_bits_uop_lrs3,
  input         io_pred_bypass_0_bits_fflags_bits_uop_ldst_val,
  input  [1:0]  io_pred_bypass_0_bits_fflags_bits_uop_dst_rtype,
  input  [1:0]  io_pred_bypass_0_bits_fflags_bits_uop_lrs1_rtype,
  input  [1:0]  io_pred_bypass_0_bits_fflags_bits_uop_lrs2_rtype,
  input         io_pred_bypass_0_bits_fflags_bits_uop_frs3_en,
  input         io_pred_bypass_0_bits_fflags_bits_uop_fp_val,
  input         io_pred_bypass_0_bits_fflags_bits_uop_fp_single,
  input         io_pred_bypass_0_bits_fflags_bits_uop_xcpt_pf_if,
  input         io_pred_bypass_0_bits_fflags_bits_uop_xcpt_ae_if,
  input         io_pred_bypass_0_bits_fflags_bits_uop_xcpt_ma_if,
  input         io_pred_bypass_0_bits_fflags_bits_uop_bp_debug_if,
  input         io_pred_bypass_0_bits_fflags_bits_uop_bp_xcpt_if,
  input  [1:0]  io_pred_bypass_0_bits_fflags_bits_uop_debug_fsrc,
  input  [1:0]  io_pred_bypass_0_bits_fflags_bits_uop_debug_tsrc,
  input  [4:0]  io_pred_bypass_0_bits_fflags_bits_flags,
  input  [3:0]  io_pred_bypass_0_bits_flagdata,
  input         io_pred_bypass_0_bits_fflagdata_valid,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_switch,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_switch_off,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_is_unicore,
  input  [2:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_shift,
  input  [1:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_lrs3_rtype,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_rflag,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_wflag,
  input  [3:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_prflag,
  input  [3:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_pwflag,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_pflag_busy,
  input  [3:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_stale_pflag,
  input  [3:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_op1_sel,
  input  [3:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_op2_sel,
  input  [5:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_split_num,
  input  [5:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_self_index,
  input  [5:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_rob_inst_idx,
  input  [5:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_address_num,
  input  [6:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_uopc,
  input  [31:0] io_pred_bypass_0_bits_fflagdata_bits_uop_inst,
  input  [31:0] io_pred_bypass_0_bits_fflagdata_bits_uop_debug_inst,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_is_rvc,
  input  [39:0] io_pred_bypass_0_bits_fflagdata_bits_uop_debug_pc,
  input  [2:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_iq_type,
  input  [9:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_fu_code,
  input  [3:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_ctrl_br_type,
  input  [1:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_ctrl_op_fcn,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_ctrl_csr_cmd,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_ctrl_is_load,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_ctrl_is_sta,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_ctrl_is_std,
  input  [1:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_ctrl_op3_sel,
  input  [1:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_iw_state,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_iw_p1_poisoned,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_iw_p2_poisoned,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_is_br,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_is_jalr,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_is_jal,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_is_sfb,
  input  [11:0] io_pred_bypass_0_bits_fflagdata_bits_uop_br_mask,
  input  [3:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_br_tag,
  input  [4:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_ftq_idx,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_edge_inst,
  input  [5:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_pc_lob,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_taken,
  input  [19:0] io_pred_bypass_0_bits_fflagdata_bits_uop_imm_packed,
  input  [11:0] io_pred_bypass_0_bits_fflagdata_bits_uop_csr_addr,
  input  [5:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_rob_idx,
  input  [4:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_ldq_idx,
  input  [4:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_stq_idx,
  input  [1:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_rxq_idx,
  input  [6:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_pdst,
  input  [6:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_prs1,
  input  [6:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_prs2,
  input  [6:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_prs3,
  input  [4:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_ppred,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_prs1_busy,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_prs2_busy,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_prs3_busy,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_ppred_busy,
  input  [6:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_stale_pdst,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_exception,
  input  [63:0] io_pred_bypass_0_bits_fflagdata_bits_uop_exc_cause,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_bypassable,
  input  [4:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_mem_cmd,
  input  [1:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_mem_size,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_mem_signed,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_is_fence,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_is_fencei,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_is_amo,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_uses_ldq,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_uses_stq,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_is_sys_pc2epc,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_is_unique,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_flush_on_commit,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_ldst_is_rs1,
  input  [5:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_ldst,
  input  [5:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_lrs1,
  input  [5:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_lrs2,
  input  [5:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_lrs3,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_ldst_val,
  input  [1:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_dst_rtype,
  input  [1:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_lrs1_rtype,
  input  [1:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_lrs2_rtype,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_frs3_en,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_fp_val,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_fp_single,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_xcpt_pf_if,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_xcpt_ae_if,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_xcpt_ma_if,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_bp_debug_if,
  input         io_pred_bypass_0_bits_fflagdata_bits_uop_bp_xcpt_if,
  input  [1:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_debug_fsrc,
  input  [1:0]  io_pred_bypass_0_bits_fflagdata_bits_uop_debug_tsrc,
  input  [31:0] io_pred_bypass_0_bits_fflagdata_bits_fflag,
  input         io_pred_bypass_1_valid,
  input         io_pred_bypass_1_bits_uop_switch,
  input         io_pred_bypass_1_bits_uop_switch_off,
  input         io_pred_bypass_1_bits_uop_is_unicore,
  input  [2:0]  io_pred_bypass_1_bits_uop_shift,
  input  [1:0]  io_pred_bypass_1_bits_uop_lrs3_rtype,
  input         io_pred_bypass_1_bits_uop_rflag,
  input         io_pred_bypass_1_bits_uop_wflag,
  input  [3:0]  io_pred_bypass_1_bits_uop_prflag,
  input  [3:0]  io_pred_bypass_1_bits_uop_pwflag,
  input         io_pred_bypass_1_bits_uop_pflag_busy,
  input  [3:0]  io_pred_bypass_1_bits_uop_stale_pflag,
  input  [3:0]  io_pred_bypass_1_bits_uop_op1_sel,
  input  [3:0]  io_pred_bypass_1_bits_uop_op2_sel,
  input  [5:0]  io_pred_bypass_1_bits_uop_split_num,
  input  [5:0]  io_pred_bypass_1_bits_uop_self_index,
  input  [5:0]  io_pred_bypass_1_bits_uop_rob_inst_idx,
  input  [5:0]  io_pred_bypass_1_bits_uop_address_num,
  input  [6:0]  io_pred_bypass_1_bits_uop_uopc,
  input  [31:0] io_pred_bypass_1_bits_uop_inst,
  input  [31:0] io_pred_bypass_1_bits_uop_debug_inst,
  input         io_pred_bypass_1_bits_uop_is_rvc,
  input  [39:0] io_pred_bypass_1_bits_uop_debug_pc,
  input  [2:0]  io_pred_bypass_1_bits_uop_iq_type,
  input  [9:0]  io_pred_bypass_1_bits_uop_fu_code,
  input  [3:0]  io_pred_bypass_1_bits_uop_ctrl_br_type,
  input  [1:0]  io_pred_bypass_1_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_pred_bypass_1_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_pred_bypass_1_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_pred_bypass_1_bits_uop_ctrl_op_fcn,
  input         io_pred_bypass_1_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_pred_bypass_1_bits_uop_ctrl_csr_cmd,
  input         io_pred_bypass_1_bits_uop_ctrl_is_load,
  input         io_pred_bypass_1_bits_uop_ctrl_is_sta,
  input         io_pred_bypass_1_bits_uop_ctrl_is_std,
  input  [1:0]  io_pred_bypass_1_bits_uop_ctrl_op3_sel,
  input  [1:0]  io_pred_bypass_1_bits_uop_iw_state,
  input         io_pred_bypass_1_bits_uop_iw_p1_poisoned,
  input         io_pred_bypass_1_bits_uop_iw_p2_poisoned,
  input         io_pred_bypass_1_bits_uop_is_br,
  input         io_pred_bypass_1_bits_uop_is_jalr,
  input         io_pred_bypass_1_bits_uop_is_jal,
  input         io_pred_bypass_1_bits_uop_is_sfb,
  input  [11:0] io_pred_bypass_1_bits_uop_br_mask,
  input  [3:0]  io_pred_bypass_1_bits_uop_br_tag,
  input  [4:0]  io_pred_bypass_1_bits_uop_ftq_idx,
  input         io_pred_bypass_1_bits_uop_edge_inst,
  input  [5:0]  io_pred_bypass_1_bits_uop_pc_lob,
  input         io_pred_bypass_1_bits_uop_taken,
  input  [19:0] io_pred_bypass_1_bits_uop_imm_packed,
  input  [11:0] io_pred_bypass_1_bits_uop_csr_addr,
  input  [5:0]  io_pred_bypass_1_bits_uop_rob_idx,
  input  [4:0]  io_pred_bypass_1_bits_uop_ldq_idx,
  input  [4:0]  io_pred_bypass_1_bits_uop_stq_idx,
  input  [1:0]  io_pred_bypass_1_bits_uop_rxq_idx,
  input  [6:0]  io_pred_bypass_1_bits_uop_pdst,
  input  [6:0]  io_pred_bypass_1_bits_uop_prs1,
  input  [6:0]  io_pred_bypass_1_bits_uop_prs2,
  input  [6:0]  io_pred_bypass_1_bits_uop_prs3,
  input  [4:0]  io_pred_bypass_1_bits_uop_ppred,
  input         io_pred_bypass_1_bits_uop_prs1_busy,
  input         io_pred_bypass_1_bits_uop_prs2_busy,
  input         io_pred_bypass_1_bits_uop_prs3_busy,
  input         io_pred_bypass_1_bits_uop_ppred_busy,
  input  [6:0]  io_pred_bypass_1_bits_uop_stale_pdst,
  input         io_pred_bypass_1_bits_uop_exception,
  input  [63:0] io_pred_bypass_1_bits_uop_exc_cause,
  input         io_pred_bypass_1_bits_uop_bypassable,
  input  [4:0]  io_pred_bypass_1_bits_uop_mem_cmd,
  input  [1:0]  io_pred_bypass_1_bits_uop_mem_size,
  input         io_pred_bypass_1_bits_uop_mem_signed,
  input         io_pred_bypass_1_bits_uop_is_fence,
  input         io_pred_bypass_1_bits_uop_is_fencei,
  input         io_pred_bypass_1_bits_uop_is_amo,
  input         io_pred_bypass_1_bits_uop_uses_ldq,
  input         io_pred_bypass_1_bits_uop_uses_stq,
  input         io_pred_bypass_1_bits_uop_is_sys_pc2epc,
  input         io_pred_bypass_1_bits_uop_is_unique,
  input         io_pred_bypass_1_bits_uop_flush_on_commit,
  input         io_pred_bypass_1_bits_uop_ldst_is_rs1,
  input  [5:0]  io_pred_bypass_1_bits_uop_ldst,
  input  [5:0]  io_pred_bypass_1_bits_uop_lrs1,
  input  [5:0]  io_pred_bypass_1_bits_uop_lrs2,
  input  [5:0]  io_pred_bypass_1_bits_uop_lrs3,
  input         io_pred_bypass_1_bits_uop_ldst_val,
  input  [1:0]  io_pred_bypass_1_bits_uop_dst_rtype,
  input  [1:0]  io_pred_bypass_1_bits_uop_lrs1_rtype,
  input  [1:0]  io_pred_bypass_1_bits_uop_lrs2_rtype,
  input         io_pred_bypass_1_bits_uop_frs3_en,
  input         io_pred_bypass_1_bits_uop_fp_val,
  input         io_pred_bypass_1_bits_uop_fp_single,
  input         io_pred_bypass_1_bits_uop_xcpt_pf_if,
  input         io_pred_bypass_1_bits_uop_xcpt_ae_if,
  input         io_pred_bypass_1_bits_uop_xcpt_ma_if,
  input         io_pred_bypass_1_bits_uop_bp_debug_if,
  input         io_pred_bypass_1_bits_uop_bp_xcpt_if,
  input  [1:0]  io_pred_bypass_1_bits_uop_debug_fsrc,
  input  [1:0]  io_pred_bypass_1_bits_uop_debug_tsrc,
  input         io_pred_bypass_1_bits_data,
  input         io_pred_bypass_1_bits_predicated,
  input         io_pred_bypass_1_bits_fflags_valid,
  input         io_pred_bypass_1_bits_fflags_bits_uop_switch,
  input         io_pred_bypass_1_bits_fflags_bits_uop_switch_off,
  input         io_pred_bypass_1_bits_fflags_bits_uop_is_unicore,
  input  [2:0]  io_pred_bypass_1_bits_fflags_bits_uop_shift,
  input  [1:0]  io_pred_bypass_1_bits_fflags_bits_uop_lrs3_rtype,
  input         io_pred_bypass_1_bits_fflags_bits_uop_rflag,
  input         io_pred_bypass_1_bits_fflags_bits_uop_wflag,
  input  [3:0]  io_pred_bypass_1_bits_fflags_bits_uop_prflag,
  input  [3:0]  io_pred_bypass_1_bits_fflags_bits_uop_pwflag,
  input         io_pred_bypass_1_bits_fflags_bits_uop_pflag_busy,
  input  [3:0]  io_pred_bypass_1_bits_fflags_bits_uop_stale_pflag,
  input  [3:0]  io_pred_bypass_1_bits_fflags_bits_uop_op1_sel,
  input  [3:0]  io_pred_bypass_1_bits_fflags_bits_uop_op2_sel,
  input  [5:0]  io_pred_bypass_1_bits_fflags_bits_uop_split_num,
  input  [5:0]  io_pred_bypass_1_bits_fflags_bits_uop_self_index,
  input  [5:0]  io_pred_bypass_1_bits_fflags_bits_uop_rob_inst_idx,
  input  [5:0]  io_pred_bypass_1_bits_fflags_bits_uop_address_num,
  input  [6:0]  io_pred_bypass_1_bits_fflags_bits_uop_uopc,
  input  [31:0] io_pred_bypass_1_bits_fflags_bits_uop_inst,
  input  [31:0] io_pred_bypass_1_bits_fflags_bits_uop_debug_inst,
  input         io_pred_bypass_1_bits_fflags_bits_uop_is_rvc,
  input  [39:0] io_pred_bypass_1_bits_fflags_bits_uop_debug_pc,
  input  [2:0]  io_pred_bypass_1_bits_fflags_bits_uop_iq_type,
  input  [9:0]  io_pred_bypass_1_bits_fflags_bits_uop_fu_code,
  input  [3:0]  io_pred_bypass_1_bits_fflags_bits_uop_ctrl_br_type,
  input  [1:0]  io_pred_bypass_1_bits_fflags_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_pred_bypass_1_bits_fflags_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_pred_bypass_1_bits_fflags_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_pred_bypass_1_bits_fflags_bits_uop_ctrl_op_fcn,
  input         io_pred_bypass_1_bits_fflags_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_pred_bypass_1_bits_fflags_bits_uop_ctrl_csr_cmd,
  input         io_pred_bypass_1_bits_fflags_bits_uop_ctrl_is_load,
  input         io_pred_bypass_1_bits_fflags_bits_uop_ctrl_is_sta,
  input         io_pred_bypass_1_bits_fflags_bits_uop_ctrl_is_std,
  input  [1:0]  io_pred_bypass_1_bits_fflags_bits_uop_ctrl_op3_sel,
  input  [1:0]  io_pred_bypass_1_bits_fflags_bits_uop_iw_state,
  input         io_pred_bypass_1_bits_fflags_bits_uop_iw_p1_poisoned,
  input         io_pred_bypass_1_bits_fflags_bits_uop_iw_p2_poisoned,
  input         io_pred_bypass_1_bits_fflags_bits_uop_is_br,
  input         io_pred_bypass_1_bits_fflags_bits_uop_is_jalr,
  input         io_pred_bypass_1_bits_fflags_bits_uop_is_jal,
  input         io_pred_bypass_1_bits_fflags_bits_uop_is_sfb,
  input  [11:0] io_pred_bypass_1_bits_fflags_bits_uop_br_mask,
  input  [3:0]  io_pred_bypass_1_bits_fflags_bits_uop_br_tag,
  input  [4:0]  io_pred_bypass_1_bits_fflags_bits_uop_ftq_idx,
  input         io_pred_bypass_1_bits_fflags_bits_uop_edge_inst,
  input  [5:0]  io_pred_bypass_1_bits_fflags_bits_uop_pc_lob,
  input         io_pred_bypass_1_bits_fflags_bits_uop_taken,
  input  [19:0] io_pred_bypass_1_bits_fflags_bits_uop_imm_packed,
  input  [11:0] io_pred_bypass_1_bits_fflags_bits_uop_csr_addr,
  input  [5:0]  io_pred_bypass_1_bits_fflags_bits_uop_rob_idx,
  input  [4:0]  io_pred_bypass_1_bits_fflags_bits_uop_ldq_idx,
  input  [4:0]  io_pred_bypass_1_bits_fflags_bits_uop_stq_idx,
  input  [1:0]  io_pred_bypass_1_bits_fflags_bits_uop_rxq_idx,
  input  [6:0]  io_pred_bypass_1_bits_fflags_bits_uop_pdst,
  input  [6:0]  io_pred_bypass_1_bits_fflags_bits_uop_prs1,
  input  [6:0]  io_pred_bypass_1_bits_fflags_bits_uop_prs2,
  input  [6:0]  io_pred_bypass_1_bits_fflags_bits_uop_prs3,
  input  [4:0]  io_pred_bypass_1_bits_fflags_bits_uop_ppred,
  input         io_pred_bypass_1_bits_fflags_bits_uop_prs1_busy,
  input         io_pred_bypass_1_bits_fflags_bits_uop_prs2_busy,
  input         io_pred_bypass_1_bits_fflags_bits_uop_prs3_busy,
  input         io_pred_bypass_1_bits_fflags_bits_uop_ppred_busy,
  input  [6:0]  io_pred_bypass_1_bits_fflags_bits_uop_stale_pdst,
  input         io_pred_bypass_1_bits_fflags_bits_uop_exception,
  input  [63:0] io_pred_bypass_1_bits_fflags_bits_uop_exc_cause,
  input         io_pred_bypass_1_bits_fflags_bits_uop_bypassable,
  input  [4:0]  io_pred_bypass_1_bits_fflags_bits_uop_mem_cmd,
  input  [1:0]  io_pred_bypass_1_bits_fflags_bits_uop_mem_size,
  input         io_pred_bypass_1_bits_fflags_bits_uop_mem_signed,
  input         io_pred_bypass_1_bits_fflags_bits_uop_is_fence,
  input         io_pred_bypass_1_bits_fflags_bits_uop_is_fencei,
  input         io_pred_bypass_1_bits_fflags_bits_uop_is_amo,
  input         io_pred_bypass_1_bits_fflags_bits_uop_uses_ldq,
  input         io_pred_bypass_1_bits_fflags_bits_uop_uses_stq,
  input         io_pred_bypass_1_bits_fflags_bits_uop_is_sys_pc2epc,
  input         io_pred_bypass_1_bits_fflags_bits_uop_is_unique,
  input         io_pred_bypass_1_bits_fflags_bits_uop_flush_on_commit,
  input         io_pred_bypass_1_bits_fflags_bits_uop_ldst_is_rs1,
  input  [5:0]  io_pred_bypass_1_bits_fflags_bits_uop_ldst,
  input  [5:0]  io_pred_bypass_1_bits_fflags_bits_uop_lrs1,
  input  [5:0]  io_pred_bypass_1_bits_fflags_bits_uop_lrs2,
  input  [5:0]  io_pred_bypass_1_bits_fflags_bits_uop_lrs3,
  input         io_pred_bypass_1_bits_fflags_bits_uop_ldst_val,
  input  [1:0]  io_pred_bypass_1_bits_fflags_bits_uop_dst_rtype,
  input  [1:0]  io_pred_bypass_1_bits_fflags_bits_uop_lrs1_rtype,
  input  [1:0]  io_pred_bypass_1_bits_fflags_bits_uop_lrs2_rtype,
  input         io_pred_bypass_1_bits_fflags_bits_uop_frs3_en,
  input         io_pred_bypass_1_bits_fflags_bits_uop_fp_val,
  input         io_pred_bypass_1_bits_fflags_bits_uop_fp_single,
  input         io_pred_bypass_1_bits_fflags_bits_uop_xcpt_pf_if,
  input         io_pred_bypass_1_bits_fflags_bits_uop_xcpt_ae_if,
  input         io_pred_bypass_1_bits_fflags_bits_uop_xcpt_ma_if,
  input         io_pred_bypass_1_bits_fflags_bits_uop_bp_debug_if,
  input         io_pred_bypass_1_bits_fflags_bits_uop_bp_xcpt_if,
  input  [1:0]  io_pred_bypass_1_bits_fflags_bits_uop_debug_fsrc,
  input  [1:0]  io_pred_bypass_1_bits_fflags_bits_uop_debug_tsrc,
  input  [4:0]  io_pred_bypass_1_bits_fflags_bits_flags,
  input  [3:0]  io_pred_bypass_1_bits_flagdata,
  input         io_pred_bypass_1_bits_fflagdata_valid,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_switch,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_switch_off,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_is_unicore,
  input  [2:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_shift,
  input  [1:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_lrs3_rtype,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_rflag,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_wflag,
  input  [3:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_prflag,
  input  [3:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_pwflag,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_pflag_busy,
  input  [3:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_stale_pflag,
  input  [3:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_op1_sel,
  input  [3:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_op2_sel,
  input  [5:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_split_num,
  input  [5:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_self_index,
  input  [5:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_rob_inst_idx,
  input  [5:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_address_num,
  input  [6:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_uopc,
  input  [31:0] io_pred_bypass_1_bits_fflagdata_bits_uop_inst,
  input  [31:0] io_pred_bypass_1_bits_fflagdata_bits_uop_debug_inst,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_is_rvc,
  input  [39:0] io_pred_bypass_1_bits_fflagdata_bits_uop_debug_pc,
  input  [2:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_iq_type,
  input  [9:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_fu_code,
  input  [3:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_ctrl_br_type,
  input  [1:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_ctrl_op_fcn,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_ctrl_csr_cmd,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_ctrl_is_load,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_ctrl_is_sta,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_ctrl_is_std,
  input  [1:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_ctrl_op3_sel,
  input  [1:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_iw_state,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_iw_p1_poisoned,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_iw_p2_poisoned,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_is_br,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_is_jalr,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_is_jal,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_is_sfb,
  input  [11:0] io_pred_bypass_1_bits_fflagdata_bits_uop_br_mask,
  input  [3:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_br_tag,
  input  [4:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_ftq_idx,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_edge_inst,
  input  [5:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_pc_lob,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_taken,
  input  [19:0] io_pred_bypass_1_bits_fflagdata_bits_uop_imm_packed,
  input  [11:0] io_pred_bypass_1_bits_fflagdata_bits_uop_csr_addr,
  input  [5:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_rob_idx,
  input  [4:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_ldq_idx,
  input  [4:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_stq_idx,
  input  [1:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_rxq_idx,
  input  [6:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_pdst,
  input  [6:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_prs1,
  input  [6:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_prs2,
  input  [6:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_prs3,
  input  [4:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_ppred,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_prs1_busy,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_prs2_busy,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_prs3_busy,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_ppred_busy,
  input  [6:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_stale_pdst,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_exception,
  input  [63:0] io_pred_bypass_1_bits_fflagdata_bits_uop_exc_cause,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_bypassable,
  input  [4:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_mem_cmd,
  input  [1:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_mem_size,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_mem_signed,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_is_fence,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_is_fencei,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_is_amo,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_uses_ldq,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_uses_stq,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_is_sys_pc2epc,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_is_unique,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_flush_on_commit,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_ldst_is_rs1,
  input  [5:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_ldst,
  input  [5:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_lrs1,
  input  [5:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_lrs2,
  input  [5:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_lrs3,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_ldst_val,
  input  [1:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_dst_rtype,
  input  [1:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_lrs1_rtype,
  input  [1:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_lrs2_rtype,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_frs3_en,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_fp_val,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_fp_single,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_xcpt_pf_if,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_xcpt_ae_if,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_xcpt_ma_if,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_bp_debug_if,
  input         io_pred_bypass_1_bits_fflagdata_bits_uop_bp_xcpt_if,
  input  [1:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_debug_fsrc,
  input  [1:0]  io_pred_bypass_1_bits_fflagdata_bits_uop_debug_tsrc,
  input  [31:0] io_pred_bypass_1_bits_fflagdata_bits_fflag,
  input         io_pred_bypass_2_valid,
  input         io_pred_bypass_2_bits_uop_switch,
  input         io_pred_bypass_2_bits_uop_switch_off,
  input         io_pred_bypass_2_bits_uop_is_unicore,
  input  [2:0]  io_pred_bypass_2_bits_uop_shift,
  input  [1:0]  io_pred_bypass_2_bits_uop_lrs3_rtype,
  input         io_pred_bypass_2_bits_uop_rflag,
  input         io_pred_bypass_2_bits_uop_wflag,
  input  [3:0]  io_pred_bypass_2_bits_uop_prflag,
  input  [3:0]  io_pred_bypass_2_bits_uop_pwflag,
  input         io_pred_bypass_2_bits_uop_pflag_busy,
  input  [3:0]  io_pred_bypass_2_bits_uop_stale_pflag,
  input  [3:0]  io_pred_bypass_2_bits_uop_op1_sel,
  input  [3:0]  io_pred_bypass_2_bits_uop_op2_sel,
  input  [5:0]  io_pred_bypass_2_bits_uop_split_num,
  input  [5:0]  io_pred_bypass_2_bits_uop_self_index,
  input  [5:0]  io_pred_bypass_2_bits_uop_rob_inst_idx,
  input  [5:0]  io_pred_bypass_2_bits_uop_address_num,
  input  [6:0]  io_pred_bypass_2_bits_uop_uopc,
  input  [31:0] io_pred_bypass_2_bits_uop_inst,
  input  [31:0] io_pred_bypass_2_bits_uop_debug_inst,
  input         io_pred_bypass_2_bits_uop_is_rvc,
  input  [39:0] io_pred_bypass_2_bits_uop_debug_pc,
  input  [2:0]  io_pred_bypass_2_bits_uop_iq_type,
  input  [9:0]  io_pred_bypass_2_bits_uop_fu_code,
  input  [3:0]  io_pred_bypass_2_bits_uop_ctrl_br_type,
  input  [1:0]  io_pred_bypass_2_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_pred_bypass_2_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_pred_bypass_2_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_pred_bypass_2_bits_uop_ctrl_op_fcn,
  input         io_pred_bypass_2_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_pred_bypass_2_bits_uop_ctrl_csr_cmd,
  input         io_pred_bypass_2_bits_uop_ctrl_is_load,
  input         io_pred_bypass_2_bits_uop_ctrl_is_sta,
  input         io_pred_bypass_2_bits_uop_ctrl_is_std,
  input  [1:0]  io_pred_bypass_2_bits_uop_ctrl_op3_sel,
  input  [1:0]  io_pred_bypass_2_bits_uop_iw_state,
  input         io_pred_bypass_2_bits_uop_iw_p1_poisoned,
  input         io_pred_bypass_2_bits_uop_iw_p2_poisoned,
  input         io_pred_bypass_2_bits_uop_is_br,
  input         io_pred_bypass_2_bits_uop_is_jalr,
  input         io_pred_bypass_2_bits_uop_is_jal,
  input         io_pred_bypass_2_bits_uop_is_sfb,
  input  [11:0] io_pred_bypass_2_bits_uop_br_mask,
  input  [3:0]  io_pred_bypass_2_bits_uop_br_tag,
  input  [4:0]  io_pred_bypass_2_bits_uop_ftq_idx,
  input         io_pred_bypass_2_bits_uop_edge_inst,
  input  [5:0]  io_pred_bypass_2_bits_uop_pc_lob,
  input         io_pred_bypass_2_bits_uop_taken,
  input  [19:0] io_pred_bypass_2_bits_uop_imm_packed,
  input  [11:0] io_pred_bypass_2_bits_uop_csr_addr,
  input  [5:0]  io_pred_bypass_2_bits_uop_rob_idx,
  input  [4:0]  io_pred_bypass_2_bits_uop_ldq_idx,
  input  [4:0]  io_pred_bypass_2_bits_uop_stq_idx,
  input  [1:0]  io_pred_bypass_2_bits_uop_rxq_idx,
  input  [6:0]  io_pred_bypass_2_bits_uop_pdst,
  input  [6:0]  io_pred_bypass_2_bits_uop_prs1,
  input  [6:0]  io_pred_bypass_2_bits_uop_prs2,
  input  [6:0]  io_pred_bypass_2_bits_uop_prs3,
  input  [4:0]  io_pred_bypass_2_bits_uop_ppred,
  input         io_pred_bypass_2_bits_uop_prs1_busy,
  input         io_pred_bypass_2_bits_uop_prs2_busy,
  input         io_pred_bypass_2_bits_uop_prs3_busy,
  input         io_pred_bypass_2_bits_uop_ppred_busy,
  input  [6:0]  io_pred_bypass_2_bits_uop_stale_pdst,
  input         io_pred_bypass_2_bits_uop_exception,
  input  [63:0] io_pred_bypass_2_bits_uop_exc_cause,
  input         io_pred_bypass_2_bits_uop_bypassable,
  input  [4:0]  io_pred_bypass_2_bits_uop_mem_cmd,
  input  [1:0]  io_pred_bypass_2_bits_uop_mem_size,
  input         io_pred_bypass_2_bits_uop_mem_signed,
  input         io_pred_bypass_2_bits_uop_is_fence,
  input         io_pred_bypass_2_bits_uop_is_fencei,
  input         io_pred_bypass_2_bits_uop_is_amo,
  input         io_pred_bypass_2_bits_uop_uses_ldq,
  input         io_pred_bypass_2_bits_uop_uses_stq,
  input         io_pred_bypass_2_bits_uop_is_sys_pc2epc,
  input         io_pred_bypass_2_bits_uop_is_unique,
  input         io_pred_bypass_2_bits_uop_flush_on_commit,
  input         io_pred_bypass_2_bits_uop_ldst_is_rs1,
  input  [5:0]  io_pred_bypass_2_bits_uop_ldst,
  input  [5:0]  io_pred_bypass_2_bits_uop_lrs1,
  input  [5:0]  io_pred_bypass_2_bits_uop_lrs2,
  input  [5:0]  io_pred_bypass_2_bits_uop_lrs3,
  input         io_pred_bypass_2_bits_uop_ldst_val,
  input  [1:0]  io_pred_bypass_2_bits_uop_dst_rtype,
  input  [1:0]  io_pred_bypass_2_bits_uop_lrs1_rtype,
  input  [1:0]  io_pred_bypass_2_bits_uop_lrs2_rtype,
  input         io_pred_bypass_2_bits_uop_frs3_en,
  input         io_pred_bypass_2_bits_uop_fp_val,
  input         io_pred_bypass_2_bits_uop_fp_single,
  input         io_pred_bypass_2_bits_uop_xcpt_pf_if,
  input         io_pred_bypass_2_bits_uop_xcpt_ae_if,
  input         io_pred_bypass_2_bits_uop_xcpt_ma_if,
  input         io_pred_bypass_2_bits_uop_bp_debug_if,
  input         io_pred_bypass_2_bits_uop_bp_xcpt_if,
  input  [1:0]  io_pred_bypass_2_bits_uop_debug_fsrc,
  input  [1:0]  io_pred_bypass_2_bits_uop_debug_tsrc,
  input         io_pred_bypass_2_bits_data,
  input         io_pred_bypass_2_bits_predicated,
  input         io_pred_bypass_2_bits_fflags_valid,
  input         io_pred_bypass_2_bits_fflags_bits_uop_switch,
  input         io_pred_bypass_2_bits_fflags_bits_uop_switch_off,
  input         io_pred_bypass_2_bits_fflags_bits_uop_is_unicore,
  input  [2:0]  io_pred_bypass_2_bits_fflags_bits_uop_shift,
  input  [1:0]  io_pred_bypass_2_bits_fflags_bits_uop_lrs3_rtype,
  input         io_pred_bypass_2_bits_fflags_bits_uop_rflag,
  input         io_pred_bypass_2_bits_fflags_bits_uop_wflag,
  input  [3:0]  io_pred_bypass_2_bits_fflags_bits_uop_prflag,
  input  [3:0]  io_pred_bypass_2_bits_fflags_bits_uop_pwflag,
  input         io_pred_bypass_2_bits_fflags_bits_uop_pflag_busy,
  input  [3:0]  io_pred_bypass_2_bits_fflags_bits_uop_stale_pflag,
  input  [3:0]  io_pred_bypass_2_bits_fflags_bits_uop_op1_sel,
  input  [3:0]  io_pred_bypass_2_bits_fflags_bits_uop_op2_sel,
  input  [5:0]  io_pred_bypass_2_bits_fflags_bits_uop_split_num,
  input  [5:0]  io_pred_bypass_2_bits_fflags_bits_uop_self_index,
  input  [5:0]  io_pred_bypass_2_bits_fflags_bits_uop_rob_inst_idx,
  input  [5:0]  io_pred_bypass_2_bits_fflags_bits_uop_address_num,
  input  [6:0]  io_pred_bypass_2_bits_fflags_bits_uop_uopc,
  input  [31:0] io_pred_bypass_2_bits_fflags_bits_uop_inst,
  input  [31:0] io_pred_bypass_2_bits_fflags_bits_uop_debug_inst,
  input         io_pred_bypass_2_bits_fflags_bits_uop_is_rvc,
  input  [39:0] io_pred_bypass_2_bits_fflags_bits_uop_debug_pc,
  input  [2:0]  io_pred_bypass_2_bits_fflags_bits_uop_iq_type,
  input  [9:0]  io_pred_bypass_2_bits_fflags_bits_uop_fu_code,
  input  [3:0]  io_pred_bypass_2_bits_fflags_bits_uop_ctrl_br_type,
  input  [1:0]  io_pred_bypass_2_bits_fflags_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_pred_bypass_2_bits_fflags_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_pred_bypass_2_bits_fflags_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_pred_bypass_2_bits_fflags_bits_uop_ctrl_op_fcn,
  input         io_pred_bypass_2_bits_fflags_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_pred_bypass_2_bits_fflags_bits_uop_ctrl_csr_cmd,
  input         io_pred_bypass_2_bits_fflags_bits_uop_ctrl_is_load,
  input         io_pred_bypass_2_bits_fflags_bits_uop_ctrl_is_sta,
  input         io_pred_bypass_2_bits_fflags_bits_uop_ctrl_is_std,
  input  [1:0]  io_pred_bypass_2_bits_fflags_bits_uop_ctrl_op3_sel,
  input  [1:0]  io_pred_bypass_2_bits_fflags_bits_uop_iw_state,
  input         io_pred_bypass_2_bits_fflags_bits_uop_iw_p1_poisoned,
  input         io_pred_bypass_2_bits_fflags_bits_uop_iw_p2_poisoned,
  input         io_pred_bypass_2_bits_fflags_bits_uop_is_br,
  input         io_pred_bypass_2_bits_fflags_bits_uop_is_jalr,
  input         io_pred_bypass_2_bits_fflags_bits_uop_is_jal,
  input         io_pred_bypass_2_bits_fflags_bits_uop_is_sfb,
  input  [11:0] io_pred_bypass_2_bits_fflags_bits_uop_br_mask,
  input  [3:0]  io_pred_bypass_2_bits_fflags_bits_uop_br_tag,
  input  [4:0]  io_pred_bypass_2_bits_fflags_bits_uop_ftq_idx,
  input         io_pred_bypass_2_bits_fflags_bits_uop_edge_inst,
  input  [5:0]  io_pred_bypass_2_bits_fflags_bits_uop_pc_lob,
  input         io_pred_bypass_2_bits_fflags_bits_uop_taken,
  input  [19:0] io_pred_bypass_2_bits_fflags_bits_uop_imm_packed,
  input  [11:0] io_pred_bypass_2_bits_fflags_bits_uop_csr_addr,
  input  [5:0]  io_pred_bypass_2_bits_fflags_bits_uop_rob_idx,
  input  [4:0]  io_pred_bypass_2_bits_fflags_bits_uop_ldq_idx,
  input  [4:0]  io_pred_bypass_2_bits_fflags_bits_uop_stq_idx,
  input  [1:0]  io_pred_bypass_2_bits_fflags_bits_uop_rxq_idx,
  input  [6:0]  io_pred_bypass_2_bits_fflags_bits_uop_pdst,
  input  [6:0]  io_pred_bypass_2_bits_fflags_bits_uop_prs1,
  input  [6:0]  io_pred_bypass_2_bits_fflags_bits_uop_prs2,
  input  [6:0]  io_pred_bypass_2_bits_fflags_bits_uop_prs3,
  input  [4:0]  io_pred_bypass_2_bits_fflags_bits_uop_ppred,
  input         io_pred_bypass_2_bits_fflags_bits_uop_prs1_busy,
  input         io_pred_bypass_2_bits_fflags_bits_uop_prs2_busy,
  input         io_pred_bypass_2_bits_fflags_bits_uop_prs3_busy,
  input         io_pred_bypass_2_bits_fflags_bits_uop_ppred_busy,
  input  [6:0]  io_pred_bypass_2_bits_fflags_bits_uop_stale_pdst,
  input         io_pred_bypass_2_bits_fflags_bits_uop_exception,
  input  [63:0] io_pred_bypass_2_bits_fflags_bits_uop_exc_cause,
  input         io_pred_bypass_2_bits_fflags_bits_uop_bypassable,
  input  [4:0]  io_pred_bypass_2_bits_fflags_bits_uop_mem_cmd,
  input  [1:0]  io_pred_bypass_2_bits_fflags_bits_uop_mem_size,
  input         io_pred_bypass_2_bits_fflags_bits_uop_mem_signed,
  input         io_pred_bypass_2_bits_fflags_bits_uop_is_fence,
  input         io_pred_bypass_2_bits_fflags_bits_uop_is_fencei,
  input         io_pred_bypass_2_bits_fflags_bits_uop_is_amo,
  input         io_pred_bypass_2_bits_fflags_bits_uop_uses_ldq,
  input         io_pred_bypass_2_bits_fflags_bits_uop_uses_stq,
  input         io_pred_bypass_2_bits_fflags_bits_uop_is_sys_pc2epc,
  input         io_pred_bypass_2_bits_fflags_bits_uop_is_unique,
  input         io_pred_bypass_2_bits_fflags_bits_uop_flush_on_commit,
  input         io_pred_bypass_2_bits_fflags_bits_uop_ldst_is_rs1,
  input  [5:0]  io_pred_bypass_2_bits_fflags_bits_uop_ldst,
  input  [5:0]  io_pred_bypass_2_bits_fflags_bits_uop_lrs1,
  input  [5:0]  io_pred_bypass_2_bits_fflags_bits_uop_lrs2,
  input  [5:0]  io_pred_bypass_2_bits_fflags_bits_uop_lrs3,
  input         io_pred_bypass_2_bits_fflags_bits_uop_ldst_val,
  input  [1:0]  io_pred_bypass_2_bits_fflags_bits_uop_dst_rtype,
  input  [1:0]  io_pred_bypass_2_bits_fflags_bits_uop_lrs1_rtype,
  input  [1:0]  io_pred_bypass_2_bits_fflags_bits_uop_lrs2_rtype,
  input         io_pred_bypass_2_bits_fflags_bits_uop_frs3_en,
  input         io_pred_bypass_2_bits_fflags_bits_uop_fp_val,
  input         io_pred_bypass_2_bits_fflags_bits_uop_fp_single,
  input         io_pred_bypass_2_bits_fflags_bits_uop_xcpt_pf_if,
  input         io_pred_bypass_2_bits_fflags_bits_uop_xcpt_ae_if,
  input         io_pred_bypass_2_bits_fflags_bits_uop_xcpt_ma_if,
  input         io_pred_bypass_2_bits_fflags_bits_uop_bp_debug_if,
  input         io_pred_bypass_2_bits_fflags_bits_uop_bp_xcpt_if,
  input  [1:0]  io_pred_bypass_2_bits_fflags_bits_uop_debug_fsrc,
  input  [1:0]  io_pred_bypass_2_bits_fflags_bits_uop_debug_tsrc,
  input  [4:0]  io_pred_bypass_2_bits_fflags_bits_flags,
  input  [3:0]  io_pred_bypass_2_bits_flagdata,
  input         io_pred_bypass_2_bits_fflagdata_valid,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_switch,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_switch_off,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_is_unicore,
  input  [2:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_shift,
  input  [1:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_lrs3_rtype,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_rflag,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_wflag,
  input  [3:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_prflag,
  input  [3:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_pwflag,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_pflag_busy,
  input  [3:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_stale_pflag,
  input  [3:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_op1_sel,
  input  [3:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_op2_sel,
  input  [5:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_split_num,
  input  [5:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_self_index,
  input  [5:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_rob_inst_idx,
  input  [5:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_address_num,
  input  [6:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_uopc,
  input  [31:0] io_pred_bypass_2_bits_fflagdata_bits_uop_inst,
  input  [31:0] io_pred_bypass_2_bits_fflagdata_bits_uop_debug_inst,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_is_rvc,
  input  [39:0] io_pred_bypass_2_bits_fflagdata_bits_uop_debug_pc,
  input  [2:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_iq_type,
  input  [9:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_fu_code,
  input  [3:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_ctrl_br_type,
  input  [1:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_ctrl_op2_sel,
  input  [2:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_ctrl_op_fcn,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_ctrl_fcn_dw,
  input  [2:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_ctrl_csr_cmd,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_ctrl_is_load,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_ctrl_is_sta,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_ctrl_is_std,
  input  [1:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_ctrl_op3_sel,
  input  [1:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_iw_state,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_iw_p1_poisoned,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_iw_p2_poisoned,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_is_br,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_is_jalr,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_is_jal,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_is_sfb,
  input  [11:0] io_pred_bypass_2_bits_fflagdata_bits_uop_br_mask,
  input  [3:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_br_tag,
  input  [4:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_ftq_idx,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_edge_inst,
  input  [5:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_pc_lob,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_taken,
  input  [19:0] io_pred_bypass_2_bits_fflagdata_bits_uop_imm_packed,
  input  [11:0] io_pred_bypass_2_bits_fflagdata_bits_uop_csr_addr,
  input  [5:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_rob_idx,
  input  [4:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_ldq_idx,
  input  [4:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_stq_idx,
  input  [1:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_rxq_idx,
  input  [6:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_pdst,
  input  [6:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_prs1,
  input  [6:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_prs2,
  input  [6:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_prs3,
  input  [4:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_ppred,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_prs1_busy,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_prs2_busy,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_prs3_busy,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_ppred_busy,
  input  [6:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_stale_pdst,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_exception,
  input  [63:0] io_pred_bypass_2_bits_fflagdata_bits_uop_exc_cause,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_bypassable,
  input  [4:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_mem_cmd,
  input  [1:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_mem_size,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_mem_signed,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_is_fence,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_is_fencei,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_is_amo,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_uses_ldq,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_uses_stq,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_is_sys_pc2epc,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_is_unique,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_flush_on_commit,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_ldst_is_rs1,
  input  [5:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_ldst,
  input  [5:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_lrs1,
  input  [5:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_lrs2,
  input  [5:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_lrs3,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_ldst_val,
  input  [1:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_dst_rtype,
  input  [1:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_lrs1_rtype,
  input  [1:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_lrs2_rtype,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_frs3_en,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_fp_val,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_fp_single,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_xcpt_pf_if,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_xcpt_ae_if,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_xcpt_ma_if,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_bp_debug_if,
  input         io_pred_bypass_2_bits_fflagdata_bits_uop_bp_xcpt_if,
  input  [1:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_debug_fsrc,
  input  [1:0]  io_pred_bypass_2_bits_fflagdata_bits_uop_debug_tsrc,
  input  [31:0] io_pred_bypass_2_bits_fflagdata_bits_fflag,
  input         io_exe_reqs_0_ready,
  output        io_exe_reqs_0_valid,
  output        io_exe_reqs_0_bits_uop_switch,
  output        io_exe_reqs_0_bits_uop_switch_off,
  output        io_exe_reqs_0_bits_uop_is_unicore,
  output [2:0]  io_exe_reqs_0_bits_uop_shift,
  output [1:0]  io_exe_reqs_0_bits_uop_lrs3_rtype,
  output        io_exe_reqs_0_bits_uop_rflag,
  output        io_exe_reqs_0_bits_uop_wflag,
  output [3:0]  io_exe_reqs_0_bits_uop_prflag,
  output [3:0]  io_exe_reqs_0_bits_uop_pwflag,
  output        io_exe_reqs_0_bits_uop_pflag_busy,
  output [3:0]  io_exe_reqs_0_bits_uop_stale_pflag,
  output [3:0]  io_exe_reqs_0_bits_uop_op1_sel,
  output [3:0]  io_exe_reqs_0_bits_uop_op2_sel,
  output [5:0]  io_exe_reqs_0_bits_uop_split_num,
  output [5:0]  io_exe_reqs_0_bits_uop_self_index,
  output [5:0]  io_exe_reqs_0_bits_uop_rob_inst_idx,
  output [5:0]  io_exe_reqs_0_bits_uop_address_num,
  output [6:0]  io_exe_reqs_0_bits_uop_uopc,
  output [31:0] io_exe_reqs_0_bits_uop_inst,
  output [31:0] io_exe_reqs_0_bits_uop_debug_inst,
  output        io_exe_reqs_0_bits_uop_is_rvc,
  output [39:0] io_exe_reqs_0_bits_uop_debug_pc,
  output [2:0]  io_exe_reqs_0_bits_uop_iq_type,
  output [9:0]  io_exe_reqs_0_bits_uop_fu_code,
  output [3:0]  io_exe_reqs_0_bits_uop_ctrl_br_type,
  output [1:0]  io_exe_reqs_0_bits_uop_ctrl_op1_sel,
  output [2:0]  io_exe_reqs_0_bits_uop_ctrl_op2_sel,
  output [2:0]  io_exe_reqs_0_bits_uop_ctrl_imm_sel,
  output [3:0]  io_exe_reqs_0_bits_uop_ctrl_op_fcn,
  output        io_exe_reqs_0_bits_uop_ctrl_fcn_dw,
  output [2:0]  io_exe_reqs_0_bits_uop_ctrl_csr_cmd,
  output        io_exe_reqs_0_bits_uop_ctrl_is_load,
  output        io_exe_reqs_0_bits_uop_ctrl_is_sta,
  output        io_exe_reqs_0_bits_uop_ctrl_is_std,
  output [1:0]  io_exe_reqs_0_bits_uop_ctrl_op3_sel,
  output [1:0]  io_exe_reqs_0_bits_uop_iw_state,
  output        io_exe_reqs_0_bits_uop_iw_p1_poisoned,
  output        io_exe_reqs_0_bits_uop_iw_p2_poisoned,
  output        io_exe_reqs_0_bits_uop_is_br,
  output        io_exe_reqs_0_bits_uop_is_jalr,
  output        io_exe_reqs_0_bits_uop_is_jal,
  output        io_exe_reqs_0_bits_uop_is_sfb,
  output [11:0] io_exe_reqs_0_bits_uop_br_mask,
  output [3:0]  io_exe_reqs_0_bits_uop_br_tag,
  output [4:0]  io_exe_reqs_0_bits_uop_ftq_idx,
  output        io_exe_reqs_0_bits_uop_edge_inst,
  output [5:0]  io_exe_reqs_0_bits_uop_pc_lob,
  output        io_exe_reqs_0_bits_uop_taken,
  output [19:0] io_exe_reqs_0_bits_uop_imm_packed,
  output [11:0] io_exe_reqs_0_bits_uop_csr_addr,
  output [5:0]  io_exe_reqs_0_bits_uop_rob_idx,
  output [4:0]  io_exe_reqs_0_bits_uop_ldq_idx,
  output [4:0]  io_exe_reqs_0_bits_uop_stq_idx,
  output [1:0]  io_exe_reqs_0_bits_uop_rxq_idx,
  output [6:0]  io_exe_reqs_0_bits_uop_pdst,
  output [6:0]  io_exe_reqs_0_bits_uop_prs1,
  output [6:0]  io_exe_reqs_0_bits_uop_prs2,
  output [6:0]  io_exe_reqs_0_bits_uop_prs3,
  output [4:0]  io_exe_reqs_0_bits_uop_ppred,
  output        io_exe_reqs_0_bits_uop_prs1_busy,
  output        io_exe_reqs_0_bits_uop_prs2_busy,
  output        io_exe_reqs_0_bits_uop_prs3_busy,
  output        io_exe_reqs_0_bits_uop_ppred_busy,
  output [6:0]  io_exe_reqs_0_bits_uop_stale_pdst,
  output        io_exe_reqs_0_bits_uop_exception,
  output [63:0] io_exe_reqs_0_bits_uop_exc_cause,
  output        io_exe_reqs_0_bits_uop_bypassable,
  output [4:0]  io_exe_reqs_0_bits_uop_mem_cmd,
  output [1:0]  io_exe_reqs_0_bits_uop_mem_size,
  output        io_exe_reqs_0_bits_uop_mem_signed,
  output        io_exe_reqs_0_bits_uop_is_fence,
  output        io_exe_reqs_0_bits_uop_is_fencei,
  output        io_exe_reqs_0_bits_uop_is_amo,
  output        io_exe_reqs_0_bits_uop_uses_ldq,
  output        io_exe_reqs_0_bits_uop_uses_stq,
  output        io_exe_reqs_0_bits_uop_is_sys_pc2epc,
  output        io_exe_reqs_0_bits_uop_is_unique,
  output        io_exe_reqs_0_bits_uop_flush_on_commit,
  output        io_exe_reqs_0_bits_uop_ldst_is_rs1,
  output [5:0]  io_exe_reqs_0_bits_uop_ldst,
  output [5:0]  io_exe_reqs_0_bits_uop_lrs1,
  output [5:0]  io_exe_reqs_0_bits_uop_lrs2,
  output [5:0]  io_exe_reqs_0_bits_uop_lrs3,
  output        io_exe_reqs_0_bits_uop_ldst_val,
  output [1:0]  io_exe_reqs_0_bits_uop_dst_rtype,
  output [1:0]  io_exe_reqs_0_bits_uop_lrs1_rtype,
  output [1:0]  io_exe_reqs_0_bits_uop_lrs2_rtype,
  output        io_exe_reqs_0_bits_uop_frs3_en,
  output        io_exe_reqs_0_bits_uop_fp_val,
  output        io_exe_reqs_0_bits_uop_fp_single,
  output        io_exe_reqs_0_bits_uop_xcpt_pf_if,
  output        io_exe_reqs_0_bits_uop_xcpt_ae_if,
  output        io_exe_reqs_0_bits_uop_xcpt_ma_if,
  output        io_exe_reqs_0_bits_uop_bp_debug_if,
  output        io_exe_reqs_0_bits_uop_bp_xcpt_if,
  output [1:0]  io_exe_reqs_0_bits_uop_debug_fsrc,
  output [1:0]  io_exe_reqs_0_bits_uop_debug_tsrc,
  output [63:0] io_exe_reqs_0_bits_rs1_data,
  output [63:0] io_exe_reqs_0_bits_rs2_data,
  output [63:0] io_exe_reqs_0_bits_rs3_data,
  output        io_exe_reqs_0_bits_pred_data,
  output [3:0]  io_exe_reqs_0_bits_flagdata,
  output [31:0] io_exe_reqs_0_bits_fflagdata,
  output        io_exe_reqs_0_bits_kill,
  input         io_exe_reqs_1_ready,
  output        io_exe_reqs_1_valid,
  output        io_exe_reqs_1_bits_uop_switch,
  output        io_exe_reqs_1_bits_uop_switch_off,
  output        io_exe_reqs_1_bits_uop_is_unicore,
  output [2:0]  io_exe_reqs_1_bits_uop_shift,
  output [1:0]  io_exe_reqs_1_bits_uop_lrs3_rtype,
  output        io_exe_reqs_1_bits_uop_rflag,
  output        io_exe_reqs_1_bits_uop_wflag,
  output [3:0]  io_exe_reqs_1_bits_uop_prflag,
  output [3:0]  io_exe_reqs_1_bits_uop_pwflag,
  output        io_exe_reqs_1_bits_uop_pflag_busy,
  output [3:0]  io_exe_reqs_1_bits_uop_stale_pflag,
  output [3:0]  io_exe_reqs_1_bits_uop_op1_sel,
  output [3:0]  io_exe_reqs_1_bits_uop_op2_sel,
  output [5:0]  io_exe_reqs_1_bits_uop_split_num,
  output [5:0]  io_exe_reqs_1_bits_uop_self_index,
  output [5:0]  io_exe_reqs_1_bits_uop_rob_inst_idx,
  output [5:0]  io_exe_reqs_1_bits_uop_address_num,
  output [6:0]  io_exe_reqs_1_bits_uop_uopc,
  output [31:0] io_exe_reqs_1_bits_uop_inst,
  output [31:0] io_exe_reqs_1_bits_uop_debug_inst,
  output        io_exe_reqs_1_bits_uop_is_rvc,
  output [39:0] io_exe_reqs_1_bits_uop_debug_pc,
  output [2:0]  io_exe_reqs_1_bits_uop_iq_type,
  output [9:0]  io_exe_reqs_1_bits_uop_fu_code,
  output [3:0]  io_exe_reqs_1_bits_uop_ctrl_br_type,
  output [1:0]  io_exe_reqs_1_bits_uop_ctrl_op1_sel,
  output [2:0]  io_exe_reqs_1_bits_uop_ctrl_op2_sel,
  output [2:0]  io_exe_reqs_1_bits_uop_ctrl_imm_sel,
  output [3:0]  io_exe_reqs_1_bits_uop_ctrl_op_fcn,
  output        io_exe_reqs_1_bits_uop_ctrl_fcn_dw,
  output [2:0]  io_exe_reqs_1_bits_uop_ctrl_csr_cmd,
  output        io_exe_reqs_1_bits_uop_ctrl_is_load,
  output        io_exe_reqs_1_bits_uop_ctrl_is_sta,
  output        io_exe_reqs_1_bits_uop_ctrl_is_std,
  output [1:0]  io_exe_reqs_1_bits_uop_ctrl_op3_sel,
  output [1:0]  io_exe_reqs_1_bits_uop_iw_state,
  output        io_exe_reqs_1_bits_uop_iw_p1_poisoned,
  output        io_exe_reqs_1_bits_uop_iw_p2_poisoned,
  output        io_exe_reqs_1_bits_uop_is_br,
  output        io_exe_reqs_1_bits_uop_is_jalr,
  output        io_exe_reqs_1_bits_uop_is_jal,
  output        io_exe_reqs_1_bits_uop_is_sfb,
  output [11:0] io_exe_reqs_1_bits_uop_br_mask,
  output [3:0]  io_exe_reqs_1_bits_uop_br_tag,
  output [4:0]  io_exe_reqs_1_bits_uop_ftq_idx,
  output        io_exe_reqs_1_bits_uop_edge_inst,
  output [5:0]  io_exe_reqs_1_bits_uop_pc_lob,
  output        io_exe_reqs_1_bits_uop_taken,
  output [19:0] io_exe_reqs_1_bits_uop_imm_packed,
  output [11:0] io_exe_reqs_1_bits_uop_csr_addr,
  output [5:0]  io_exe_reqs_1_bits_uop_rob_idx,
  output [4:0]  io_exe_reqs_1_bits_uop_ldq_idx,
  output [4:0]  io_exe_reqs_1_bits_uop_stq_idx,
  output [1:0]  io_exe_reqs_1_bits_uop_rxq_idx,
  output [6:0]  io_exe_reqs_1_bits_uop_pdst,
  output [6:0]  io_exe_reqs_1_bits_uop_prs1,
  output [6:0]  io_exe_reqs_1_bits_uop_prs2,
  output [6:0]  io_exe_reqs_1_bits_uop_prs3,
  output [4:0]  io_exe_reqs_1_bits_uop_ppred,
  output        io_exe_reqs_1_bits_uop_prs1_busy,
  output        io_exe_reqs_1_bits_uop_prs2_busy,
  output        io_exe_reqs_1_bits_uop_prs3_busy,
  output        io_exe_reqs_1_bits_uop_ppred_busy,
  output [6:0]  io_exe_reqs_1_bits_uop_stale_pdst,
  output        io_exe_reqs_1_bits_uop_exception,
  output [63:0] io_exe_reqs_1_bits_uop_exc_cause,
  output        io_exe_reqs_1_bits_uop_bypassable,
  output [4:0]  io_exe_reqs_1_bits_uop_mem_cmd,
  output [1:0]  io_exe_reqs_1_bits_uop_mem_size,
  output        io_exe_reqs_1_bits_uop_mem_signed,
  output        io_exe_reqs_1_bits_uop_is_fence,
  output        io_exe_reqs_1_bits_uop_is_fencei,
  output        io_exe_reqs_1_bits_uop_is_amo,
  output        io_exe_reqs_1_bits_uop_uses_ldq,
  output        io_exe_reqs_1_bits_uop_uses_stq,
  output        io_exe_reqs_1_bits_uop_is_sys_pc2epc,
  output        io_exe_reqs_1_bits_uop_is_unique,
  output        io_exe_reqs_1_bits_uop_flush_on_commit,
  output        io_exe_reqs_1_bits_uop_ldst_is_rs1,
  output [5:0]  io_exe_reqs_1_bits_uop_ldst,
  output [5:0]  io_exe_reqs_1_bits_uop_lrs1,
  output [5:0]  io_exe_reqs_1_bits_uop_lrs2,
  output [5:0]  io_exe_reqs_1_bits_uop_lrs3,
  output        io_exe_reqs_1_bits_uop_ldst_val,
  output [1:0]  io_exe_reqs_1_bits_uop_dst_rtype,
  output [1:0]  io_exe_reqs_1_bits_uop_lrs1_rtype,
  output [1:0]  io_exe_reqs_1_bits_uop_lrs2_rtype,
  output        io_exe_reqs_1_bits_uop_frs3_en,
  output        io_exe_reqs_1_bits_uop_fp_val,
  output        io_exe_reqs_1_bits_uop_fp_single,
  output        io_exe_reqs_1_bits_uop_xcpt_pf_if,
  output        io_exe_reqs_1_bits_uop_xcpt_ae_if,
  output        io_exe_reqs_1_bits_uop_xcpt_ma_if,
  output        io_exe_reqs_1_bits_uop_bp_debug_if,
  output        io_exe_reqs_1_bits_uop_bp_xcpt_if,
  output [1:0]  io_exe_reqs_1_bits_uop_debug_fsrc,
  output [1:0]  io_exe_reqs_1_bits_uop_debug_tsrc,
  output [63:0] io_exe_reqs_1_bits_rs1_data,
  output [63:0] io_exe_reqs_1_bits_rs2_data,
  output [63:0] io_exe_reqs_1_bits_rs3_data,
  output        io_exe_reqs_1_bits_pred_data,
  output [3:0]  io_exe_reqs_1_bits_flagdata,
  output [31:0] io_exe_reqs_1_bits_fflagdata,
  output        io_exe_reqs_1_bits_kill,
  input         io_exe_reqs_2_ready,
  output        io_exe_reqs_2_valid,
  output        io_exe_reqs_2_bits_uop_switch,
  output        io_exe_reqs_2_bits_uop_switch_off,
  output        io_exe_reqs_2_bits_uop_is_unicore,
  output [2:0]  io_exe_reqs_2_bits_uop_shift,
  output [1:0]  io_exe_reqs_2_bits_uop_lrs3_rtype,
  output        io_exe_reqs_2_bits_uop_rflag,
  output        io_exe_reqs_2_bits_uop_wflag,
  output [3:0]  io_exe_reqs_2_bits_uop_prflag,
  output [3:0]  io_exe_reqs_2_bits_uop_pwflag,
  output        io_exe_reqs_2_bits_uop_pflag_busy,
  output [3:0]  io_exe_reqs_2_bits_uop_stale_pflag,
  output [3:0]  io_exe_reqs_2_bits_uop_op1_sel,
  output [3:0]  io_exe_reqs_2_bits_uop_op2_sel,
  output [5:0]  io_exe_reqs_2_bits_uop_split_num,
  output [5:0]  io_exe_reqs_2_bits_uop_self_index,
  output [5:0]  io_exe_reqs_2_bits_uop_rob_inst_idx,
  output [5:0]  io_exe_reqs_2_bits_uop_address_num,
  output [6:0]  io_exe_reqs_2_bits_uop_uopc,
  output [31:0] io_exe_reqs_2_bits_uop_inst,
  output [31:0] io_exe_reqs_2_bits_uop_debug_inst,
  output        io_exe_reqs_2_bits_uop_is_rvc,
  output [39:0] io_exe_reqs_2_bits_uop_debug_pc,
  output [2:0]  io_exe_reqs_2_bits_uop_iq_type,
  output [9:0]  io_exe_reqs_2_bits_uop_fu_code,
  output [3:0]  io_exe_reqs_2_bits_uop_ctrl_br_type,
  output [1:0]  io_exe_reqs_2_bits_uop_ctrl_op1_sel,
  output [2:0]  io_exe_reqs_2_bits_uop_ctrl_op2_sel,
  output [2:0]  io_exe_reqs_2_bits_uop_ctrl_imm_sel,
  output [3:0]  io_exe_reqs_2_bits_uop_ctrl_op_fcn,
  output        io_exe_reqs_2_bits_uop_ctrl_fcn_dw,
  output [2:0]  io_exe_reqs_2_bits_uop_ctrl_csr_cmd,
  output        io_exe_reqs_2_bits_uop_ctrl_is_load,
  output        io_exe_reqs_2_bits_uop_ctrl_is_sta,
  output        io_exe_reqs_2_bits_uop_ctrl_is_std,
  output [1:0]  io_exe_reqs_2_bits_uop_ctrl_op3_sel,
  output [1:0]  io_exe_reqs_2_bits_uop_iw_state,
  output        io_exe_reqs_2_bits_uop_iw_p1_poisoned,
  output        io_exe_reqs_2_bits_uop_iw_p2_poisoned,
  output        io_exe_reqs_2_bits_uop_is_br,
  output        io_exe_reqs_2_bits_uop_is_jalr,
  output        io_exe_reqs_2_bits_uop_is_jal,
  output        io_exe_reqs_2_bits_uop_is_sfb,
  output [11:0] io_exe_reqs_2_bits_uop_br_mask,
  output [3:0]  io_exe_reqs_2_bits_uop_br_tag,
  output [4:0]  io_exe_reqs_2_bits_uop_ftq_idx,
  output        io_exe_reqs_2_bits_uop_edge_inst,
  output [5:0]  io_exe_reqs_2_bits_uop_pc_lob,
  output        io_exe_reqs_2_bits_uop_taken,
  output [19:0] io_exe_reqs_2_bits_uop_imm_packed,
  output [11:0] io_exe_reqs_2_bits_uop_csr_addr,
  output [5:0]  io_exe_reqs_2_bits_uop_rob_idx,
  output [4:0]  io_exe_reqs_2_bits_uop_ldq_idx,
  output [4:0]  io_exe_reqs_2_bits_uop_stq_idx,
  output [1:0]  io_exe_reqs_2_bits_uop_rxq_idx,
  output [6:0]  io_exe_reqs_2_bits_uop_pdst,
  output [6:0]  io_exe_reqs_2_bits_uop_prs1,
  output [6:0]  io_exe_reqs_2_bits_uop_prs2,
  output [6:0]  io_exe_reqs_2_bits_uop_prs3,
  output [4:0]  io_exe_reqs_2_bits_uop_ppred,
  output        io_exe_reqs_2_bits_uop_prs1_busy,
  output        io_exe_reqs_2_bits_uop_prs2_busy,
  output        io_exe_reqs_2_bits_uop_prs3_busy,
  output        io_exe_reqs_2_bits_uop_ppred_busy,
  output [6:0]  io_exe_reqs_2_bits_uop_stale_pdst,
  output        io_exe_reqs_2_bits_uop_exception,
  output [63:0] io_exe_reqs_2_bits_uop_exc_cause,
  output        io_exe_reqs_2_bits_uop_bypassable,
  output [4:0]  io_exe_reqs_2_bits_uop_mem_cmd,
  output [1:0]  io_exe_reqs_2_bits_uop_mem_size,
  output        io_exe_reqs_2_bits_uop_mem_signed,
  output        io_exe_reqs_2_bits_uop_is_fence,
  output        io_exe_reqs_2_bits_uop_is_fencei,
  output        io_exe_reqs_2_bits_uop_is_amo,
  output        io_exe_reqs_2_bits_uop_uses_ldq,
  output        io_exe_reqs_2_bits_uop_uses_stq,
  output        io_exe_reqs_2_bits_uop_is_sys_pc2epc,
  output        io_exe_reqs_2_bits_uop_is_unique,
  output        io_exe_reqs_2_bits_uop_flush_on_commit,
  output        io_exe_reqs_2_bits_uop_ldst_is_rs1,
  output [5:0]  io_exe_reqs_2_bits_uop_ldst,
  output [5:0]  io_exe_reqs_2_bits_uop_lrs1,
  output [5:0]  io_exe_reqs_2_bits_uop_lrs2,
  output [5:0]  io_exe_reqs_2_bits_uop_lrs3,
  output        io_exe_reqs_2_bits_uop_ldst_val,
  output [1:0]  io_exe_reqs_2_bits_uop_dst_rtype,
  output [1:0]  io_exe_reqs_2_bits_uop_lrs1_rtype,
  output [1:0]  io_exe_reqs_2_bits_uop_lrs2_rtype,
  output        io_exe_reqs_2_bits_uop_frs3_en,
  output        io_exe_reqs_2_bits_uop_fp_val,
  output        io_exe_reqs_2_bits_uop_fp_single,
  output        io_exe_reqs_2_bits_uop_xcpt_pf_if,
  output        io_exe_reqs_2_bits_uop_xcpt_ae_if,
  output        io_exe_reqs_2_bits_uop_xcpt_ma_if,
  output        io_exe_reqs_2_bits_uop_bp_debug_if,
  output        io_exe_reqs_2_bits_uop_bp_xcpt_if,
  output [1:0]  io_exe_reqs_2_bits_uop_debug_fsrc,
  output [1:0]  io_exe_reqs_2_bits_uop_debug_tsrc,
  output [63:0] io_exe_reqs_2_bits_rs1_data,
  output [63:0] io_exe_reqs_2_bits_rs2_data,
  output [63:0] io_exe_reqs_2_bits_rs3_data,
  output        io_exe_reqs_2_bits_pred_data,
  output [3:0]  io_exe_reqs_2_bits_flagdata,
  output [31:0] io_exe_reqs_2_bits_fflagdata,
  output        io_exe_reqs_2_bits_kill,
  input         io_kill,
  input  [11:0] io_brupdate_b1_resolve_mask,
  input  [11:0] io_brupdate_b1_mispredict_mask,
  input         io_brupdate_b2_uop_switch,
  input         io_brupdate_b2_uop_switch_off,
  input         io_brupdate_b2_uop_is_unicore,
  input  [2:0]  io_brupdate_b2_uop_shift,
  input  [1:0]  io_brupdate_b2_uop_lrs3_rtype,
  input         io_brupdate_b2_uop_rflag,
  input         io_brupdate_b2_uop_wflag,
  input  [3:0]  io_brupdate_b2_uop_prflag,
  input  [3:0]  io_brupdate_b2_uop_pwflag,
  input         io_brupdate_b2_uop_pflag_busy,
  input  [3:0]  io_brupdate_b2_uop_stale_pflag,
  input  [3:0]  io_brupdate_b2_uop_op1_sel,
  input  [3:0]  io_brupdate_b2_uop_op2_sel,
  input  [5:0]  io_brupdate_b2_uop_split_num,
  input  [5:0]  io_brupdate_b2_uop_self_index,
  input  [5:0]  io_brupdate_b2_uop_rob_inst_idx,
  input  [5:0]  io_brupdate_b2_uop_address_num,
  input  [6:0]  io_brupdate_b2_uop_uopc,
  input  [31:0] io_brupdate_b2_uop_inst,
  input  [31:0] io_brupdate_b2_uop_debug_inst,
  input         io_brupdate_b2_uop_is_rvc,
  input  [39:0] io_brupdate_b2_uop_debug_pc,
  input  [2:0]  io_brupdate_b2_uop_iq_type,
  input  [9:0]  io_brupdate_b2_uop_fu_code,
  input  [3:0]  io_brupdate_b2_uop_ctrl_br_type,
  input  [1:0]  io_brupdate_b2_uop_ctrl_op1_sel,
  input  [2:0]  io_brupdate_b2_uop_ctrl_op2_sel,
  input  [2:0]  io_brupdate_b2_uop_ctrl_imm_sel,
  input  [3:0]  io_brupdate_b2_uop_ctrl_op_fcn,
  input         io_brupdate_b2_uop_ctrl_fcn_dw,
  input  [2:0]  io_brupdate_b2_uop_ctrl_csr_cmd,
  input         io_brupdate_b2_uop_ctrl_is_load,
  input         io_brupdate_b2_uop_ctrl_is_sta,
  input         io_brupdate_b2_uop_ctrl_is_std,
  input  [1:0]  io_brupdate_b2_uop_ctrl_op3_sel,
  input  [1:0]  io_brupdate_b2_uop_iw_state,
  input         io_brupdate_b2_uop_iw_p1_poisoned,
  input         io_brupdate_b2_uop_iw_p2_poisoned,
  input         io_brupdate_b2_uop_is_br,
  input         io_brupdate_b2_uop_is_jalr,
  input         io_brupdate_b2_uop_is_jal,
  input         io_brupdate_b2_uop_is_sfb,
  input  [11:0] io_brupdate_b2_uop_br_mask,
  input  [3:0]  io_brupdate_b2_uop_br_tag,
  input  [4:0]  io_brupdate_b2_uop_ftq_idx,
  input         io_brupdate_b2_uop_edge_inst,
  input  [5:0]  io_brupdate_b2_uop_pc_lob,
  input         io_brupdate_b2_uop_taken,
  input  [19:0] io_brupdate_b2_uop_imm_packed,
  input  [11:0] io_brupdate_b2_uop_csr_addr,
  input  [5:0]  io_brupdate_b2_uop_rob_idx,
  input  [4:0]  io_brupdate_b2_uop_ldq_idx,
  input  [4:0]  io_brupdate_b2_uop_stq_idx,
  input  [1:0]  io_brupdate_b2_uop_rxq_idx,
  input  [6:0]  io_brupdate_b2_uop_pdst,
  input  [6:0]  io_brupdate_b2_uop_prs1,
  input  [6:0]  io_brupdate_b2_uop_prs2,
  input  [6:0]  io_brupdate_b2_uop_prs3,
  input  [4:0]  io_brupdate_b2_uop_ppred,
  input         io_brupdate_b2_uop_prs1_busy,
  input         io_brupdate_b2_uop_prs2_busy,
  input         io_brupdate_b2_uop_prs3_busy,
  input         io_brupdate_b2_uop_ppred_busy,
  input  [6:0]  io_brupdate_b2_uop_stale_pdst,
  input         io_brupdate_b2_uop_exception,
  input  [63:0] io_brupdate_b2_uop_exc_cause,
  input         io_brupdate_b2_uop_bypassable,
  input  [4:0]  io_brupdate_b2_uop_mem_cmd,
  input  [1:0]  io_brupdate_b2_uop_mem_size,
  input         io_brupdate_b2_uop_mem_signed,
  input         io_brupdate_b2_uop_is_fence,
  input         io_brupdate_b2_uop_is_fencei,
  input         io_brupdate_b2_uop_is_amo,
  input         io_brupdate_b2_uop_uses_ldq,
  input         io_brupdate_b2_uop_uses_stq,
  input         io_brupdate_b2_uop_is_sys_pc2epc,
  input         io_brupdate_b2_uop_is_unique,
  input         io_brupdate_b2_uop_flush_on_commit,
  input         io_brupdate_b2_uop_ldst_is_rs1,
  input  [5:0]  io_brupdate_b2_uop_ldst,
  input  [5:0]  io_brupdate_b2_uop_lrs1,
  input  [5:0]  io_brupdate_b2_uop_lrs2,
  input  [5:0]  io_brupdate_b2_uop_lrs3,
  input         io_brupdate_b2_uop_ldst_val,
  input  [1:0]  io_brupdate_b2_uop_dst_rtype,
  input  [1:0]  io_brupdate_b2_uop_lrs1_rtype,
  input  [1:0]  io_brupdate_b2_uop_lrs2_rtype,
  input         io_brupdate_b2_uop_frs3_en,
  input         io_brupdate_b2_uop_fp_val,
  input         io_brupdate_b2_uop_fp_single,
  input         io_brupdate_b2_uop_xcpt_pf_if,
  input         io_brupdate_b2_uop_xcpt_ae_if,
  input         io_brupdate_b2_uop_xcpt_ma_if,
  input         io_brupdate_b2_uop_bp_debug_if,
  input         io_brupdate_b2_uop_bp_xcpt_if,
  input  [1:0]  io_brupdate_b2_uop_debug_fsrc,
  input  [1:0]  io_brupdate_b2_uop_debug_tsrc,
  input         io_brupdate_b2_valid,
  input         io_brupdate_b2_mispredict,
  input         io_brupdate_b2_taken,
  input  [2:0]  io_brupdate_b2_cfi_type,
  input  [1:0]  io_brupdate_b2_pc_sel,
  input  [39:0] io_brupdate_b2_jalr_target,
  input  [31:0] io_brupdate_b2_target_offset
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [63:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [63:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [63:0] _RAND_294;
  reg [63:0] _RAND_295;
  reg [63:0] _RAND_296;
  reg [63:0] _RAND_297;
  reg [63:0] _RAND_298;
  reg [63:0] _RAND_299;
  reg [63:0] _RAND_300;
  reg [63:0] _RAND_301;
  reg [63:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [63:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [63:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [63:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [63:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [63:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [63:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
`endif // RANDOMIZE_REG_INIT
  wire  RegisterReadDecode_clock; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_reset; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_valid; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_switch; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_switch_off; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_is_unicore; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_io_iss_uop_shift; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_iss_uop_lrs3_rtype; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_rflag; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_wflag; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_io_iss_uop_prflag; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_io_iss_uop_pwflag; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_pflag_busy; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_io_iss_uop_stale_pflag; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_io_iss_uop_op1_sel; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_io_iss_uop_op2_sel; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_io_iss_uop_split_num; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_io_iss_uop_self_index; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_io_iss_uop_rob_inst_idx; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_io_iss_uop_address_num; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_io_iss_uop_uopc; // @[register-read.scala 86:33]
  wire [31:0] RegisterReadDecode_io_iss_uop_inst; // @[register-read.scala 86:33]
  wire [31:0] RegisterReadDecode_io_iss_uop_debug_inst; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_is_rvc; // @[register-read.scala 86:33]
  wire [39:0] RegisterReadDecode_io_iss_uop_debug_pc; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_io_iss_uop_iq_type; // @[register-read.scala 86:33]
  wire [9:0] RegisterReadDecode_io_iss_uop_fu_code; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_io_iss_uop_ctrl_br_type; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_iss_uop_ctrl_op1_sel; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_io_iss_uop_ctrl_op2_sel; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_io_iss_uop_ctrl_imm_sel; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_io_iss_uop_ctrl_op_fcn; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_ctrl_fcn_dw; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_io_iss_uop_ctrl_csr_cmd; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_ctrl_is_load; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_ctrl_is_sta; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_ctrl_is_std; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_iss_uop_ctrl_op3_sel; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_iss_uop_iw_state; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_iw_p1_poisoned; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_iw_p2_poisoned; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_is_br; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_is_jalr; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_is_jal; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_is_sfb; // @[register-read.scala 86:33]
  wire [11:0] RegisterReadDecode_io_iss_uop_br_mask; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_io_iss_uop_br_tag; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_io_iss_uop_ftq_idx; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_edge_inst; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_io_iss_uop_pc_lob; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_taken; // @[register-read.scala 86:33]
  wire [19:0] RegisterReadDecode_io_iss_uop_imm_packed; // @[register-read.scala 86:33]
  wire [11:0] RegisterReadDecode_io_iss_uop_csr_addr; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_io_iss_uop_rob_idx; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_io_iss_uop_ldq_idx; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_io_iss_uop_stq_idx; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_iss_uop_rxq_idx; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_io_iss_uop_pdst; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_io_iss_uop_prs1; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_io_iss_uop_prs2; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_io_iss_uop_prs3; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_io_iss_uop_ppred; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_prs1_busy; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_prs2_busy; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_prs3_busy; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_ppred_busy; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_io_iss_uop_stale_pdst; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_exception; // @[register-read.scala 86:33]
  wire [63:0] RegisterReadDecode_io_iss_uop_exc_cause; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_bypassable; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_io_iss_uop_mem_cmd; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_iss_uop_mem_size; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_mem_signed; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_is_fence; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_is_fencei; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_is_amo; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_uses_ldq; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_uses_stq; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_is_sys_pc2epc; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_is_unique; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_flush_on_commit; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_ldst_is_rs1; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_io_iss_uop_ldst; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_io_iss_uop_lrs1; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_io_iss_uop_lrs2; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_io_iss_uop_lrs3; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_ldst_val; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_iss_uop_dst_rtype; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_iss_uop_lrs1_rtype; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_iss_uop_lrs2_rtype; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_frs3_en; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_fp_val; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_fp_single; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_xcpt_pf_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_xcpt_ae_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_xcpt_ma_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_bp_debug_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_iss_uop_bp_xcpt_if; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_iss_uop_debug_fsrc; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_iss_uop_debug_tsrc; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_valid; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_switch; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_switch_off; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_is_unicore; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_io_rrd_uop_shift; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_rrd_uop_lrs3_rtype; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_rflag; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_wflag; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_io_rrd_uop_prflag; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_io_rrd_uop_pwflag; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_pflag_busy; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_io_rrd_uop_stale_pflag; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_io_rrd_uop_op1_sel; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_io_rrd_uop_op2_sel; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_io_rrd_uop_split_num; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_io_rrd_uop_self_index; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_io_rrd_uop_rob_inst_idx; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_io_rrd_uop_address_num; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_io_rrd_uop_uopc; // @[register-read.scala 86:33]
  wire [31:0] RegisterReadDecode_io_rrd_uop_inst; // @[register-read.scala 86:33]
  wire [31:0] RegisterReadDecode_io_rrd_uop_debug_inst; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_is_rvc; // @[register-read.scala 86:33]
  wire [39:0] RegisterReadDecode_io_rrd_uop_debug_pc; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_io_rrd_uop_iq_type; // @[register-read.scala 86:33]
  wire [9:0] RegisterReadDecode_io_rrd_uop_fu_code; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_io_rrd_uop_ctrl_br_type; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_rrd_uop_ctrl_op1_sel; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_io_rrd_uop_ctrl_op2_sel; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_io_rrd_uop_ctrl_imm_sel; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_io_rrd_uop_ctrl_op_fcn; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_ctrl_fcn_dw; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_io_rrd_uop_ctrl_csr_cmd; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_ctrl_is_load; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_ctrl_is_sta; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_ctrl_is_std; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_rrd_uop_ctrl_op3_sel; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_rrd_uop_iw_state; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_iw_p1_poisoned; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_iw_p2_poisoned; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_is_br; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_is_jalr; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_is_jal; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_is_sfb; // @[register-read.scala 86:33]
  wire [11:0] RegisterReadDecode_io_rrd_uop_br_mask; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_io_rrd_uop_br_tag; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_io_rrd_uop_ftq_idx; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_edge_inst; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_io_rrd_uop_pc_lob; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_taken; // @[register-read.scala 86:33]
  wire [19:0] RegisterReadDecode_io_rrd_uop_imm_packed; // @[register-read.scala 86:33]
  wire [11:0] RegisterReadDecode_io_rrd_uop_csr_addr; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_io_rrd_uop_rob_idx; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_io_rrd_uop_ldq_idx; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_io_rrd_uop_stq_idx; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_rrd_uop_rxq_idx; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_io_rrd_uop_pdst; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_io_rrd_uop_prs1; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_io_rrd_uop_prs2; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_io_rrd_uop_prs3; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_io_rrd_uop_ppred; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_prs1_busy; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_prs2_busy; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_prs3_busy; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_ppred_busy; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_io_rrd_uop_stale_pdst; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_exception; // @[register-read.scala 86:33]
  wire [63:0] RegisterReadDecode_io_rrd_uop_exc_cause; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_bypassable; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_io_rrd_uop_mem_cmd; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_rrd_uop_mem_size; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_mem_signed; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_is_fence; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_is_fencei; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_is_amo; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_uses_ldq; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_uses_stq; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_is_sys_pc2epc; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_is_unique; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_flush_on_commit; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_ldst_is_rs1; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_io_rrd_uop_ldst; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_io_rrd_uop_lrs1; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_io_rrd_uop_lrs2; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_io_rrd_uop_lrs3; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_ldst_val; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_rrd_uop_dst_rtype; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_rrd_uop_lrs1_rtype; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_rrd_uop_lrs2_rtype; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_frs3_en; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_fp_val; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_fp_single; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_xcpt_pf_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_xcpt_ae_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_xcpt_ma_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_bp_debug_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_io_rrd_uop_bp_xcpt_if; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_rrd_uop_debug_fsrc; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_io_rrd_uop_debug_tsrc; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_clock; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_reset; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_valid; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_switch; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_switch_off; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_is_unicore; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_1_io_iss_uop_shift; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_iss_uop_lrs3_rtype; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_rflag; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_wflag; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_1_io_iss_uop_prflag; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_1_io_iss_uop_pwflag; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_pflag_busy; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_1_io_iss_uop_stale_pflag; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_1_io_iss_uop_op1_sel; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_1_io_iss_uop_op2_sel; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_1_io_iss_uop_split_num; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_1_io_iss_uop_self_index; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_1_io_iss_uop_rob_inst_idx; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_1_io_iss_uop_address_num; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_1_io_iss_uop_uopc; // @[register-read.scala 86:33]
  wire [31:0] RegisterReadDecode_1_io_iss_uop_inst; // @[register-read.scala 86:33]
  wire [31:0] RegisterReadDecode_1_io_iss_uop_debug_inst; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_is_rvc; // @[register-read.scala 86:33]
  wire [39:0] RegisterReadDecode_1_io_iss_uop_debug_pc; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_1_io_iss_uop_iq_type; // @[register-read.scala 86:33]
  wire [9:0] RegisterReadDecode_1_io_iss_uop_fu_code; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_1_io_iss_uop_ctrl_br_type; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_iss_uop_ctrl_op1_sel; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_1_io_iss_uop_ctrl_op2_sel; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_1_io_iss_uop_ctrl_imm_sel; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_1_io_iss_uop_ctrl_op_fcn; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_ctrl_fcn_dw; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_1_io_iss_uop_ctrl_csr_cmd; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_ctrl_is_load; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_ctrl_is_sta; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_ctrl_is_std; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_iss_uop_ctrl_op3_sel; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_iss_uop_iw_state; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_iw_p1_poisoned; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_iw_p2_poisoned; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_is_br; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_is_jalr; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_is_jal; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_is_sfb; // @[register-read.scala 86:33]
  wire [11:0] RegisterReadDecode_1_io_iss_uop_br_mask; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_1_io_iss_uop_br_tag; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_1_io_iss_uop_ftq_idx; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_edge_inst; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_1_io_iss_uop_pc_lob; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_taken; // @[register-read.scala 86:33]
  wire [19:0] RegisterReadDecode_1_io_iss_uop_imm_packed; // @[register-read.scala 86:33]
  wire [11:0] RegisterReadDecode_1_io_iss_uop_csr_addr; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_1_io_iss_uop_rob_idx; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_1_io_iss_uop_ldq_idx; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_1_io_iss_uop_stq_idx; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_iss_uop_rxq_idx; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_1_io_iss_uop_pdst; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_1_io_iss_uop_prs1; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_1_io_iss_uop_prs2; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_1_io_iss_uop_prs3; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_1_io_iss_uop_ppred; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_prs1_busy; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_prs2_busy; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_prs3_busy; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_ppred_busy; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_1_io_iss_uop_stale_pdst; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_exception; // @[register-read.scala 86:33]
  wire [63:0] RegisterReadDecode_1_io_iss_uop_exc_cause; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_bypassable; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_1_io_iss_uop_mem_cmd; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_iss_uop_mem_size; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_mem_signed; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_is_fence; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_is_fencei; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_is_amo; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_uses_ldq; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_uses_stq; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_is_sys_pc2epc; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_is_unique; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_flush_on_commit; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_ldst_is_rs1; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_1_io_iss_uop_ldst; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_1_io_iss_uop_lrs1; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_1_io_iss_uop_lrs2; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_1_io_iss_uop_lrs3; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_ldst_val; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_iss_uop_dst_rtype; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_iss_uop_lrs1_rtype; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_iss_uop_lrs2_rtype; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_frs3_en; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_fp_val; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_fp_single; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_xcpt_pf_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_xcpt_ae_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_xcpt_ma_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_bp_debug_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_iss_uop_bp_xcpt_if; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_iss_uop_debug_fsrc; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_iss_uop_debug_tsrc; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_valid; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_switch; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_switch_off; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_is_unicore; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_1_io_rrd_uop_shift; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_rrd_uop_lrs3_rtype; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_rflag; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_wflag; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_1_io_rrd_uop_prflag; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_1_io_rrd_uop_pwflag; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_pflag_busy; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_1_io_rrd_uop_stale_pflag; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_1_io_rrd_uop_op1_sel; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_1_io_rrd_uop_op2_sel; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_1_io_rrd_uop_split_num; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_1_io_rrd_uop_self_index; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_1_io_rrd_uop_rob_inst_idx; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_1_io_rrd_uop_address_num; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_1_io_rrd_uop_uopc; // @[register-read.scala 86:33]
  wire [31:0] RegisterReadDecode_1_io_rrd_uop_inst; // @[register-read.scala 86:33]
  wire [31:0] RegisterReadDecode_1_io_rrd_uop_debug_inst; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_is_rvc; // @[register-read.scala 86:33]
  wire [39:0] RegisterReadDecode_1_io_rrd_uop_debug_pc; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_1_io_rrd_uop_iq_type; // @[register-read.scala 86:33]
  wire [9:0] RegisterReadDecode_1_io_rrd_uop_fu_code; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_1_io_rrd_uop_ctrl_br_type; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_rrd_uop_ctrl_op1_sel; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_1_io_rrd_uop_ctrl_op2_sel; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_1_io_rrd_uop_ctrl_imm_sel; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_1_io_rrd_uop_ctrl_op_fcn; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_ctrl_fcn_dw; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_1_io_rrd_uop_ctrl_csr_cmd; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_ctrl_is_load; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_ctrl_is_sta; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_ctrl_is_std; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_rrd_uop_ctrl_op3_sel; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_rrd_uop_iw_state; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_iw_p1_poisoned; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_iw_p2_poisoned; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_is_br; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_is_jalr; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_is_jal; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_is_sfb; // @[register-read.scala 86:33]
  wire [11:0] RegisterReadDecode_1_io_rrd_uop_br_mask; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_1_io_rrd_uop_br_tag; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_1_io_rrd_uop_ftq_idx; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_edge_inst; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_1_io_rrd_uop_pc_lob; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_taken; // @[register-read.scala 86:33]
  wire [19:0] RegisterReadDecode_1_io_rrd_uop_imm_packed; // @[register-read.scala 86:33]
  wire [11:0] RegisterReadDecode_1_io_rrd_uop_csr_addr; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_1_io_rrd_uop_rob_idx; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_1_io_rrd_uop_ldq_idx; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_1_io_rrd_uop_stq_idx; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_rrd_uop_rxq_idx; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_1_io_rrd_uop_pdst; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_1_io_rrd_uop_prs1; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_1_io_rrd_uop_prs2; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_1_io_rrd_uop_prs3; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_1_io_rrd_uop_ppred; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_prs1_busy; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_prs2_busy; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_prs3_busy; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_ppred_busy; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_1_io_rrd_uop_stale_pdst; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_exception; // @[register-read.scala 86:33]
  wire [63:0] RegisterReadDecode_1_io_rrd_uop_exc_cause; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_bypassable; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_1_io_rrd_uop_mem_cmd; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_rrd_uop_mem_size; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_mem_signed; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_is_fence; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_is_fencei; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_is_amo; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_uses_ldq; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_uses_stq; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_is_sys_pc2epc; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_is_unique; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_flush_on_commit; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_ldst_is_rs1; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_1_io_rrd_uop_ldst; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_1_io_rrd_uop_lrs1; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_1_io_rrd_uop_lrs2; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_1_io_rrd_uop_lrs3; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_ldst_val; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_rrd_uop_dst_rtype; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_rrd_uop_lrs1_rtype; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_rrd_uop_lrs2_rtype; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_frs3_en; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_fp_val; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_fp_single; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_xcpt_pf_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_xcpt_ae_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_xcpt_ma_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_bp_debug_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_1_io_rrd_uop_bp_xcpt_if; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_rrd_uop_debug_fsrc; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_1_io_rrd_uop_debug_tsrc; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_clock; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_reset; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_valid; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_switch; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_switch_off; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_is_unicore; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_2_io_iss_uop_shift; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_iss_uop_lrs3_rtype; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_rflag; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_wflag; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_2_io_iss_uop_prflag; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_2_io_iss_uop_pwflag; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_pflag_busy; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_2_io_iss_uop_stale_pflag; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_2_io_iss_uop_op1_sel; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_2_io_iss_uop_op2_sel; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_2_io_iss_uop_split_num; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_2_io_iss_uop_self_index; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_2_io_iss_uop_rob_inst_idx; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_2_io_iss_uop_address_num; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_2_io_iss_uop_uopc; // @[register-read.scala 86:33]
  wire [31:0] RegisterReadDecode_2_io_iss_uop_inst; // @[register-read.scala 86:33]
  wire [31:0] RegisterReadDecode_2_io_iss_uop_debug_inst; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_is_rvc; // @[register-read.scala 86:33]
  wire [39:0] RegisterReadDecode_2_io_iss_uop_debug_pc; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_2_io_iss_uop_iq_type; // @[register-read.scala 86:33]
  wire [9:0] RegisterReadDecode_2_io_iss_uop_fu_code; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_2_io_iss_uop_ctrl_br_type; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_iss_uop_ctrl_op1_sel; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_2_io_iss_uop_ctrl_op2_sel; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_2_io_iss_uop_ctrl_imm_sel; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_2_io_iss_uop_ctrl_op_fcn; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_ctrl_fcn_dw; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_2_io_iss_uop_ctrl_csr_cmd; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_ctrl_is_load; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_ctrl_is_sta; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_ctrl_is_std; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_iss_uop_ctrl_op3_sel; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_iss_uop_iw_state; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_iw_p1_poisoned; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_iw_p2_poisoned; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_is_br; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_is_jalr; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_is_jal; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_is_sfb; // @[register-read.scala 86:33]
  wire [11:0] RegisterReadDecode_2_io_iss_uop_br_mask; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_2_io_iss_uop_br_tag; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_2_io_iss_uop_ftq_idx; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_edge_inst; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_2_io_iss_uop_pc_lob; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_taken; // @[register-read.scala 86:33]
  wire [19:0] RegisterReadDecode_2_io_iss_uop_imm_packed; // @[register-read.scala 86:33]
  wire [11:0] RegisterReadDecode_2_io_iss_uop_csr_addr; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_2_io_iss_uop_rob_idx; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_2_io_iss_uop_ldq_idx; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_2_io_iss_uop_stq_idx; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_iss_uop_rxq_idx; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_2_io_iss_uop_pdst; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_2_io_iss_uop_prs1; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_2_io_iss_uop_prs2; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_2_io_iss_uop_prs3; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_2_io_iss_uop_ppred; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_prs1_busy; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_prs2_busy; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_prs3_busy; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_ppred_busy; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_2_io_iss_uop_stale_pdst; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_exception; // @[register-read.scala 86:33]
  wire [63:0] RegisterReadDecode_2_io_iss_uop_exc_cause; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_bypassable; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_2_io_iss_uop_mem_cmd; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_iss_uop_mem_size; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_mem_signed; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_is_fence; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_is_fencei; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_is_amo; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_uses_ldq; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_uses_stq; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_is_sys_pc2epc; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_is_unique; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_flush_on_commit; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_ldst_is_rs1; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_2_io_iss_uop_ldst; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_2_io_iss_uop_lrs1; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_2_io_iss_uop_lrs2; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_2_io_iss_uop_lrs3; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_ldst_val; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_iss_uop_dst_rtype; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_iss_uop_lrs1_rtype; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_iss_uop_lrs2_rtype; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_frs3_en; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_fp_val; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_fp_single; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_xcpt_pf_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_xcpt_ae_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_xcpt_ma_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_bp_debug_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_iss_uop_bp_xcpt_if; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_iss_uop_debug_fsrc; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_iss_uop_debug_tsrc; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_valid; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_switch; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_switch_off; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_is_unicore; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_2_io_rrd_uop_shift; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_rrd_uop_lrs3_rtype; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_rflag; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_wflag; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_2_io_rrd_uop_prflag; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_2_io_rrd_uop_pwflag; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_pflag_busy; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_2_io_rrd_uop_stale_pflag; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_2_io_rrd_uop_op1_sel; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_2_io_rrd_uop_op2_sel; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_2_io_rrd_uop_split_num; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_2_io_rrd_uop_self_index; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_2_io_rrd_uop_rob_inst_idx; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_2_io_rrd_uop_address_num; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_2_io_rrd_uop_uopc; // @[register-read.scala 86:33]
  wire [31:0] RegisterReadDecode_2_io_rrd_uop_inst; // @[register-read.scala 86:33]
  wire [31:0] RegisterReadDecode_2_io_rrd_uop_debug_inst; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_is_rvc; // @[register-read.scala 86:33]
  wire [39:0] RegisterReadDecode_2_io_rrd_uop_debug_pc; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_2_io_rrd_uop_iq_type; // @[register-read.scala 86:33]
  wire [9:0] RegisterReadDecode_2_io_rrd_uop_fu_code; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_2_io_rrd_uop_ctrl_br_type; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_rrd_uop_ctrl_op1_sel; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_2_io_rrd_uop_ctrl_op2_sel; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_2_io_rrd_uop_ctrl_imm_sel; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_2_io_rrd_uop_ctrl_op_fcn; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_ctrl_fcn_dw; // @[register-read.scala 86:33]
  wire [2:0] RegisterReadDecode_2_io_rrd_uop_ctrl_csr_cmd; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_ctrl_is_load; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_ctrl_is_sta; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_ctrl_is_std; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_rrd_uop_ctrl_op3_sel; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_rrd_uop_iw_state; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_iw_p1_poisoned; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_iw_p2_poisoned; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_is_br; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_is_jalr; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_is_jal; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_is_sfb; // @[register-read.scala 86:33]
  wire [11:0] RegisterReadDecode_2_io_rrd_uop_br_mask; // @[register-read.scala 86:33]
  wire [3:0] RegisterReadDecode_2_io_rrd_uop_br_tag; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_2_io_rrd_uop_ftq_idx; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_edge_inst; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_2_io_rrd_uop_pc_lob; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_taken; // @[register-read.scala 86:33]
  wire [19:0] RegisterReadDecode_2_io_rrd_uop_imm_packed; // @[register-read.scala 86:33]
  wire [11:0] RegisterReadDecode_2_io_rrd_uop_csr_addr; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_2_io_rrd_uop_rob_idx; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_2_io_rrd_uop_ldq_idx; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_2_io_rrd_uop_stq_idx; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_rrd_uop_rxq_idx; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_2_io_rrd_uop_pdst; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_2_io_rrd_uop_prs1; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_2_io_rrd_uop_prs2; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_2_io_rrd_uop_prs3; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_2_io_rrd_uop_ppred; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_prs1_busy; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_prs2_busy; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_prs3_busy; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_ppred_busy; // @[register-read.scala 86:33]
  wire [6:0] RegisterReadDecode_2_io_rrd_uop_stale_pdst; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_exception; // @[register-read.scala 86:33]
  wire [63:0] RegisterReadDecode_2_io_rrd_uop_exc_cause; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_bypassable; // @[register-read.scala 86:33]
  wire [4:0] RegisterReadDecode_2_io_rrd_uop_mem_cmd; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_rrd_uop_mem_size; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_mem_signed; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_is_fence; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_is_fencei; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_is_amo; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_uses_ldq; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_uses_stq; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_is_sys_pc2epc; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_is_unique; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_flush_on_commit; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_ldst_is_rs1; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_2_io_rrd_uop_ldst; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_2_io_rrd_uop_lrs1; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_2_io_rrd_uop_lrs2; // @[register-read.scala 86:33]
  wire [5:0] RegisterReadDecode_2_io_rrd_uop_lrs3; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_ldst_val; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_rrd_uop_dst_rtype; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_rrd_uop_lrs1_rtype; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_rrd_uop_lrs2_rtype; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_frs3_en; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_fp_val; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_fp_single; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_xcpt_pf_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_xcpt_ae_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_xcpt_ma_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_bp_debug_if; // @[register-read.scala 86:33]
  wire  RegisterReadDecode_2_io_rrd_uop_bp_xcpt_if; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_rrd_uop_debug_fsrc; // @[register-read.scala 86:33]
  wire [1:0] RegisterReadDecode_2_io_rrd_uop_debug_tsrc; // @[register-read.scala 86:33]
  reg  exe_reg_valids_0; // @[register-read.scala 72:33]
  reg  exe_reg_valids_1; // @[register-read.scala 72:33]
  reg  exe_reg_valids_2; // @[register-read.scala 72:33]
  reg  exe_reg_uops_0_switch; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_switch_off; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_is_unicore; // @[register-read.scala 73:29]
  reg [2:0] exe_reg_uops_0_shift; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_0_lrs3_rtype; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_rflag; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_wflag; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_0_prflag; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_0_pwflag; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_pflag_busy; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_0_stale_pflag; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_0_op1_sel; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_0_op2_sel; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_0_split_num; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_0_self_index; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_0_rob_inst_idx; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_0_address_num; // @[register-read.scala 73:29]
  reg [6:0] exe_reg_uops_0_uopc; // @[register-read.scala 73:29]
  reg [31:0] exe_reg_uops_0_inst; // @[register-read.scala 73:29]
  reg [31:0] exe_reg_uops_0_debug_inst; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_is_rvc; // @[register-read.scala 73:29]
  reg [39:0] exe_reg_uops_0_debug_pc; // @[register-read.scala 73:29]
  reg [2:0] exe_reg_uops_0_iq_type; // @[register-read.scala 73:29]
  reg [9:0] exe_reg_uops_0_fu_code; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_0_ctrl_br_type; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_0_ctrl_op1_sel; // @[register-read.scala 73:29]
  reg [2:0] exe_reg_uops_0_ctrl_op2_sel; // @[register-read.scala 73:29]
  reg [2:0] exe_reg_uops_0_ctrl_imm_sel; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_0_ctrl_op_fcn; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_ctrl_fcn_dw; // @[register-read.scala 73:29]
  reg [2:0] exe_reg_uops_0_ctrl_csr_cmd; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_ctrl_is_load; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_ctrl_is_sta; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_ctrl_is_std; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_0_ctrl_op3_sel; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_0_iw_state; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_iw_p1_poisoned; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_iw_p2_poisoned; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_is_br; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_is_jalr; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_is_jal; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_is_sfb; // @[register-read.scala 73:29]
  reg [11:0] exe_reg_uops_0_br_mask; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_0_br_tag; // @[register-read.scala 73:29]
  reg [4:0] exe_reg_uops_0_ftq_idx; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_edge_inst; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_0_pc_lob; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_taken; // @[register-read.scala 73:29]
  reg [19:0] exe_reg_uops_0_imm_packed; // @[register-read.scala 73:29]
  reg [11:0] exe_reg_uops_0_csr_addr; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_0_rob_idx; // @[register-read.scala 73:29]
  reg [4:0] exe_reg_uops_0_ldq_idx; // @[register-read.scala 73:29]
  reg [4:0] exe_reg_uops_0_stq_idx; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_0_rxq_idx; // @[register-read.scala 73:29]
  reg [6:0] exe_reg_uops_0_pdst; // @[register-read.scala 73:29]
  reg [6:0] exe_reg_uops_0_prs1; // @[register-read.scala 73:29]
  reg [6:0] exe_reg_uops_0_prs2; // @[register-read.scala 73:29]
  reg [6:0] exe_reg_uops_0_prs3; // @[register-read.scala 73:29]
  reg [4:0] exe_reg_uops_0_ppred; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_prs1_busy; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_prs2_busy; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_prs3_busy; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_ppred_busy; // @[register-read.scala 73:29]
  reg [6:0] exe_reg_uops_0_stale_pdst; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_exception; // @[register-read.scala 73:29]
  reg [63:0] exe_reg_uops_0_exc_cause; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_bypassable; // @[register-read.scala 73:29]
  reg [4:0] exe_reg_uops_0_mem_cmd; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_0_mem_size; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_mem_signed; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_is_fence; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_is_fencei; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_is_amo; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_uses_ldq; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_uses_stq; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_is_sys_pc2epc; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_is_unique; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_flush_on_commit; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_ldst_is_rs1; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_0_ldst; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_0_lrs1; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_0_lrs2; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_0_lrs3; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_ldst_val; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_0_dst_rtype; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_0_lrs1_rtype; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_0_lrs2_rtype; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_frs3_en; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_fp_val; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_fp_single; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_xcpt_pf_if; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_xcpt_ae_if; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_xcpt_ma_if; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_bp_debug_if; // @[register-read.scala 73:29]
  reg  exe_reg_uops_0_bp_xcpt_if; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_0_debug_fsrc; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_0_debug_tsrc; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_switch; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_switch_off; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_is_unicore; // @[register-read.scala 73:29]
  reg [2:0] exe_reg_uops_1_shift; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_1_lrs3_rtype; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_rflag; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_wflag; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_1_prflag; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_1_pwflag; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_pflag_busy; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_1_stale_pflag; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_1_op1_sel; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_1_op2_sel; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_1_split_num; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_1_self_index; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_1_rob_inst_idx; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_1_address_num; // @[register-read.scala 73:29]
  reg [6:0] exe_reg_uops_1_uopc; // @[register-read.scala 73:29]
  reg [31:0] exe_reg_uops_1_inst; // @[register-read.scala 73:29]
  reg [31:0] exe_reg_uops_1_debug_inst; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_is_rvc; // @[register-read.scala 73:29]
  reg [39:0] exe_reg_uops_1_debug_pc; // @[register-read.scala 73:29]
  reg [2:0] exe_reg_uops_1_iq_type; // @[register-read.scala 73:29]
  reg [9:0] exe_reg_uops_1_fu_code; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_1_ctrl_br_type; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_1_ctrl_op1_sel; // @[register-read.scala 73:29]
  reg [2:0] exe_reg_uops_1_ctrl_op2_sel; // @[register-read.scala 73:29]
  reg [2:0] exe_reg_uops_1_ctrl_imm_sel; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_1_ctrl_op_fcn; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_ctrl_fcn_dw; // @[register-read.scala 73:29]
  reg [2:0] exe_reg_uops_1_ctrl_csr_cmd; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_ctrl_is_load; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_ctrl_is_sta; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_ctrl_is_std; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_1_ctrl_op3_sel; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_1_iw_state; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_iw_p1_poisoned; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_iw_p2_poisoned; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_is_br; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_is_jalr; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_is_jal; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_is_sfb; // @[register-read.scala 73:29]
  reg [11:0] exe_reg_uops_1_br_mask; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_1_br_tag; // @[register-read.scala 73:29]
  reg [4:0] exe_reg_uops_1_ftq_idx; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_edge_inst; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_1_pc_lob; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_taken; // @[register-read.scala 73:29]
  reg [19:0] exe_reg_uops_1_imm_packed; // @[register-read.scala 73:29]
  reg [11:0] exe_reg_uops_1_csr_addr; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_1_rob_idx; // @[register-read.scala 73:29]
  reg [4:0] exe_reg_uops_1_ldq_idx; // @[register-read.scala 73:29]
  reg [4:0] exe_reg_uops_1_stq_idx; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_1_rxq_idx; // @[register-read.scala 73:29]
  reg [6:0] exe_reg_uops_1_pdst; // @[register-read.scala 73:29]
  reg [6:0] exe_reg_uops_1_prs1; // @[register-read.scala 73:29]
  reg [6:0] exe_reg_uops_1_prs2; // @[register-read.scala 73:29]
  reg [6:0] exe_reg_uops_1_prs3; // @[register-read.scala 73:29]
  reg [4:0] exe_reg_uops_1_ppred; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_prs1_busy; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_prs2_busy; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_prs3_busy; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_ppred_busy; // @[register-read.scala 73:29]
  reg [6:0] exe_reg_uops_1_stale_pdst; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_exception; // @[register-read.scala 73:29]
  reg [63:0] exe_reg_uops_1_exc_cause; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_bypassable; // @[register-read.scala 73:29]
  reg [4:0] exe_reg_uops_1_mem_cmd; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_1_mem_size; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_mem_signed; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_is_fence; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_is_fencei; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_is_amo; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_uses_ldq; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_uses_stq; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_is_sys_pc2epc; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_is_unique; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_flush_on_commit; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_ldst_is_rs1; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_1_ldst; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_1_lrs1; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_1_lrs2; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_1_lrs3; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_ldst_val; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_1_dst_rtype; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_1_lrs1_rtype; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_1_lrs2_rtype; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_frs3_en; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_fp_val; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_fp_single; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_xcpt_pf_if; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_xcpt_ae_if; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_xcpt_ma_if; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_bp_debug_if; // @[register-read.scala 73:29]
  reg  exe_reg_uops_1_bp_xcpt_if; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_1_debug_fsrc; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_1_debug_tsrc; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_switch; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_switch_off; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_is_unicore; // @[register-read.scala 73:29]
  reg [2:0] exe_reg_uops_2_shift; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_2_lrs3_rtype; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_rflag; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_wflag; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_2_prflag; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_2_pwflag; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_pflag_busy; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_2_stale_pflag; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_2_op1_sel; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_2_op2_sel; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_2_split_num; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_2_self_index; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_2_rob_inst_idx; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_2_address_num; // @[register-read.scala 73:29]
  reg [6:0] exe_reg_uops_2_uopc; // @[register-read.scala 73:29]
  reg [31:0] exe_reg_uops_2_inst; // @[register-read.scala 73:29]
  reg [31:0] exe_reg_uops_2_debug_inst; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_is_rvc; // @[register-read.scala 73:29]
  reg [39:0] exe_reg_uops_2_debug_pc; // @[register-read.scala 73:29]
  reg [2:0] exe_reg_uops_2_iq_type; // @[register-read.scala 73:29]
  reg [9:0] exe_reg_uops_2_fu_code; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_2_ctrl_br_type; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_2_ctrl_op1_sel; // @[register-read.scala 73:29]
  reg [2:0] exe_reg_uops_2_ctrl_op2_sel; // @[register-read.scala 73:29]
  reg [2:0] exe_reg_uops_2_ctrl_imm_sel; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_2_ctrl_op_fcn; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_ctrl_fcn_dw; // @[register-read.scala 73:29]
  reg [2:0] exe_reg_uops_2_ctrl_csr_cmd; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_ctrl_is_load; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_ctrl_is_sta; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_ctrl_is_std; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_2_ctrl_op3_sel; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_2_iw_state; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_iw_p1_poisoned; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_iw_p2_poisoned; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_is_br; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_is_jalr; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_is_jal; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_is_sfb; // @[register-read.scala 73:29]
  reg [11:0] exe_reg_uops_2_br_mask; // @[register-read.scala 73:29]
  reg [3:0] exe_reg_uops_2_br_tag; // @[register-read.scala 73:29]
  reg [4:0] exe_reg_uops_2_ftq_idx; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_edge_inst; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_2_pc_lob; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_taken; // @[register-read.scala 73:29]
  reg [19:0] exe_reg_uops_2_imm_packed; // @[register-read.scala 73:29]
  reg [11:0] exe_reg_uops_2_csr_addr; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_2_rob_idx; // @[register-read.scala 73:29]
  reg [4:0] exe_reg_uops_2_ldq_idx; // @[register-read.scala 73:29]
  reg [4:0] exe_reg_uops_2_stq_idx; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_2_rxq_idx; // @[register-read.scala 73:29]
  reg [6:0] exe_reg_uops_2_pdst; // @[register-read.scala 73:29]
  reg [6:0] exe_reg_uops_2_prs1; // @[register-read.scala 73:29]
  reg [6:0] exe_reg_uops_2_prs2; // @[register-read.scala 73:29]
  reg [6:0] exe_reg_uops_2_prs3; // @[register-read.scala 73:29]
  reg [4:0] exe_reg_uops_2_ppred; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_prs1_busy; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_prs2_busy; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_prs3_busy; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_ppred_busy; // @[register-read.scala 73:29]
  reg [6:0] exe_reg_uops_2_stale_pdst; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_exception; // @[register-read.scala 73:29]
  reg [63:0] exe_reg_uops_2_exc_cause; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_bypassable; // @[register-read.scala 73:29]
  reg [4:0] exe_reg_uops_2_mem_cmd; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_2_mem_size; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_mem_signed; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_is_fence; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_is_fencei; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_is_amo; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_uses_ldq; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_uses_stq; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_is_sys_pc2epc; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_is_unique; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_flush_on_commit; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_ldst_is_rs1; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_2_ldst; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_2_lrs1; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_2_lrs2; // @[register-read.scala 73:29]
  reg [5:0] exe_reg_uops_2_lrs3; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_ldst_val; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_2_dst_rtype; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_2_lrs1_rtype; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_2_lrs2_rtype; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_frs3_en; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_fp_val; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_fp_single; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_xcpt_pf_if; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_xcpt_ae_if; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_xcpt_ma_if; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_bp_debug_if; // @[register-read.scala 73:29]
  reg  exe_reg_uops_2_bp_xcpt_if; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_2_debug_fsrc; // @[register-read.scala 73:29]
  reg [1:0] exe_reg_uops_2_debug_tsrc; // @[register-read.scala 73:29]
  reg [63:0] exe_reg_rs1_data_0; // @[register-read.scala 74:29]
  reg [63:0] exe_reg_rs1_data_1; // @[register-read.scala 74:29]
  reg [63:0] exe_reg_rs1_data_2; // @[register-read.scala 74:29]
  reg [63:0] exe_reg_rs2_data_0; // @[register-read.scala 75:29]
  reg [63:0] exe_reg_rs2_data_1; // @[register-read.scala 75:29]
  reg [63:0] exe_reg_rs2_data_2; // @[register-read.scala 75:29]
  reg [63:0] exe_reg_rs3_data_0; // @[register-read.scala 76:29]
  reg [63:0] exe_reg_rs3_data_1; // @[register-read.scala 76:29]
  reg [63:0] exe_reg_rs3_data_2; // @[register-read.scala 76:29]
  reg [3:0] exe_reg_flag_data_0; // @[register-read.scala 79:30]
  reg [3:0] exe_reg_flag_data_1; // @[register-read.scala 79:30]
  reg [3:0] exe_reg_flag_data_2; // @[register-read.scala 79:30]
  wire [11:0] _T = io_brupdate_b1_mispredict_mask & RegisterReadDecode_io_rrd_uop_br_mask; // @[util.scala 175:51]
  wire  _T_1 = _T != 12'h0; // @[util.scala 175:59]
  wire  _T_2 = ~_T_1; // @[register-read.scala 91:17]
  reg  REG; // @[register-read.scala 90:29]
  wire [11:0] _T_4 = ~io_brupdate_b1_resolve_mask; // @[util.scala 131:37]
  reg  REG_1_switch; // @[register-read.scala 92:29]
  reg  REG_1_switch_off; // @[register-read.scala 92:29]
  reg  REG_1_is_unicore; // @[register-read.scala 92:29]
  reg [2:0] REG_1_shift; // @[register-read.scala 92:29]
  reg [1:0] REG_1_lrs3_rtype; // @[register-read.scala 92:29]
  reg  REG_1_rflag; // @[register-read.scala 92:29]
  reg  REG_1_wflag; // @[register-read.scala 92:29]
  reg [3:0] REG_1_prflag; // @[register-read.scala 92:29]
  reg [3:0] REG_1_pwflag; // @[register-read.scala 92:29]
  reg  REG_1_pflag_busy; // @[register-read.scala 92:29]
  reg [3:0] REG_1_stale_pflag; // @[register-read.scala 92:29]
  reg [3:0] REG_1_op1_sel; // @[register-read.scala 92:29]
  reg [3:0] REG_1_op2_sel; // @[register-read.scala 92:29]
  reg [5:0] REG_1_split_num; // @[register-read.scala 92:29]
  reg [5:0] REG_1_self_index; // @[register-read.scala 92:29]
  reg [5:0] REG_1_rob_inst_idx; // @[register-read.scala 92:29]
  reg [5:0] REG_1_address_num; // @[register-read.scala 92:29]
  reg [6:0] REG_1_uopc; // @[register-read.scala 92:29]
  reg [31:0] REG_1_inst; // @[register-read.scala 92:29]
  reg [31:0] REG_1_debug_inst; // @[register-read.scala 92:29]
  reg  REG_1_is_rvc; // @[register-read.scala 92:29]
  reg [39:0] REG_1_debug_pc; // @[register-read.scala 92:29]
  reg [2:0] REG_1_iq_type; // @[register-read.scala 92:29]
  reg [9:0] REG_1_fu_code; // @[register-read.scala 92:29]
  reg [3:0] REG_1_ctrl_br_type; // @[register-read.scala 92:29]
  reg [1:0] REG_1_ctrl_op1_sel; // @[register-read.scala 92:29]
  reg [2:0] REG_1_ctrl_op2_sel; // @[register-read.scala 92:29]
  reg [2:0] REG_1_ctrl_imm_sel; // @[register-read.scala 92:29]
  reg [3:0] REG_1_ctrl_op_fcn; // @[register-read.scala 92:29]
  reg  REG_1_ctrl_fcn_dw; // @[register-read.scala 92:29]
  reg [2:0] REG_1_ctrl_csr_cmd; // @[register-read.scala 92:29]
  reg  REG_1_ctrl_is_load; // @[register-read.scala 92:29]
  reg  REG_1_ctrl_is_sta; // @[register-read.scala 92:29]
  reg  REG_1_ctrl_is_std; // @[register-read.scala 92:29]
  reg [1:0] REG_1_ctrl_op3_sel; // @[register-read.scala 92:29]
  reg [1:0] REG_1_iw_state; // @[register-read.scala 92:29]
  reg  REG_1_iw_p1_poisoned; // @[register-read.scala 92:29]
  reg  REG_1_iw_p2_poisoned; // @[register-read.scala 92:29]
  reg  REG_1_is_br; // @[register-read.scala 92:29]
  reg  REG_1_is_jalr; // @[register-read.scala 92:29]
  reg  REG_1_is_jal; // @[register-read.scala 92:29]
  reg  REG_1_is_sfb; // @[register-read.scala 92:29]
  reg [11:0] REG_1_br_mask; // @[register-read.scala 92:29]
  reg [3:0] REG_1_br_tag; // @[register-read.scala 92:29]
  reg [4:0] REG_1_ftq_idx; // @[register-read.scala 92:29]
  reg  REG_1_edge_inst; // @[register-read.scala 92:29]
  reg [5:0] REG_1_pc_lob; // @[register-read.scala 92:29]
  reg  REG_1_taken; // @[register-read.scala 92:29]
  reg [19:0] REG_1_imm_packed; // @[register-read.scala 92:29]
  reg [11:0] REG_1_csr_addr; // @[register-read.scala 92:29]
  reg [5:0] REG_1_rob_idx; // @[register-read.scala 92:29]
  reg [4:0] REG_1_ldq_idx; // @[register-read.scala 92:29]
  reg [4:0] REG_1_stq_idx; // @[register-read.scala 92:29]
  reg [1:0] REG_1_rxq_idx; // @[register-read.scala 92:29]
  reg [6:0] REG_1_pdst; // @[register-read.scala 92:29]
  reg [6:0] REG_1_prs1; // @[register-read.scala 92:29]
  reg [6:0] REG_1_prs2; // @[register-read.scala 92:29]
  reg [6:0] REG_1_prs3; // @[register-read.scala 92:29]
  reg [4:0] REG_1_ppred; // @[register-read.scala 92:29]
  reg  REG_1_prs1_busy; // @[register-read.scala 92:29]
  reg  REG_1_prs2_busy; // @[register-read.scala 92:29]
  reg  REG_1_prs3_busy; // @[register-read.scala 92:29]
  reg  REG_1_ppred_busy; // @[register-read.scala 92:29]
  reg [6:0] REG_1_stale_pdst; // @[register-read.scala 92:29]
  reg  REG_1_exception; // @[register-read.scala 92:29]
  reg [63:0] REG_1_exc_cause; // @[register-read.scala 92:29]
  reg  REG_1_bypassable; // @[register-read.scala 92:29]
  reg [4:0] REG_1_mem_cmd; // @[register-read.scala 92:29]
  reg [1:0] REG_1_mem_size; // @[register-read.scala 92:29]
  reg  REG_1_mem_signed; // @[register-read.scala 92:29]
  reg  REG_1_is_fence; // @[register-read.scala 92:29]
  reg  REG_1_is_fencei; // @[register-read.scala 92:29]
  reg  REG_1_is_amo; // @[register-read.scala 92:29]
  reg  REG_1_uses_ldq; // @[register-read.scala 92:29]
  reg  REG_1_uses_stq; // @[register-read.scala 92:29]
  reg  REG_1_is_sys_pc2epc; // @[register-read.scala 92:29]
  reg  REG_1_is_unique; // @[register-read.scala 92:29]
  reg  REG_1_flush_on_commit; // @[register-read.scala 92:29]
  reg  REG_1_ldst_is_rs1; // @[register-read.scala 92:29]
  reg [5:0] REG_1_ldst; // @[register-read.scala 92:29]
  reg [5:0] REG_1_lrs1; // @[register-read.scala 92:29]
  reg [5:0] REG_1_lrs2; // @[register-read.scala 92:29]
  reg [5:0] REG_1_lrs3; // @[register-read.scala 92:29]
  reg  REG_1_ldst_val; // @[register-read.scala 92:29]
  reg [1:0] REG_1_dst_rtype; // @[register-read.scala 92:29]
  reg [1:0] REG_1_lrs1_rtype; // @[register-read.scala 92:29]
  reg [1:0] REG_1_lrs2_rtype; // @[register-read.scala 92:29]
  reg  REG_1_frs3_en; // @[register-read.scala 92:29]
  reg  REG_1_fp_val; // @[register-read.scala 92:29]
  reg  REG_1_fp_single; // @[register-read.scala 92:29]
  reg  REG_1_xcpt_pf_if; // @[register-read.scala 92:29]
  reg  REG_1_xcpt_ae_if; // @[register-read.scala 92:29]
  reg  REG_1_xcpt_ma_if; // @[register-read.scala 92:29]
  reg  REG_1_bp_debug_if; // @[register-read.scala 92:29]
  reg  REG_1_bp_xcpt_if; // @[register-read.scala 92:29]
  reg [1:0] REG_1_debug_fsrc; // @[register-read.scala 92:29]
  reg [1:0] REG_1_debug_tsrc; // @[register-read.scala 92:29]
  wire [11:0] _T_6 = io_brupdate_b1_mispredict_mask & RegisterReadDecode_1_io_rrd_uop_br_mask; // @[util.scala 175:51]
  wire  _T_7 = _T_6 != 12'h0; // @[util.scala 175:59]
  wire  _T_8 = ~_T_7; // @[register-read.scala 91:17]
  reg  REG_2; // @[register-read.scala 90:29]
  reg  REG_3_switch; // @[register-read.scala 92:29]
  reg  REG_3_switch_off; // @[register-read.scala 92:29]
  reg  REG_3_is_unicore; // @[register-read.scala 92:29]
  reg [2:0] REG_3_shift; // @[register-read.scala 92:29]
  reg [1:0] REG_3_lrs3_rtype; // @[register-read.scala 92:29]
  reg  REG_3_rflag; // @[register-read.scala 92:29]
  reg  REG_3_wflag; // @[register-read.scala 92:29]
  reg [3:0] REG_3_prflag; // @[register-read.scala 92:29]
  reg [3:0] REG_3_pwflag; // @[register-read.scala 92:29]
  reg  REG_3_pflag_busy; // @[register-read.scala 92:29]
  reg [3:0] REG_3_stale_pflag; // @[register-read.scala 92:29]
  reg [3:0] REG_3_op1_sel; // @[register-read.scala 92:29]
  reg [3:0] REG_3_op2_sel; // @[register-read.scala 92:29]
  reg [5:0] REG_3_split_num; // @[register-read.scala 92:29]
  reg [5:0] REG_3_self_index; // @[register-read.scala 92:29]
  reg [5:0] REG_3_rob_inst_idx; // @[register-read.scala 92:29]
  reg [5:0] REG_3_address_num; // @[register-read.scala 92:29]
  reg [6:0] REG_3_uopc; // @[register-read.scala 92:29]
  reg [31:0] REG_3_inst; // @[register-read.scala 92:29]
  reg [31:0] REG_3_debug_inst; // @[register-read.scala 92:29]
  reg  REG_3_is_rvc; // @[register-read.scala 92:29]
  reg [39:0] REG_3_debug_pc; // @[register-read.scala 92:29]
  reg [2:0] REG_3_iq_type; // @[register-read.scala 92:29]
  reg [9:0] REG_3_fu_code; // @[register-read.scala 92:29]
  reg [3:0] REG_3_ctrl_br_type; // @[register-read.scala 92:29]
  reg [1:0] REG_3_ctrl_op1_sel; // @[register-read.scala 92:29]
  reg [2:0] REG_3_ctrl_op2_sel; // @[register-read.scala 92:29]
  reg [2:0] REG_3_ctrl_imm_sel; // @[register-read.scala 92:29]
  reg [3:0] REG_3_ctrl_op_fcn; // @[register-read.scala 92:29]
  reg  REG_3_ctrl_fcn_dw; // @[register-read.scala 92:29]
  reg [2:0] REG_3_ctrl_csr_cmd; // @[register-read.scala 92:29]
  reg  REG_3_ctrl_is_load; // @[register-read.scala 92:29]
  reg  REG_3_ctrl_is_sta; // @[register-read.scala 92:29]
  reg  REG_3_ctrl_is_std; // @[register-read.scala 92:29]
  reg [1:0] REG_3_ctrl_op3_sel; // @[register-read.scala 92:29]
  reg [1:0] REG_3_iw_state; // @[register-read.scala 92:29]
  reg  REG_3_iw_p1_poisoned; // @[register-read.scala 92:29]
  reg  REG_3_iw_p2_poisoned; // @[register-read.scala 92:29]
  reg  REG_3_is_br; // @[register-read.scala 92:29]
  reg  REG_3_is_jalr; // @[register-read.scala 92:29]
  reg  REG_3_is_jal; // @[register-read.scala 92:29]
  reg  REG_3_is_sfb; // @[register-read.scala 92:29]
  reg [11:0] REG_3_br_mask; // @[register-read.scala 92:29]
  reg [3:0] REG_3_br_tag; // @[register-read.scala 92:29]
  reg [4:0] REG_3_ftq_idx; // @[register-read.scala 92:29]
  reg  REG_3_edge_inst; // @[register-read.scala 92:29]
  reg [5:0] REG_3_pc_lob; // @[register-read.scala 92:29]
  reg  REG_3_taken; // @[register-read.scala 92:29]
  reg [19:0] REG_3_imm_packed; // @[register-read.scala 92:29]
  reg [11:0] REG_3_csr_addr; // @[register-read.scala 92:29]
  reg [5:0] REG_3_rob_idx; // @[register-read.scala 92:29]
  reg [4:0] REG_3_ldq_idx; // @[register-read.scala 92:29]
  reg [4:0] REG_3_stq_idx; // @[register-read.scala 92:29]
  reg [1:0] REG_3_rxq_idx; // @[register-read.scala 92:29]
  reg [6:0] REG_3_pdst; // @[register-read.scala 92:29]
  reg [6:0] REG_3_prs1; // @[register-read.scala 92:29]
  reg [6:0] REG_3_prs2; // @[register-read.scala 92:29]
  reg [6:0] REG_3_prs3; // @[register-read.scala 92:29]
  reg [4:0] REG_3_ppred; // @[register-read.scala 92:29]
  reg  REG_3_prs1_busy; // @[register-read.scala 92:29]
  reg  REG_3_prs2_busy; // @[register-read.scala 92:29]
  reg  REG_3_prs3_busy; // @[register-read.scala 92:29]
  reg  REG_3_ppred_busy; // @[register-read.scala 92:29]
  reg [6:0] REG_3_stale_pdst; // @[register-read.scala 92:29]
  reg  REG_3_exception; // @[register-read.scala 92:29]
  reg [63:0] REG_3_exc_cause; // @[register-read.scala 92:29]
  reg  REG_3_bypassable; // @[register-read.scala 92:29]
  reg [4:0] REG_3_mem_cmd; // @[register-read.scala 92:29]
  reg [1:0] REG_3_mem_size; // @[register-read.scala 92:29]
  reg  REG_3_mem_signed; // @[register-read.scala 92:29]
  reg  REG_3_is_fence; // @[register-read.scala 92:29]
  reg  REG_3_is_fencei; // @[register-read.scala 92:29]
  reg  REG_3_is_amo; // @[register-read.scala 92:29]
  reg  REG_3_uses_ldq; // @[register-read.scala 92:29]
  reg  REG_3_uses_stq; // @[register-read.scala 92:29]
  reg  REG_3_is_sys_pc2epc; // @[register-read.scala 92:29]
  reg  REG_3_is_unique; // @[register-read.scala 92:29]
  reg  REG_3_flush_on_commit; // @[register-read.scala 92:29]
  reg  REG_3_ldst_is_rs1; // @[register-read.scala 92:29]
  reg [5:0] REG_3_ldst; // @[register-read.scala 92:29]
  reg [5:0] REG_3_lrs1; // @[register-read.scala 92:29]
  reg [5:0] REG_3_lrs2; // @[register-read.scala 92:29]
  reg [5:0] REG_3_lrs3; // @[register-read.scala 92:29]
  reg  REG_3_ldst_val; // @[register-read.scala 92:29]
  reg [1:0] REG_3_dst_rtype; // @[register-read.scala 92:29]
  reg [1:0] REG_3_lrs1_rtype; // @[register-read.scala 92:29]
  reg [1:0] REG_3_lrs2_rtype; // @[register-read.scala 92:29]
  reg  REG_3_frs3_en; // @[register-read.scala 92:29]
  reg  REG_3_fp_val; // @[register-read.scala 92:29]
  reg  REG_3_fp_single; // @[register-read.scala 92:29]
  reg  REG_3_xcpt_pf_if; // @[register-read.scala 92:29]
  reg  REG_3_xcpt_ae_if; // @[register-read.scala 92:29]
  reg  REG_3_xcpt_ma_if; // @[register-read.scala 92:29]
  reg  REG_3_bp_debug_if; // @[register-read.scala 92:29]
  reg  REG_3_bp_xcpt_if; // @[register-read.scala 92:29]
  reg [1:0] REG_3_debug_fsrc; // @[register-read.scala 92:29]
  reg [1:0] REG_3_debug_tsrc; // @[register-read.scala 92:29]
  wire [11:0] _T_12 = io_brupdate_b1_mispredict_mask & RegisterReadDecode_2_io_rrd_uop_br_mask; // @[util.scala 175:51]
  wire  _T_13 = _T_12 != 12'h0; // @[util.scala 175:59]
  wire  _T_14 = ~_T_13; // @[register-read.scala 91:17]
  reg  REG_4; // @[register-read.scala 90:29]
  reg  REG_5_switch; // @[register-read.scala 92:29]
  reg  REG_5_switch_off; // @[register-read.scala 92:29]
  reg  REG_5_is_unicore; // @[register-read.scala 92:29]
  reg [2:0] REG_5_shift; // @[register-read.scala 92:29]
  reg [1:0] REG_5_lrs3_rtype; // @[register-read.scala 92:29]
  reg  REG_5_rflag; // @[register-read.scala 92:29]
  reg  REG_5_wflag; // @[register-read.scala 92:29]
  reg [3:0] REG_5_prflag; // @[register-read.scala 92:29]
  reg [3:0] REG_5_pwflag; // @[register-read.scala 92:29]
  reg  REG_5_pflag_busy; // @[register-read.scala 92:29]
  reg [3:0] REG_5_stale_pflag; // @[register-read.scala 92:29]
  reg [3:0] REG_5_op1_sel; // @[register-read.scala 92:29]
  reg [3:0] REG_5_op2_sel; // @[register-read.scala 92:29]
  reg [5:0] REG_5_split_num; // @[register-read.scala 92:29]
  reg [5:0] REG_5_self_index; // @[register-read.scala 92:29]
  reg [5:0] REG_5_rob_inst_idx; // @[register-read.scala 92:29]
  reg [5:0] REG_5_address_num; // @[register-read.scala 92:29]
  reg [6:0] REG_5_uopc; // @[register-read.scala 92:29]
  reg [31:0] REG_5_inst; // @[register-read.scala 92:29]
  reg [31:0] REG_5_debug_inst; // @[register-read.scala 92:29]
  reg  REG_5_is_rvc; // @[register-read.scala 92:29]
  reg [39:0] REG_5_debug_pc; // @[register-read.scala 92:29]
  reg [2:0] REG_5_iq_type; // @[register-read.scala 92:29]
  reg [9:0] REG_5_fu_code; // @[register-read.scala 92:29]
  reg [3:0] REG_5_ctrl_br_type; // @[register-read.scala 92:29]
  reg [1:0] REG_5_ctrl_op1_sel; // @[register-read.scala 92:29]
  reg [2:0] REG_5_ctrl_op2_sel; // @[register-read.scala 92:29]
  reg [2:0] REG_5_ctrl_imm_sel; // @[register-read.scala 92:29]
  reg [3:0] REG_5_ctrl_op_fcn; // @[register-read.scala 92:29]
  reg  REG_5_ctrl_fcn_dw; // @[register-read.scala 92:29]
  reg [2:0] REG_5_ctrl_csr_cmd; // @[register-read.scala 92:29]
  reg  REG_5_ctrl_is_load; // @[register-read.scala 92:29]
  reg  REG_5_ctrl_is_sta; // @[register-read.scala 92:29]
  reg  REG_5_ctrl_is_std; // @[register-read.scala 92:29]
  reg [1:0] REG_5_ctrl_op3_sel; // @[register-read.scala 92:29]
  reg [1:0] REG_5_iw_state; // @[register-read.scala 92:29]
  reg  REG_5_iw_p1_poisoned; // @[register-read.scala 92:29]
  reg  REG_5_iw_p2_poisoned; // @[register-read.scala 92:29]
  reg  REG_5_is_br; // @[register-read.scala 92:29]
  reg  REG_5_is_jalr; // @[register-read.scala 92:29]
  reg  REG_5_is_jal; // @[register-read.scala 92:29]
  reg  REG_5_is_sfb; // @[register-read.scala 92:29]
  reg [11:0] REG_5_br_mask; // @[register-read.scala 92:29]
  reg [3:0] REG_5_br_tag; // @[register-read.scala 92:29]
  reg [4:0] REG_5_ftq_idx; // @[register-read.scala 92:29]
  reg  REG_5_edge_inst; // @[register-read.scala 92:29]
  reg [5:0] REG_5_pc_lob; // @[register-read.scala 92:29]
  reg  REG_5_taken; // @[register-read.scala 92:29]
  reg [19:0] REG_5_imm_packed; // @[register-read.scala 92:29]
  reg [11:0] REG_5_csr_addr; // @[register-read.scala 92:29]
  reg [5:0] REG_5_rob_idx; // @[register-read.scala 92:29]
  reg [4:0] REG_5_ldq_idx; // @[register-read.scala 92:29]
  reg [4:0] REG_5_stq_idx; // @[register-read.scala 92:29]
  reg [1:0] REG_5_rxq_idx; // @[register-read.scala 92:29]
  reg [6:0] REG_5_pdst; // @[register-read.scala 92:29]
  reg [6:0] REG_5_prs1; // @[register-read.scala 92:29]
  reg [6:0] REG_5_prs2; // @[register-read.scala 92:29]
  reg [6:0] REG_5_prs3; // @[register-read.scala 92:29]
  reg [4:0] REG_5_ppred; // @[register-read.scala 92:29]
  reg  REG_5_prs1_busy; // @[register-read.scala 92:29]
  reg  REG_5_prs2_busy; // @[register-read.scala 92:29]
  reg  REG_5_prs3_busy; // @[register-read.scala 92:29]
  reg  REG_5_ppred_busy; // @[register-read.scala 92:29]
  reg [6:0] REG_5_stale_pdst; // @[register-read.scala 92:29]
  reg  REG_5_exception; // @[register-read.scala 92:29]
  reg [63:0] REG_5_exc_cause; // @[register-read.scala 92:29]
  reg  REG_5_bypassable; // @[register-read.scala 92:29]
  reg [4:0] REG_5_mem_cmd; // @[register-read.scala 92:29]
  reg [1:0] REG_5_mem_size; // @[register-read.scala 92:29]
  reg  REG_5_mem_signed; // @[register-read.scala 92:29]
  reg  REG_5_is_fence; // @[register-read.scala 92:29]
  reg  REG_5_is_fencei; // @[register-read.scala 92:29]
  reg  REG_5_is_amo; // @[register-read.scala 92:29]
  reg  REG_5_uses_ldq; // @[register-read.scala 92:29]
  reg  REG_5_uses_stq; // @[register-read.scala 92:29]
  reg  REG_5_is_sys_pc2epc; // @[register-read.scala 92:29]
  reg  REG_5_is_unique; // @[register-read.scala 92:29]
  reg  REG_5_flush_on_commit; // @[register-read.scala 92:29]
  reg  REG_5_ldst_is_rs1; // @[register-read.scala 92:29]
  reg [5:0] REG_5_ldst; // @[register-read.scala 92:29]
  reg [5:0] REG_5_lrs1; // @[register-read.scala 92:29]
  reg [5:0] REG_5_lrs2; // @[register-read.scala 92:29]
  reg [5:0] REG_5_lrs3; // @[register-read.scala 92:29]
  reg  REG_5_ldst_val; // @[register-read.scala 92:29]
  reg [1:0] REG_5_dst_rtype; // @[register-read.scala 92:29]
  reg [1:0] REG_5_lrs1_rtype; // @[register-read.scala 92:29]
  reg [1:0] REG_5_lrs2_rtype; // @[register-read.scala 92:29]
  reg  REG_5_frs3_en; // @[register-read.scala 92:29]
  reg  REG_5_fp_val; // @[register-read.scala 92:29]
  reg  REG_5_fp_single; // @[register-read.scala 92:29]
  reg  REG_5_xcpt_pf_if; // @[register-read.scala 92:29]
  reg  REG_5_xcpt_ae_if; // @[register-read.scala 92:29]
  reg  REG_5_xcpt_ma_if; // @[register-read.scala 92:29]
  reg  REG_5_bp_debug_if; // @[register-read.scala 92:29]
  reg  REG_5_bp_xcpt_if; // @[register-read.scala 92:29]
  reg [1:0] REG_5_debug_fsrc; // @[register-read.scala 92:29]
  reg [1:0] REG_5_debug_tsrc; // @[register-read.scala 92:29]
  wire  _T_19 = ~io_iss_uops_0_is_unicore; // @[register-read.scala 134:79]
  reg  REG_6; // @[register-read.scala 134:57]
  wire [63:0] rrd_rs1_data_0 = REG_6 ? 64'h0 : io_rf_read_ports_0_data; // @[register-read.scala 134:49]
  reg  REG_7; // @[register-read.scala 135:57]
  wire [63:0] rrd_rs2_data_0 = REG_7 ? 64'h0 : io_rf_read_ports_1_data; // @[register-read.scala 135:49]
  reg  REG_8; // @[register-read.scala 136:57]
  wire [63:0] rrd_rs3_data_0 = REG_8 ? 64'h0 : io_rf_read_ports_2_data; // @[register-read.scala 136:49]
  reg  REG_9; // @[register-read.scala 143:36]
  wire [3:0] rrd_flag_data_0 = REG_9 ? io_flag_rf_read_ports_0_data : 4'h0; // @[register-read.scala 143:28]
  wire [11:0] _T_32 = io_brupdate_b1_mispredict_mask & REG_1_br_mask; // @[util.scala 175:51]
  wire  _T_33 = _T_32 != 12'h0; // @[util.scala 175:59]
  wire  _T_34 = io_kill | _T_33; // @[register-read.scala 145:28]
  wire  _T_40 = ~io_iss_uops_1_is_unicore; // @[register-read.scala 134:79]
  reg  REG_10; // @[register-read.scala 134:57]
  wire [63:0] rrd_rs1_data_1 = REG_10 ? 64'h0 : io_rf_read_ports_3_data; // @[register-read.scala 134:49]
  reg  REG_11; // @[register-read.scala 135:57]
  wire [63:0] rrd_rs2_data_1 = REG_11 ? 64'h0 : io_rf_read_ports_4_data; // @[register-read.scala 135:49]
  reg  REG_12; // @[register-read.scala 136:57]
  wire [63:0] rrd_rs3_data_1 = REG_12 ? 64'h0 : io_rf_read_ports_5_data; // @[register-read.scala 136:49]
  reg  REG_13; // @[register-read.scala 143:36]
  wire [3:0] rrd_flag_data_1 = REG_13 ? io_flag_rf_read_ports_1_data : 4'h0; // @[register-read.scala 143:28]
  wire [11:0] _T_53 = io_brupdate_b1_mispredict_mask & REG_3_br_mask; // @[util.scala 175:51]
  wire  _T_54 = _T_53 != 12'h0; // @[util.scala 175:59]
  wire  _T_55 = io_kill | _T_54; // @[register-read.scala 145:28]
  wire  _T_61 = ~io_iss_uops_2_is_unicore; // @[register-read.scala 134:79]
  reg  REG_14; // @[register-read.scala 134:57]
  wire [63:0] rrd_rs1_data_2 = REG_14 ? 64'h0 : io_rf_read_ports_6_data; // @[register-read.scala 134:49]
  reg  REG_15; // @[register-read.scala 135:57]
  wire [63:0] rrd_rs2_data_2 = REG_15 ? 64'h0 : io_rf_read_ports_7_data; // @[register-read.scala 135:49]
  reg  REG_16; // @[register-read.scala 136:57]
  wire [63:0] rrd_rs3_data_2 = REG_16 ? 64'h0 : io_rf_read_ports_8_data; // @[register-read.scala 136:49]
  reg  REG_17; // @[register-read.scala 143:36]
  wire [3:0] rrd_flag_data_2 = REG_17 ? io_flag_rf_read_ports_2_data : 4'h0; // @[register-read.scala 143:28]
  wire [11:0] _T_74 = io_brupdate_b1_mispredict_mask & REG_5_br_mask; // @[util.scala 175:51]
  wire  _T_75 = _T_74 != 12'h0; // @[util.scala 175:59]
  wire  _T_76 = io_kill | _T_75; // @[register-read.scala 145:28]
  wire  _T_83 = io_bypass_0_bits_uop_dst_rtype != 2'h2; // @[micro-op.scala 184:36]
  wire  _T_84 = io_bypass_0_valid & REG_1_prs1 == io_bypass_0_bits_uop_pdst & _T_83; // @[register-read.scala 200:76]
  wire  _T_85 = io_bypass_0_bits_uop_dst_rtype == 2'h0; // @[register-read.scala 201:38]
  wire  _T_90 = _T_84 & io_bypass_0_bits_uop_dst_rtype == 2'h0 & REG_1_lrs1_rtype == 2'h0 & REG_1_prs1 != 7'h0; // @[register-read.scala 201:74]
  wire  _T_94 = io_bypass_0_valid & REG_1_prs2 == io_bypass_0_bits_uop_pdst & _T_83; // @[register-read.scala 202:76]
  wire  _T_100 = _T_94 & _T_85 & REG_1_lrs2_rtype == 2'h0 & REG_1_prs2 != 7'h0; // @[register-read.scala 203:74]
  wire  _T_104 = io_bypass_0_valid & REG_1_prs3 == io_bypass_0_bits_uop_pdst & _T_83; // @[register-read.scala 207:76]
  wire  _T_110 = _T_104 & _T_85 & REG_1_lrs3_rtype == 2'h0 & REG_1_prs3 != 7'h0; // @[register-read.scala 208:74]
  wire  _T_116 = io_bypass_0_valid & REG_1_prflag == io_bypass_0_bits_uop_pwflag & io_bypass_0_bits_uop_wflag &
    REG_1_rflag & io_bypass_0_bits_uop_is_unicore & REG_1_is_unicore; // @[register-read.scala 210:157]
  wire  _T_119 = io_bypass_1_bits_uop_dst_rtype != 2'h2; // @[micro-op.scala 184:36]
  wire  _T_120 = io_bypass_1_valid & REG_1_prs1 == io_bypass_1_bits_uop_pdst & _T_119; // @[register-read.scala 200:76]
  wire  _T_121 = io_bypass_1_bits_uop_dst_rtype == 2'h0; // @[register-read.scala 201:38]
  wire  _T_126 = _T_120 & io_bypass_1_bits_uop_dst_rtype == 2'h0 & REG_1_lrs1_rtype == 2'h0 & REG_1_prs1 != 7'h0; // @[register-read.scala 201:74]
  wire  _T_130 = io_bypass_1_valid & REG_1_prs2 == io_bypass_1_bits_uop_pdst & _T_119; // @[register-read.scala 202:76]
  wire  _T_136 = _T_130 & _T_121 & REG_1_lrs2_rtype == 2'h0 & REG_1_prs2 != 7'h0; // @[register-read.scala 203:74]
  wire  _T_140 = io_bypass_1_valid & REG_1_prs3 == io_bypass_1_bits_uop_pdst & _T_119; // @[register-read.scala 207:76]
  wire  _T_146 = _T_140 & _T_121 & REG_1_lrs3_rtype == 2'h0 & REG_1_prs3 != 7'h0; // @[register-read.scala 208:74]
  wire  _T_152 = io_bypass_1_valid & REG_1_prflag == io_bypass_1_bits_uop_pwflag & io_bypass_1_bits_uop_wflag &
    REG_1_rflag & io_bypass_1_bits_uop_is_unicore & REG_1_is_unicore; // @[register-read.scala 210:157]
  wire  _T_155 = io_bypass_2_bits_uop_dst_rtype != 2'h2; // @[micro-op.scala 184:36]
  wire  _T_156 = io_bypass_2_valid & REG_1_prs1 == io_bypass_2_bits_uop_pdst & _T_155; // @[register-read.scala 200:76]
  wire  _T_157 = io_bypass_2_bits_uop_dst_rtype == 2'h0; // @[register-read.scala 201:38]
  wire  _T_162 = _T_156 & io_bypass_2_bits_uop_dst_rtype == 2'h0 & REG_1_lrs1_rtype == 2'h0 & REG_1_prs1 != 7'h0; // @[register-read.scala 201:74]
  wire  _T_166 = io_bypass_2_valid & REG_1_prs2 == io_bypass_2_bits_uop_pdst & _T_155; // @[register-read.scala 202:76]
  wire  _T_172 = _T_166 & _T_157 & REG_1_lrs2_rtype == 2'h0 & REG_1_prs2 != 7'h0; // @[register-read.scala 203:74]
  wire  _T_176 = io_bypass_2_valid & REG_1_prs3 == io_bypass_2_bits_uop_pdst & _T_155; // @[register-read.scala 207:76]
  wire  _T_182 = _T_176 & _T_157 & REG_1_lrs3_rtype == 2'h0 & REG_1_prs3 != 7'h0; // @[register-read.scala 208:74]
  wire  _T_188 = io_bypass_2_valid & REG_1_prflag == io_bypass_2_bits_uop_pwflag & io_bypass_2_bits_uop_wflag &
    REG_1_rflag & io_bypass_2_bits_uop_is_unicore & REG_1_is_unicore; // @[register-read.scala 210:157]
  wire  _T_191 = io_bypass_3_bits_uop_dst_rtype != 2'h2; // @[micro-op.scala 184:36]
  wire  _T_192 = io_bypass_3_valid & REG_1_prs1 == io_bypass_3_bits_uop_pdst & _T_191; // @[register-read.scala 200:76]
  wire  _T_193 = io_bypass_3_bits_uop_dst_rtype == 2'h0; // @[register-read.scala 201:38]
  wire  _T_198 = _T_192 & io_bypass_3_bits_uop_dst_rtype == 2'h0 & REG_1_lrs1_rtype == 2'h0 & REG_1_prs1 != 7'h0; // @[register-read.scala 201:74]
  wire  _T_202 = io_bypass_3_valid & REG_1_prs2 == io_bypass_3_bits_uop_pdst & _T_191; // @[register-read.scala 202:76]
  wire  _T_208 = _T_202 & _T_193 & REG_1_lrs2_rtype == 2'h0 & REG_1_prs2 != 7'h0; // @[register-read.scala 203:74]
  wire  _T_212 = io_bypass_3_valid & REG_1_prs3 == io_bypass_3_bits_uop_pdst & _T_191; // @[register-read.scala 207:76]
  wire  _T_218 = _T_212 & _T_193 & REG_1_lrs3_rtype == 2'h0 & REG_1_prs3 != 7'h0; // @[register-read.scala 208:74]
  wire  _T_224 = io_bypass_3_valid & REG_1_prflag == io_bypass_3_bits_uop_pwflag & io_bypass_3_bits_uop_wflag &
    REG_1_rflag & io_bypass_3_bits_uop_is_unicore & REG_1_is_unicore; // @[register-read.scala 210:157]
  wire  _T_263 = io_bypass_0_valid & REG_3_prs1 == io_bypass_0_bits_uop_pdst & _T_83; // @[register-read.scala 200:76]
  wire  _T_269 = _T_263 & io_bypass_0_bits_uop_dst_rtype == 2'h0 & REG_3_lrs1_rtype == 2'h0 & REG_3_prs1 != 7'h0; // @[register-read.scala 201:74]
  wire  _T_273 = io_bypass_0_valid & REG_3_prs2 == io_bypass_0_bits_uop_pdst & _T_83; // @[register-read.scala 202:76]
  wire  _T_279 = _T_273 & _T_85 & REG_3_lrs2_rtype == 2'h0 & REG_3_prs2 != 7'h0; // @[register-read.scala 203:74]
  wire  _T_283 = io_bypass_0_valid & REG_3_prs3 == io_bypass_0_bits_uop_pdst & _T_83; // @[register-read.scala 207:76]
  wire  _T_289 = _T_283 & _T_85 & REG_3_lrs3_rtype == 2'h0 & REG_3_prs3 != 7'h0; // @[register-read.scala 208:74]
  wire  _T_295 = io_bypass_0_valid & REG_3_prflag == io_bypass_0_bits_uop_pwflag & io_bypass_0_bits_uop_wflag &
    REG_3_rflag & io_bypass_0_bits_uop_is_unicore & REG_3_is_unicore; // @[register-read.scala 210:157]
  wire  _T_299 = io_bypass_1_valid & REG_3_prs1 == io_bypass_1_bits_uop_pdst & _T_119; // @[register-read.scala 200:76]
  wire  _T_305 = _T_299 & io_bypass_1_bits_uop_dst_rtype == 2'h0 & REG_3_lrs1_rtype == 2'h0 & REG_3_prs1 != 7'h0; // @[register-read.scala 201:74]
  wire  _T_309 = io_bypass_1_valid & REG_3_prs2 == io_bypass_1_bits_uop_pdst & _T_119; // @[register-read.scala 202:76]
  wire  _T_315 = _T_309 & _T_121 & REG_3_lrs2_rtype == 2'h0 & REG_3_prs2 != 7'h0; // @[register-read.scala 203:74]
  wire  _T_319 = io_bypass_1_valid & REG_3_prs3 == io_bypass_1_bits_uop_pdst & _T_119; // @[register-read.scala 207:76]
  wire  _T_325 = _T_319 & _T_121 & REG_3_lrs3_rtype == 2'h0 & REG_3_prs3 != 7'h0; // @[register-read.scala 208:74]
  wire  _T_331 = io_bypass_1_valid & REG_3_prflag == io_bypass_1_bits_uop_pwflag & io_bypass_1_bits_uop_wflag &
    REG_3_rflag & io_bypass_1_bits_uop_is_unicore & REG_3_is_unicore; // @[register-read.scala 210:157]
  wire  _T_335 = io_bypass_2_valid & REG_3_prs1 == io_bypass_2_bits_uop_pdst & _T_155; // @[register-read.scala 200:76]
  wire  _T_341 = _T_335 & io_bypass_2_bits_uop_dst_rtype == 2'h0 & REG_3_lrs1_rtype == 2'h0 & REG_3_prs1 != 7'h0; // @[register-read.scala 201:74]
  wire  _T_345 = io_bypass_2_valid & REG_3_prs2 == io_bypass_2_bits_uop_pdst & _T_155; // @[register-read.scala 202:76]
  wire  _T_351 = _T_345 & _T_157 & REG_3_lrs2_rtype == 2'h0 & REG_3_prs2 != 7'h0; // @[register-read.scala 203:74]
  wire  _T_355 = io_bypass_2_valid & REG_3_prs3 == io_bypass_2_bits_uop_pdst & _T_155; // @[register-read.scala 207:76]
  wire  _T_361 = _T_355 & _T_157 & REG_3_lrs3_rtype == 2'h0 & REG_3_prs3 != 7'h0; // @[register-read.scala 208:74]
  wire  _T_367 = io_bypass_2_valid & REG_3_prflag == io_bypass_2_bits_uop_pwflag & io_bypass_2_bits_uop_wflag &
    REG_3_rflag & io_bypass_2_bits_uop_is_unicore & REG_3_is_unicore; // @[register-read.scala 210:157]
  wire  _T_371 = io_bypass_3_valid & REG_3_prs1 == io_bypass_3_bits_uop_pdst & _T_191; // @[register-read.scala 200:76]
  wire  _T_377 = _T_371 & io_bypass_3_bits_uop_dst_rtype == 2'h0 & REG_3_lrs1_rtype == 2'h0 & REG_3_prs1 != 7'h0; // @[register-read.scala 201:74]
  wire  _T_381 = io_bypass_3_valid & REG_3_prs2 == io_bypass_3_bits_uop_pdst & _T_191; // @[register-read.scala 202:76]
  wire  _T_387 = _T_381 & _T_193 & REG_3_lrs2_rtype == 2'h0 & REG_3_prs2 != 7'h0; // @[register-read.scala 203:74]
  wire  _T_391 = io_bypass_3_valid & REG_3_prs3 == io_bypass_3_bits_uop_pdst & _T_191; // @[register-read.scala 207:76]
  wire  _T_397 = _T_391 & _T_193 & REG_3_lrs3_rtype == 2'h0 & REG_3_prs3 != 7'h0; // @[register-read.scala 208:74]
  wire  _T_403 = io_bypass_3_valid & REG_3_prflag == io_bypass_3_bits_uop_pwflag & io_bypass_3_bits_uop_wflag &
    REG_3_rflag & io_bypass_3_bits_uop_is_unicore & REG_3_is_unicore; // @[register-read.scala 210:157]
  wire  _T_442 = io_bypass_0_valid & REG_5_prs1 == io_bypass_0_bits_uop_pdst & _T_83; // @[register-read.scala 200:76]
  wire  _T_448 = _T_442 & io_bypass_0_bits_uop_dst_rtype == 2'h0 & REG_5_lrs1_rtype == 2'h0 & REG_5_prs1 != 7'h0; // @[register-read.scala 201:74]
  wire  _T_452 = io_bypass_0_valid & REG_5_prs2 == io_bypass_0_bits_uop_pdst & _T_83; // @[register-read.scala 202:76]
  wire  _T_458 = _T_452 & _T_85 & REG_5_lrs2_rtype == 2'h0 & REG_5_prs2 != 7'h0; // @[register-read.scala 203:74]
  wire  _T_462 = io_bypass_0_valid & REG_5_prs3 == io_bypass_0_bits_uop_pdst & _T_83; // @[register-read.scala 207:76]
  wire  _T_468 = _T_462 & _T_85 & REG_5_lrs3_rtype == 2'h0 & REG_5_prs3 != 7'h0; // @[register-read.scala 208:74]
  wire  _T_474 = io_bypass_0_valid & REG_5_prflag == io_bypass_0_bits_uop_pwflag & io_bypass_0_bits_uop_wflag &
    REG_5_rflag & io_bypass_0_bits_uop_is_unicore & REG_5_is_unicore; // @[register-read.scala 210:157]
  wire  _T_478 = io_bypass_1_valid & REG_5_prs1 == io_bypass_1_bits_uop_pdst & _T_119; // @[register-read.scala 200:76]
  wire  _T_484 = _T_478 & io_bypass_1_bits_uop_dst_rtype == 2'h0 & REG_5_lrs1_rtype == 2'h0 & REG_5_prs1 != 7'h0; // @[register-read.scala 201:74]
  wire  _T_488 = io_bypass_1_valid & REG_5_prs2 == io_bypass_1_bits_uop_pdst & _T_119; // @[register-read.scala 202:76]
  wire  _T_494 = _T_488 & _T_121 & REG_5_lrs2_rtype == 2'h0 & REG_5_prs2 != 7'h0; // @[register-read.scala 203:74]
  wire  _T_498 = io_bypass_1_valid & REG_5_prs3 == io_bypass_1_bits_uop_pdst & _T_119; // @[register-read.scala 207:76]
  wire  _T_504 = _T_498 & _T_121 & REG_5_lrs3_rtype == 2'h0 & REG_5_prs3 != 7'h0; // @[register-read.scala 208:74]
  wire  _T_510 = io_bypass_1_valid & REG_5_prflag == io_bypass_1_bits_uop_pwflag & io_bypass_1_bits_uop_wflag &
    REG_5_rflag & io_bypass_1_bits_uop_is_unicore & REG_5_is_unicore; // @[register-read.scala 210:157]
  wire  _T_514 = io_bypass_2_valid & REG_5_prs1 == io_bypass_2_bits_uop_pdst & _T_155; // @[register-read.scala 200:76]
  wire  _T_520 = _T_514 & io_bypass_2_bits_uop_dst_rtype == 2'h0 & REG_5_lrs1_rtype == 2'h0 & REG_5_prs1 != 7'h0; // @[register-read.scala 201:74]
  wire  _T_524 = io_bypass_2_valid & REG_5_prs2 == io_bypass_2_bits_uop_pdst & _T_155; // @[register-read.scala 202:76]
  wire  _T_530 = _T_524 & _T_157 & REG_5_lrs2_rtype == 2'h0 & REG_5_prs2 != 7'h0; // @[register-read.scala 203:74]
  wire  _T_534 = io_bypass_2_valid & REG_5_prs3 == io_bypass_2_bits_uop_pdst & _T_155; // @[register-read.scala 207:76]
  wire  _T_540 = _T_534 & _T_157 & REG_5_lrs3_rtype == 2'h0 & REG_5_prs3 != 7'h0; // @[register-read.scala 208:74]
  wire  _T_546 = io_bypass_2_valid & REG_5_prflag == io_bypass_2_bits_uop_pwflag & io_bypass_2_bits_uop_wflag &
    REG_5_rflag & io_bypass_2_bits_uop_is_unicore & REG_5_is_unicore; // @[register-read.scala 210:157]
  wire  _T_550 = io_bypass_3_valid & REG_5_prs1 == io_bypass_3_bits_uop_pdst & _T_191; // @[register-read.scala 200:76]
  wire  _T_556 = _T_550 & io_bypass_3_bits_uop_dst_rtype == 2'h0 & REG_5_lrs1_rtype == 2'h0 & REG_5_prs1 != 7'h0; // @[register-read.scala 201:74]
  wire  _T_560 = io_bypass_3_valid & REG_5_prs2 == io_bypass_3_bits_uop_pdst & _T_191; // @[register-read.scala 202:76]
  wire  _T_566 = _T_560 & _T_193 & REG_5_lrs2_rtype == 2'h0 & REG_5_prs2 != 7'h0; // @[register-read.scala 203:74]
  wire  _T_570 = io_bypass_3_valid & REG_5_prs3 == io_bypass_3_bits_uop_pdst & _T_191; // @[register-read.scala 207:76]
  wire  _T_576 = _T_570 & _T_193 & REG_5_lrs3_rtype == 2'h0 & REG_5_prs3 != 7'h0; // @[register-read.scala 208:74]
  wire  _T_582 = io_bypass_3_valid & REG_5_prflag == io_bypass_3_bits_uop_pwflag & io_bypass_3_bits_uop_wflag &
    REG_5_rflag & io_bypass_3_bits_uop_is_unicore & REG_5_is_unicore; // @[register-read.scala 210:157]
  RegisterReadDecode_1 RegisterReadDecode ( // @[register-read.scala 86:33]
    .clock(RegisterReadDecode_clock),
    .reset(RegisterReadDecode_reset),
    .io_iss_valid(RegisterReadDecode_io_iss_valid),
    .io_iss_uop_switch(RegisterReadDecode_io_iss_uop_switch),
    .io_iss_uop_switch_off(RegisterReadDecode_io_iss_uop_switch_off),
    .io_iss_uop_is_unicore(RegisterReadDecode_io_iss_uop_is_unicore),
    .io_iss_uop_shift(RegisterReadDecode_io_iss_uop_shift),
    .io_iss_uop_lrs3_rtype(RegisterReadDecode_io_iss_uop_lrs3_rtype),
    .io_iss_uop_rflag(RegisterReadDecode_io_iss_uop_rflag),
    .io_iss_uop_wflag(RegisterReadDecode_io_iss_uop_wflag),
    .io_iss_uop_prflag(RegisterReadDecode_io_iss_uop_prflag),
    .io_iss_uop_pwflag(RegisterReadDecode_io_iss_uop_pwflag),
    .io_iss_uop_pflag_busy(RegisterReadDecode_io_iss_uop_pflag_busy),
    .io_iss_uop_stale_pflag(RegisterReadDecode_io_iss_uop_stale_pflag),
    .io_iss_uop_op1_sel(RegisterReadDecode_io_iss_uop_op1_sel),
    .io_iss_uop_op2_sel(RegisterReadDecode_io_iss_uop_op2_sel),
    .io_iss_uop_split_num(RegisterReadDecode_io_iss_uop_split_num),
    .io_iss_uop_self_index(RegisterReadDecode_io_iss_uop_self_index),
    .io_iss_uop_rob_inst_idx(RegisterReadDecode_io_iss_uop_rob_inst_idx),
    .io_iss_uop_address_num(RegisterReadDecode_io_iss_uop_address_num),
    .io_iss_uop_uopc(RegisterReadDecode_io_iss_uop_uopc),
    .io_iss_uop_inst(RegisterReadDecode_io_iss_uop_inst),
    .io_iss_uop_debug_inst(RegisterReadDecode_io_iss_uop_debug_inst),
    .io_iss_uop_is_rvc(RegisterReadDecode_io_iss_uop_is_rvc),
    .io_iss_uop_debug_pc(RegisterReadDecode_io_iss_uop_debug_pc),
    .io_iss_uop_iq_type(RegisterReadDecode_io_iss_uop_iq_type),
    .io_iss_uop_fu_code(RegisterReadDecode_io_iss_uop_fu_code),
    .io_iss_uop_ctrl_br_type(RegisterReadDecode_io_iss_uop_ctrl_br_type),
    .io_iss_uop_ctrl_op1_sel(RegisterReadDecode_io_iss_uop_ctrl_op1_sel),
    .io_iss_uop_ctrl_op2_sel(RegisterReadDecode_io_iss_uop_ctrl_op2_sel),
    .io_iss_uop_ctrl_imm_sel(RegisterReadDecode_io_iss_uop_ctrl_imm_sel),
    .io_iss_uop_ctrl_op_fcn(RegisterReadDecode_io_iss_uop_ctrl_op_fcn),
    .io_iss_uop_ctrl_fcn_dw(RegisterReadDecode_io_iss_uop_ctrl_fcn_dw),
    .io_iss_uop_ctrl_csr_cmd(RegisterReadDecode_io_iss_uop_ctrl_csr_cmd),
    .io_iss_uop_ctrl_is_load(RegisterReadDecode_io_iss_uop_ctrl_is_load),
    .io_iss_uop_ctrl_is_sta(RegisterReadDecode_io_iss_uop_ctrl_is_sta),
    .io_iss_uop_ctrl_is_std(RegisterReadDecode_io_iss_uop_ctrl_is_std),
    .io_iss_uop_ctrl_op3_sel(RegisterReadDecode_io_iss_uop_ctrl_op3_sel),
    .io_iss_uop_iw_state(RegisterReadDecode_io_iss_uop_iw_state),
    .io_iss_uop_iw_p1_poisoned(RegisterReadDecode_io_iss_uop_iw_p1_poisoned),
    .io_iss_uop_iw_p2_poisoned(RegisterReadDecode_io_iss_uop_iw_p2_poisoned),
    .io_iss_uop_is_br(RegisterReadDecode_io_iss_uop_is_br),
    .io_iss_uop_is_jalr(RegisterReadDecode_io_iss_uop_is_jalr),
    .io_iss_uop_is_jal(RegisterReadDecode_io_iss_uop_is_jal),
    .io_iss_uop_is_sfb(RegisterReadDecode_io_iss_uop_is_sfb),
    .io_iss_uop_br_mask(RegisterReadDecode_io_iss_uop_br_mask),
    .io_iss_uop_br_tag(RegisterReadDecode_io_iss_uop_br_tag),
    .io_iss_uop_ftq_idx(RegisterReadDecode_io_iss_uop_ftq_idx),
    .io_iss_uop_edge_inst(RegisterReadDecode_io_iss_uop_edge_inst),
    .io_iss_uop_pc_lob(RegisterReadDecode_io_iss_uop_pc_lob),
    .io_iss_uop_taken(RegisterReadDecode_io_iss_uop_taken),
    .io_iss_uop_imm_packed(RegisterReadDecode_io_iss_uop_imm_packed),
    .io_iss_uop_csr_addr(RegisterReadDecode_io_iss_uop_csr_addr),
    .io_iss_uop_rob_idx(RegisterReadDecode_io_iss_uop_rob_idx),
    .io_iss_uop_ldq_idx(RegisterReadDecode_io_iss_uop_ldq_idx),
    .io_iss_uop_stq_idx(RegisterReadDecode_io_iss_uop_stq_idx),
    .io_iss_uop_rxq_idx(RegisterReadDecode_io_iss_uop_rxq_idx),
    .io_iss_uop_pdst(RegisterReadDecode_io_iss_uop_pdst),
    .io_iss_uop_prs1(RegisterReadDecode_io_iss_uop_prs1),
    .io_iss_uop_prs2(RegisterReadDecode_io_iss_uop_prs2),
    .io_iss_uop_prs3(RegisterReadDecode_io_iss_uop_prs3),
    .io_iss_uop_ppred(RegisterReadDecode_io_iss_uop_ppred),
    .io_iss_uop_prs1_busy(RegisterReadDecode_io_iss_uop_prs1_busy),
    .io_iss_uop_prs2_busy(RegisterReadDecode_io_iss_uop_prs2_busy),
    .io_iss_uop_prs3_busy(RegisterReadDecode_io_iss_uop_prs3_busy),
    .io_iss_uop_ppred_busy(RegisterReadDecode_io_iss_uop_ppred_busy),
    .io_iss_uop_stale_pdst(RegisterReadDecode_io_iss_uop_stale_pdst),
    .io_iss_uop_exception(RegisterReadDecode_io_iss_uop_exception),
    .io_iss_uop_exc_cause(RegisterReadDecode_io_iss_uop_exc_cause),
    .io_iss_uop_bypassable(RegisterReadDecode_io_iss_uop_bypassable),
    .io_iss_uop_mem_cmd(RegisterReadDecode_io_iss_uop_mem_cmd),
    .io_iss_uop_mem_size(RegisterReadDecode_io_iss_uop_mem_size),
    .io_iss_uop_mem_signed(RegisterReadDecode_io_iss_uop_mem_signed),
    .io_iss_uop_is_fence(RegisterReadDecode_io_iss_uop_is_fence),
    .io_iss_uop_is_fencei(RegisterReadDecode_io_iss_uop_is_fencei),
    .io_iss_uop_is_amo(RegisterReadDecode_io_iss_uop_is_amo),
    .io_iss_uop_uses_ldq(RegisterReadDecode_io_iss_uop_uses_ldq),
    .io_iss_uop_uses_stq(RegisterReadDecode_io_iss_uop_uses_stq),
    .io_iss_uop_is_sys_pc2epc(RegisterReadDecode_io_iss_uop_is_sys_pc2epc),
    .io_iss_uop_is_unique(RegisterReadDecode_io_iss_uop_is_unique),
    .io_iss_uop_flush_on_commit(RegisterReadDecode_io_iss_uop_flush_on_commit),
    .io_iss_uop_ldst_is_rs1(RegisterReadDecode_io_iss_uop_ldst_is_rs1),
    .io_iss_uop_ldst(RegisterReadDecode_io_iss_uop_ldst),
    .io_iss_uop_lrs1(RegisterReadDecode_io_iss_uop_lrs1),
    .io_iss_uop_lrs2(RegisterReadDecode_io_iss_uop_lrs2),
    .io_iss_uop_lrs3(RegisterReadDecode_io_iss_uop_lrs3),
    .io_iss_uop_ldst_val(RegisterReadDecode_io_iss_uop_ldst_val),
    .io_iss_uop_dst_rtype(RegisterReadDecode_io_iss_uop_dst_rtype),
    .io_iss_uop_lrs1_rtype(RegisterReadDecode_io_iss_uop_lrs1_rtype),
    .io_iss_uop_lrs2_rtype(RegisterReadDecode_io_iss_uop_lrs2_rtype),
    .io_iss_uop_frs3_en(RegisterReadDecode_io_iss_uop_frs3_en),
    .io_iss_uop_fp_val(RegisterReadDecode_io_iss_uop_fp_val),
    .io_iss_uop_fp_single(RegisterReadDecode_io_iss_uop_fp_single),
    .io_iss_uop_xcpt_pf_if(RegisterReadDecode_io_iss_uop_xcpt_pf_if),
    .io_iss_uop_xcpt_ae_if(RegisterReadDecode_io_iss_uop_xcpt_ae_if),
    .io_iss_uop_xcpt_ma_if(RegisterReadDecode_io_iss_uop_xcpt_ma_if),
    .io_iss_uop_bp_debug_if(RegisterReadDecode_io_iss_uop_bp_debug_if),
    .io_iss_uop_bp_xcpt_if(RegisterReadDecode_io_iss_uop_bp_xcpt_if),
    .io_iss_uop_debug_fsrc(RegisterReadDecode_io_iss_uop_debug_fsrc),
    .io_iss_uop_debug_tsrc(RegisterReadDecode_io_iss_uop_debug_tsrc),
    .io_rrd_valid(RegisterReadDecode_io_rrd_valid),
    .io_rrd_uop_switch(RegisterReadDecode_io_rrd_uop_switch),
    .io_rrd_uop_switch_off(RegisterReadDecode_io_rrd_uop_switch_off),
    .io_rrd_uop_is_unicore(RegisterReadDecode_io_rrd_uop_is_unicore),
    .io_rrd_uop_shift(RegisterReadDecode_io_rrd_uop_shift),
    .io_rrd_uop_lrs3_rtype(RegisterReadDecode_io_rrd_uop_lrs3_rtype),
    .io_rrd_uop_rflag(RegisterReadDecode_io_rrd_uop_rflag),
    .io_rrd_uop_wflag(RegisterReadDecode_io_rrd_uop_wflag),
    .io_rrd_uop_prflag(RegisterReadDecode_io_rrd_uop_prflag),
    .io_rrd_uop_pwflag(RegisterReadDecode_io_rrd_uop_pwflag),
    .io_rrd_uop_pflag_busy(RegisterReadDecode_io_rrd_uop_pflag_busy),
    .io_rrd_uop_stale_pflag(RegisterReadDecode_io_rrd_uop_stale_pflag),
    .io_rrd_uop_op1_sel(RegisterReadDecode_io_rrd_uop_op1_sel),
    .io_rrd_uop_op2_sel(RegisterReadDecode_io_rrd_uop_op2_sel),
    .io_rrd_uop_split_num(RegisterReadDecode_io_rrd_uop_split_num),
    .io_rrd_uop_self_index(RegisterReadDecode_io_rrd_uop_self_index),
    .io_rrd_uop_rob_inst_idx(RegisterReadDecode_io_rrd_uop_rob_inst_idx),
    .io_rrd_uop_address_num(RegisterReadDecode_io_rrd_uop_address_num),
    .io_rrd_uop_uopc(RegisterReadDecode_io_rrd_uop_uopc),
    .io_rrd_uop_inst(RegisterReadDecode_io_rrd_uop_inst),
    .io_rrd_uop_debug_inst(RegisterReadDecode_io_rrd_uop_debug_inst),
    .io_rrd_uop_is_rvc(RegisterReadDecode_io_rrd_uop_is_rvc),
    .io_rrd_uop_debug_pc(RegisterReadDecode_io_rrd_uop_debug_pc),
    .io_rrd_uop_iq_type(RegisterReadDecode_io_rrd_uop_iq_type),
    .io_rrd_uop_fu_code(RegisterReadDecode_io_rrd_uop_fu_code),
    .io_rrd_uop_ctrl_br_type(RegisterReadDecode_io_rrd_uop_ctrl_br_type),
    .io_rrd_uop_ctrl_op1_sel(RegisterReadDecode_io_rrd_uop_ctrl_op1_sel),
    .io_rrd_uop_ctrl_op2_sel(RegisterReadDecode_io_rrd_uop_ctrl_op2_sel),
    .io_rrd_uop_ctrl_imm_sel(RegisterReadDecode_io_rrd_uop_ctrl_imm_sel),
    .io_rrd_uop_ctrl_op_fcn(RegisterReadDecode_io_rrd_uop_ctrl_op_fcn),
    .io_rrd_uop_ctrl_fcn_dw(RegisterReadDecode_io_rrd_uop_ctrl_fcn_dw),
    .io_rrd_uop_ctrl_csr_cmd(RegisterReadDecode_io_rrd_uop_ctrl_csr_cmd),
    .io_rrd_uop_ctrl_is_load(RegisterReadDecode_io_rrd_uop_ctrl_is_load),
    .io_rrd_uop_ctrl_is_sta(RegisterReadDecode_io_rrd_uop_ctrl_is_sta),
    .io_rrd_uop_ctrl_is_std(RegisterReadDecode_io_rrd_uop_ctrl_is_std),
    .io_rrd_uop_ctrl_op3_sel(RegisterReadDecode_io_rrd_uop_ctrl_op3_sel),
    .io_rrd_uop_iw_state(RegisterReadDecode_io_rrd_uop_iw_state),
    .io_rrd_uop_iw_p1_poisoned(RegisterReadDecode_io_rrd_uop_iw_p1_poisoned),
    .io_rrd_uop_iw_p2_poisoned(RegisterReadDecode_io_rrd_uop_iw_p2_poisoned),
    .io_rrd_uop_is_br(RegisterReadDecode_io_rrd_uop_is_br),
    .io_rrd_uop_is_jalr(RegisterReadDecode_io_rrd_uop_is_jalr),
    .io_rrd_uop_is_jal(RegisterReadDecode_io_rrd_uop_is_jal),
    .io_rrd_uop_is_sfb(RegisterReadDecode_io_rrd_uop_is_sfb),
    .io_rrd_uop_br_mask(RegisterReadDecode_io_rrd_uop_br_mask),
    .io_rrd_uop_br_tag(RegisterReadDecode_io_rrd_uop_br_tag),
    .io_rrd_uop_ftq_idx(RegisterReadDecode_io_rrd_uop_ftq_idx),
    .io_rrd_uop_edge_inst(RegisterReadDecode_io_rrd_uop_edge_inst),
    .io_rrd_uop_pc_lob(RegisterReadDecode_io_rrd_uop_pc_lob),
    .io_rrd_uop_taken(RegisterReadDecode_io_rrd_uop_taken),
    .io_rrd_uop_imm_packed(RegisterReadDecode_io_rrd_uop_imm_packed),
    .io_rrd_uop_csr_addr(RegisterReadDecode_io_rrd_uop_csr_addr),
    .io_rrd_uop_rob_idx(RegisterReadDecode_io_rrd_uop_rob_idx),
    .io_rrd_uop_ldq_idx(RegisterReadDecode_io_rrd_uop_ldq_idx),
    .io_rrd_uop_stq_idx(RegisterReadDecode_io_rrd_uop_stq_idx),
    .io_rrd_uop_rxq_idx(RegisterReadDecode_io_rrd_uop_rxq_idx),
    .io_rrd_uop_pdst(RegisterReadDecode_io_rrd_uop_pdst),
    .io_rrd_uop_prs1(RegisterReadDecode_io_rrd_uop_prs1),
    .io_rrd_uop_prs2(RegisterReadDecode_io_rrd_uop_prs2),
    .io_rrd_uop_prs3(RegisterReadDecode_io_rrd_uop_prs3),
    .io_rrd_uop_ppred(RegisterReadDecode_io_rrd_uop_ppred),
    .io_rrd_uop_prs1_busy(RegisterReadDecode_io_rrd_uop_prs1_busy),
    .io_rrd_uop_prs2_busy(RegisterReadDecode_io_rrd_uop_prs2_busy),
    .io_rrd_uop_prs3_busy(RegisterReadDecode_io_rrd_uop_prs3_busy),
    .io_rrd_uop_ppred_busy(RegisterReadDecode_io_rrd_uop_ppred_busy),
    .io_rrd_uop_stale_pdst(RegisterReadDecode_io_rrd_uop_stale_pdst),
    .io_rrd_uop_exception(RegisterReadDecode_io_rrd_uop_exception),
    .io_rrd_uop_exc_cause(RegisterReadDecode_io_rrd_uop_exc_cause),
    .io_rrd_uop_bypassable(RegisterReadDecode_io_rrd_uop_bypassable),
    .io_rrd_uop_mem_cmd(RegisterReadDecode_io_rrd_uop_mem_cmd),
    .io_rrd_uop_mem_size(RegisterReadDecode_io_rrd_uop_mem_size),
    .io_rrd_uop_mem_signed(RegisterReadDecode_io_rrd_uop_mem_signed),
    .io_rrd_uop_is_fence(RegisterReadDecode_io_rrd_uop_is_fence),
    .io_rrd_uop_is_fencei(RegisterReadDecode_io_rrd_uop_is_fencei),
    .io_rrd_uop_is_amo(RegisterReadDecode_io_rrd_uop_is_amo),
    .io_rrd_uop_uses_ldq(RegisterReadDecode_io_rrd_uop_uses_ldq),
    .io_rrd_uop_uses_stq(RegisterReadDecode_io_rrd_uop_uses_stq),
    .io_rrd_uop_is_sys_pc2epc(RegisterReadDecode_io_rrd_uop_is_sys_pc2epc),
    .io_rrd_uop_is_unique(RegisterReadDecode_io_rrd_uop_is_unique),
    .io_rrd_uop_flush_on_commit(RegisterReadDecode_io_rrd_uop_flush_on_commit),
    .io_rrd_uop_ldst_is_rs1(RegisterReadDecode_io_rrd_uop_ldst_is_rs1),
    .io_rrd_uop_ldst(RegisterReadDecode_io_rrd_uop_ldst),
    .io_rrd_uop_lrs1(RegisterReadDecode_io_rrd_uop_lrs1),
    .io_rrd_uop_lrs2(RegisterReadDecode_io_rrd_uop_lrs2),
    .io_rrd_uop_lrs3(RegisterReadDecode_io_rrd_uop_lrs3),
    .io_rrd_uop_ldst_val(RegisterReadDecode_io_rrd_uop_ldst_val),
    .io_rrd_uop_dst_rtype(RegisterReadDecode_io_rrd_uop_dst_rtype),
    .io_rrd_uop_lrs1_rtype(RegisterReadDecode_io_rrd_uop_lrs1_rtype),
    .io_rrd_uop_lrs2_rtype(RegisterReadDecode_io_rrd_uop_lrs2_rtype),
    .io_rrd_uop_frs3_en(RegisterReadDecode_io_rrd_uop_frs3_en),
    .io_rrd_uop_fp_val(RegisterReadDecode_io_rrd_uop_fp_val),
    .io_rrd_uop_fp_single(RegisterReadDecode_io_rrd_uop_fp_single),
    .io_rrd_uop_xcpt_pf_if(RegisterReadDecode_io_rrd_uop_xcpt_pf_if),
    .io_rrd_uop_xcpt_ae_if(RegisterReadDecode_io_rrd_uop_xcpt_ae_if),
    .io_rrd_uop_xcpt_ma_if(RegisterReadDecode_io_rrd_uop_xcpt_ma_if),
    .io_rrd_uop_bp_debug_if(RegisterReadDecode_io_rrd_uop_bp_debug_if),
    .io_rrd_uop_bp_xcpt_if(RegisterReadDecode_io_rrd_uop_bp_xcpt_if),
    .io_rrd_uop_debug_fsrc(RegisterReadDecode_io_rrd_uop_debug_fsrc),
    .io_rrd_uop_debug_tsrc(RegisterReadDecode_io_rrd_uop_debug_tsrc)
  );
  RegisterReadDecode_2 RegisterReadDecode_1 ( // @[register-read.scala 86:33]
    .clock(RegisterReadDecode_1_clock),
    .reset(RegisterReadDecode_1_reset),
    .io_iss_valid(RegisterReadDecode_1_io_iss_valid),
    .io_iss_uop_switch(RegisterReadDecode_1_io_iss_uop_switch),
    .io_iss_uop_switch_off(RegisterReadDecode_1_io_iss_uop_switch_off),
    .io_iss_uop_is_unicore(RegisterReadDecode_1_io_iss_uop_is_unicore),
    .io_iss_uop_shift(RegisterReadDecode_1_io_iss_uop_shift),
    .io_iss_uop_lrs3_rtype(RegisterReadDecode_1_io_iss_uop_lrs3_rtype),
    .io_iss_uop_rflag(RegisterReadDecode_1_io_iss_uop_rflag),
    .io_iss_uop_wflag(RegisterReadDecode_1_io_iss_uop_wflag),
    .io_iss_uop_prflag(RegisterReadDecode_1_io_iss_uop_prflag),
    .io_iss_uop_pwflag(RegisterReadDecode_1_io_iss_uop_pwflag),
    .io_iss_uop_pflag_busy(RegisterReadDecode_1_io_iss_uop_pflag_busy),
    .io_iss_uop_stale_pflag(RegisterReadDecode_1_io_iss_uop_stale_pflag),
    .io_iss_uop_op1_sel(RegisterReadDecode_1_io_iss_uop_op1_sel),
    .io_iss_uop_op2_sel(RegisterReadDecode_1_io_iss_uop_op2_sel),
    .io_iss_uop_split_num(RegisterReadDecode_1_io_iss_uop_split_num),
    .io_iss_uop_self_index(RegisterReadDecode_1_io_iss_uop_self_index),
    .io_iss_uop_rob_inst_idx(RegisterReadDecode_1_io_iss_uop_rob_inst_idx),
    .io_iss_uop_address_num(RegisterReadDecode_1_io_iss_uop_address_num),
    .io_iss_uop_uopc(RegisterReadDecode_1_io_iss_uop_uopc),
    .io_iss_uop_inst(RegisterReadDecode_1_io_iss_uop_inst),
    .io_iss_uop_debug_inst(RegisterReadDecode_1_io_iss_uop_debug_inst),
    .io_iss_uop_is_rvc(RegisterReadDecode_1_io_iss_uop_is_rvc),
    .io_iss_uop_debug_pc(RegisterReadDecode_1_io_iss_uop_debug_pc),
    .io_iss_uop_iq_type(RegisterReadDecode_1_io_iss_uop_iq_type),
    .io_iss_uop_fu_code(RegisterReadDecode_1_io_iss_uop_fu_code),
    .io_iss_uop_ctrl_br_type(RegisterReadDecode_1_io_iss_uop_ctrl_br_type),
    .io_iss_uop_ctrl_op1_sel(RegisterReadDecode_1_io_iss_uop_ctrl_op1_sel),
    .io_iss_uop_ctrl_op2_sel(RegisterReadDecode_1_io_iss_uop_ctrl_op2_sel),
    .io_iss_uop_ctrl_imm_sel(RegisterReadDecode_1_io_iss_uop_ctrl_imm_sel),
    .io_iss_uop_ctrl_op_fcn(RegisterReadDecode_1_io_iss_uop_ctrl_op_fcn),
    .io_iss_uop_ctrl_fcn_dw(RegisterReadDecode_1_io_iss_uop_ctrl_fcn_dw),
    .io_iss_uop_ctrl_csr_cmd(RegisterReadDecode_1_io_iss_uop_ctrl_csr_cmd),
    .io_iss_uop_ctrl_is_load(RegisterReadDecode_1_io_iss_uop_ctrl_is_load),
    .io_iss_uop_ctrl_is_sta(RegisterReadDecode_1_io_iss_uop_ctrl_is_sta),
    .io_iss_uop_ctrl_is_std(RegisterReadDecode_1_io_iss_uop_ctrl_is_std),
    .io_iss_uop_ctrl_op3_sel(RegisterReadDecode_1_io_iss_uop_ctrl_op3_sel),
    .io_iss_uop_iw_state(RegisterReadDecode_1_io_iss_uop_iw_state),
    .io_iss_uop_iw_p1_poisoned(RegisterReadDecode_1_io_iss_uop_iw_p1_poisoned),
    .io_iss_uop_iw_p2_poisoned(RegisterReadDecode_1_io_iss_uop_iw_p2_poisoned),
    .io_iss_uop_is_br(RegisterReadDecode_1_io_iss_uop_is_br),
    .io_iss_uop_is_jalr(RegisterReadDecode_1_io_iss_uop_is_jalr),
    .io_iss_uop_is_jal(RegisterReadDecode_1_io_iss_uop_is_jal),
    .io_iss_uop_is_sfb(RegisterReadDecode_1_io_iss_uop_is_sfb),
    .io_iss_uop_br_mask(RegisterReadDecode_1_io_iss_uop_br_mask),
    .io_iss_uop_br_tag(RegisterReadDecode_1_io_iss_uop_br_tag),
    .io_iss_uop_ftq_idx(RegisterReadDecode_1_io_iss_uop_ftq_idx),
    .io_iss_uop_edge_inst(RegisterReadDecode_1_io_iss_uop_edge_inst),
    .io_iss_uop_pc_lob(RegisterReadDecode_1_io_iss_uop_pc_lob),
    .io_iss_uop_taken(RegisterReadDecode_1_io_iss_uop_taken),
    .io_iss_uop_imm_packed(RegisterReadDecode_1_io_iss_uop_imm_packed),
    .io_iss_uop_csr_addr(RegisterReadDecode_1_io_iss_uop_csr_addr),
    .io_iss_uop_rob_idx(RegisterReadDecode_1_io_iss_uop_rob_idx),
    .io_iss_uop_ldq_idx(RegisterReadDecode_1_io_iss_uop_ldq_idx),
    .io_iss_uop_stq_idx(RegisterReadDecode_1_io_iss_uop_stq_idx),
    .io_iss_uop_rxq_idx(RegisterReadDecode_1_io_iss_uop_rxq_idx),
    .io_iss_uop_pdst(RegisterReadDecode_1_io_iss_uop_pdst),
    .io_iss_uop_prs1(RegisterReadDecode_1_io_iss_uop_prs1),
    .io_iss_uop_prs2(RegisterReadDecode_1_io_iss_uop_prs2),
    .io_iss_uop_prs3(RegisterReadDecode_1_io_iss_uop_prs3),
    .io_iss_uop_ppred(RegisterReadDecode_1_io_iss_uop_ppred),
    .io_iss_uop_prs1_busy(RegisterReadDecode_1_io_iss_uop_prs1_busy),
    .io_iss_uop_prs2_busy(RegisterReadDecode_1_io_iss_uop_prs2_busy),
    .io_iss_uop_prs3_busy(RegisterReadDecode_1_io_iss_uop_prs3_busy),
    .io_iss_uop_ppred_busy(RegisterReadDecode_1_io_iss_uop_ppred_busy),
    .io_iss_uop_stale_pdst(RegisterReadDecode_1_io_iss_uop_stale_pdst),
    .io_iss_uop_exception(RegisterReadDecode_1_io_iss_uop_exception),
    .io_iss_uop_exc_cause(RegisterReadDecode_1_io_iss_uop_exc_cause),
    .io_iss_uop_bypassable(RegisterReadDecode_1_io_iss_uop_bypassable),
    .io_iss_uop_mem_cmd(RegisterReadDecode_1_io_iss_uop_mem_cmd),
    .io_iss_uop_mem_size(RegisterReadDecode_1_io_iss_uop_mem_size),
    .io_iss_uop_mem_signed(RegisterReadDecode_1_io_iss_uop_mem_signed),
    .io_iss_uop_is_fence(RegisterReadDecode_1_io_iss_uop_is_fence),
    .io_iss_uop_is_fencei(RegisterReadDecode_1_io_iss_uop_is_fencei),
    .io_iss_uop_is_amo(RegisterReadDecode_1_io_iss_uop_is_amo),
    .io_iss_uop_uses_ldq(RegisterReadDecode_1_io_iss_uop_uses_ldq),
    .io_iss_uop_uses_stq(RegisterReadDecode_1_io_iss_uop_uses_stq),
    .io_iss_uop_is_sys_pc2epc(RegisterReadDecode_1_io_iss_uop_is_sys_pc2epc),
    .io_iss_uop_is_unique(RegisterReadDecode_1_io_iss_uop_is_unique),
    .io_iss_uop_flush_on_commit(RegisterReadDecode_1_io_iss_uop_flush_on_commit),
    .io_iss_uop_ldst_is_rs1(RegisterReadDecode_1_io_iss_uop_ldst_is_rs1),
    .io_iss_uop_ldst(RegisterReadDecode_1_io_iss_uop_ldst),
    .io_iss_uop_lrs1(RegisterReadDecode_1_io_iss_uop_lrs1),
    .io_iss_uop_lrs2(RegisterReadDecode_1_io_iss_uop_lrs2),
    .io_iss_uop_lrs3(RegisterReadDecode_1_io_iss_uop_lrs3),
    .io_iss_uop_ldst_val(RegisterReadDecode_1_io_iss_uop_ldst_val),
    .io_iss_uop_dst_rtype(RegisterReadDecode_1_io_iss_uop_dst_rtype),
    .io_iss_uop_lrs1_rtype(RegisterReadDecode_1_io_iss_uop_lrs1_rtype),
    .io_iss_uop_lrs2_rtype(RegisterReadDecode_1_io_iss_uop_lrs2_rtype),
    .io_iss_uop_frs3_en(RegisterReadDecode_1_io_iss_uop_frs3_en),
    .io_iss_uop_fp_val(RegisterReadDecode_1_io_iss_uop_fp_val),
    .io_iss_uop_fp_single(RegisterReadDecode_1_io_iss_uop_fp_single),
    .io_iss_uop_xcpt_pf_if(RegisterReadDecode_1_io_iss_uop_xcpt_pf_if),
    .io_iss_uop_xcpt_ae_if(RegisterReadDecode_1_io_iss_uop_xcpt_ae_if),
    .io_iss_uop_xcpt_ma_if(RegisterReadDecode_1_io_iss_uop_xcpt_ma_if),
    .io_iss_uop_bp_debug_if(RegisterReadDecode_1_io_iss_uop_bp_debug_if),
    .io_iss_uop_bp_xcpt_if(RegisterReadDecode_1_io_iss_uop_bp_xcpt_if),
    .io_iss_uop_debug_fsrc(RegisterReadDecode_1_io_iss_uop_debug_fsrc),
    .io_iss_uop_debug_tsrc(RegisterReadDecode_1_io_iss_uop_debug_tsrc),
    .io_rrd_valid(RegisterReadDecode_1_io_rrd_valid),
    .io_rrd_uop_switch(RegisterReadDecode_1_io_rrd_uop_switch),
    .io_rrd_uop_switch_off(RegisterReadDecode_1_io_rrd_uop_switch_off),
    .io_rrd_uop_is_unicore(RegisterReadDecode_1_io_rrd_uop_is_unicore),
    .io_rrd_uop_shift(RegisterReadDecode_1_io_rrd_uop_shift),
    .io_rrd_uop_lrs3_rtype(RegisterReadDecode_1_io_rrd_uop_lrs3_rtype),
    .io_rrd_uop_rflag(RegisterReadDecode_1_io_rrd_uop_rflag),
    .io_rrd_uop_wflag(RegisterReadDecode_1_io_rrd_uop_wflag),
    .io_rrd_uop_prflag(RegisterReadDecode_1_io_rrd_uop_prflag),
    .io_rrd_uop_pwflag(RegisterReadDecode_1_io_rrd_uop_pwflag),
    .io_rrd_uop_pflag_busy(RegisterReadDecode_1_io_rrd_uop_pflag_busy),
    .io_rrd_uop_stale_pflag(RegisterReadDecode_1_io_rrd_uop_stale_pflag),
    .io_rrd_uop_op1_sel(RegisterReadDecode_1_io_rrd_uop_op1_sel),
    .io_rrd_uop_op2_sel(RegisterReadDecode_1_io_rrd_uop_op2_sel),
    .io_rrd_uop_split_num(RegisterReadDecode_1_io_rrd_uop_split_num),
    .io_rrd_uop_self_index(RegisterReadDecode_1_io_rrd_uop_self_index),
    .io_rrd_uop_rob_inst_idx(RegisterReadDecode_1_io_rrd_uop_rob_inst_idx),
    .io_rrd_uop_address_num(RegisterReadDecode_1_io_rrd_uop_address_num),
    .io_rrd_uop_uopc(RegisterReadDecode_1_io_rrd_uop_uopc),
    .io_rrd_uop_inst(RegisterReadDecode_1_io_rrd_uop_inst),
    .io_rrd_uop_debug_inst(RegisterReadDecode_1_io_rrd_uop_debug_inst),
    .io_rrd_uop_is_rvc(RegisterReadDecode_1_io_rrd_uop_is_rvc),
    .io_rrd_uop_debug_pc(RegisterReadDecode_1_io_rrd_uop_debug_pc),
    .io_rrd_uop_iq_type(RegisterReadDecode_1_io_rrd_uop_iq_type),
    .io_rrd_uop_fu_code(RegisterReadDecode_1_io_rrd_uop_fu_code),
    .io_rrd_uop_ctrl_br_type(RegisterReadDecode_1_io_rrd_uop_ctrl_br_type),
    .io_rrd_uop_ctrl_op1_sel(RegisterReadDecode_1_io_rrd_uop_ctrl_op1_sel),
    .io_rrd_uop_ctrl_op2_sel(RegisterReadDecode_1_io_rrd_uop_ctrl_op2_sel),
    .io_rrd_uop_ctrl_imm_sel(RegisterReadDecode_1_io_rrd_uop_ctrl_imm_sel),
    .io_rrd_uop_ctrl_op_fcn(RegisterReadDecode_1_io_rrd_uop_ctrl_op_fcn),
    .io_rrd_uop_ctrl_fcn_dw(RegisterReadDecode_1_io_rrd_uop_ctrl_fcn_dw),
    .io_rrd_uop_ctrl_csr_cmd(RegisterReadDecode_1_io_rrd_uop_ctrl_csr_cmd),
    .io_rrd_uop_ctrl_is_load(RegisterReadDecode_1_io_rrd_uop_ctrl_is_load),
    .io_rrd_uop_ctrl_is_sta(RegisterReadDecode_1_io_rrd_uop_ctrl_is_sta),
    .io_rrd_uop_ctrl_is_std(RegisterReadDecode_1_io_rrd_uop_ctrl_is_std),
    .io_rrd_uop_ctrl_op3_sel(RegisterReadDecode_1_io_rrd_uop_ctrl_op3_sel),
    .io_rrd_uop_iw_state(RegisterReadDecode_1_io_rrd_uop_iw_state),
    .io_rrd_uop_iw_p1_poisoned(RegisterReadDecode_1_io_rrd_uop_iw_p1_poisoned),
    .io_rrd_uop_iw_p2_poisoned(RegisterReadDecode_1_io_rrd_uop_iw_p2_poisoned),
    .io_rrd_uop_is_br(RegisterReadDecode_1_io_rrd_uop_is_br),
    .io_rrd_uop_is_jalr(RegisterReadDecode_1_io_rrd_uop_is_jalr),
    .io_rrd_uop_is_jal(RegisterReadDecode_1_io_rrd_uop_is_jal),
    .io_rrd_uop_is_sfb(RegisterReadDecode_1_io_rrd_uop_is_sfb),
    .io_rrd_uop_br_mask(RegisterReadDecode_1_io_rrd_uop_br_mask),
    .io_rrd_uop_br_tag(RegisterReadDecode_1_io_rrd_uop_br_tag),
    .io_rrd_uop_ftq_idx(RegisterReadDecode_1_io_rrd_uop_ftq_idx),
    .io_rrd_uop_edge_inst(RegisterReadDecode_1_io_rrd_uop_edge_inst),
    .io_rrd_uop_pc_lob(RegisterReadDecode_1_io_rrd_uop_pc_lob),
    .io_rrd_uop_taken(RegisterReadDecode_1_io_rrd_uop_taken),
    .io_rrd_uop_imm_packed(RegisterReadDecode_1_io_rrd_uop_imm_packed),
    .io_rrd_uop_csr_addr(RegisterReadDecode_1_io_rrd_uop_csr_addr),
    .io_rrd_uop_rob_idx(RegisterReadDecode_1_io_rrd_uop_rob_idx),
    .io_rrd_uop_ldq_idx(RegisterReadDecode_1_io_rrd_uop_ldq_idx),
    .io_rrd_uop_stq_idx(RegisterReadDecode_1_io_rrd_uop_stq_idx),
    .io_rrd_uop_rxq_idx(RegisterReadDecode_1_io_rrd_uop_rxq_idx),
    .io_rrd_uop_pdst(RegisterReadDecode_1_io_rrd_uop_pdst),
    .io_rrd_uop_prs1(RegisterReadDecode_1_io_rrd_uop_prs1),
    .io_rrd_uop_prs2(RegisterReadDecode_1_io_rrd_uop_prs2),
    .io_rrd_uop_prs3(RegisterReadDecode_1_io_rrd_uop_prs3),
    .io_rrd_uop_ppred(RegisterReadDecode_1_io_rrd_uop_ppred),
    .io_rrd_uop_prs1_busy(RegisterReadDecode_1_io_rrd_uop_prs1_busy),
    .io_rrd_uop_prs2_busy(RegisterReadDecode_1_io_rrd_uop_prs2_busy),
    .io_rrd_uop_prs3_busy(RegisterReadDecode_1_io_rrd_uop_prs3_busy),
    .io_rrd_uop_ppred_busy(RegisterReadDecode_1_io_rrd_uop_ppred_busy),
    .io_rrd_uop_stale_pdst(RegisterReadDecode_1_io_rrd_uop_stale_pdst),
    .io_rrd_uop_exception(RegisterReadDecode_1_io_rrd_uop_exception),
    .io_rrd_uop_exc_cause(RegisterReadDecode_1_io_rrd_uop_exc_cause),
    .io_rrd_uop_bypassable(RegisterReadDecode_1_io_rrd_uop_bypassable),
    .io_rrd_uop_mem_cmd(RegisterReadDecode_1_io_rrd_uop_mem_cmd),
    .io_rrd_uop_mem_size(RegisterReadDecode_1_io_rrd_uop_mem_size),
    .io_rrd_uop_mem_signed(RegisterReadDecode_1_io_rrd_uop_mem_signed),
    .io_rrd_uop_is_fence(RegisterReadDecode_1_io_rrd_uop_is_fence),
    .io_rrd_uop_is_fencei(RegisterReadDecode_1_io_rrd_uop_is_fencei),
    .io_rrd_uop_is_amo(RegisterReadDecode_1_io_rrd_uop_is_amo),
    .io_rrd_uop_uses_ldq(RegisterReadDecode_1_io_rrd_uop_uses_ldq),
    .io_rrd_uop_uses_stq(RegisterReadDecode_1_io_rrd_uop_uses_stq),
    .io_rrd_uop_is_sys_pc2epc(RegisterReadDecode_1_io_rrd_uop_is_sys_pc2epc),
    .io_rrd_uop_is_unique(RegisterReadDecode_1_io_rrd_uop_is_unique),
    .io_rrd_uop_flush_on_commit(RegisterReadDecode_1_io_rrd_uop_flush_on_commit),
    .io_rrd_uop_ldst_is_rs1(RegisterReadDecode_1_io_rrd_uop_ldst_is_rs1),
    .io_rrd_uop_ldst(RegisterReadDecode_1_io_rrd_uop_ldst),
    .io_rrd_uop_lrs1(RegisterReadDecode_1_io_rrd_uop_lrs1),
    .io_rrd_uop_lrs2(RegisterReadDecode_1_io_rrd_uop_lrs2),
    .io_rrd_uop_lrs3(RegisterReadDecode_1_io_rrd_uop_lrs3),
    .io_rrd_uop_ldst_val(RegisterReadDecode_1_io_rrd_uop_ldst_val),
    .io_rrd_uop_dst_rtype(RegisterReadDecode_1_io_rrd_uop_dst_rtype),
    .io_rrd_uop_lrs1_rtype(RegisterReadDecode_1_io_rrd_uop_lrs1_rtype),
    .io_rrd_uop_lrs2_rtype(RegisterReadDecode_1_io_rrd_uop_lrs2_rtype),
    .io_rrd_uop_frs3_en(RegisterReadDecode_1_io_rrd_uop_frs3_en),
    .io_rrd_uop_fp_val(RegisterReadDecode_1_io_rrd_uop_fp_val),
    .io_rrd_uop_fp_single(RegisterReadDecode_1_io_rrd_uop_fp_single),
    .io_rrd_uop_xcpt_pf_if(RegisterReadDecode_1_io_rrd_uop_xcpt_pf_if),
    .io_rrd_uop_xcpt_ae_if(RegisterReadDecode_1_io_rrd_uop_xcpt_ae_if),
    .io_rrd_uop_xcpt_ma_if(RegisterReadDecode_1_io_rrd_uop_xcpt_ma_if),
    .io_rrd_uop_bp_debug_if(RegisterReadDecode_1_io_rrd_uop_bp_debug_if),
    .io_rrd_uop_bp_xcpt_if(RegisterReadDecode_1_io_rrd_uop_bp_xcpt_if),
    .io_rrd_uop_debug_fsrc(RegisterReadDecode_1_io_rrd_uop_debug_fsrc),
    .io_rrd_uop_debug_tsrc(RegisterReadDecode_1_io_rrd_uop_debug_tsrc)
  );
  RegisterReadDecode_3 RegisterReadDecode_2 ( // @[register-read.scala 86:33]
    .clock(RegisterReadDecode_2_clock),
    .reset(RegisterReadDecode_2_reset),
    .io_iss_valid(RegisterReadDecode_2_io_iss_valid),
    .io_iss_uop_switch(RegisterReadDecode_2_io_iss_uop_switch),
    .io_iss_uop_switch_off(RegisterReadDecode_2_io_iss_uop_switch_off),
    .io_iss_uop_is_unicore(RegisterReadDecode_2_io_iss_uop_is_unicore),
    .io_iss_uop_shift(RegisterReadDecode_2_io_iss_uop_shift),
    .io_iss_uop_lrs3_rtype(RegisterReadDecode_2_io_iss_uop_lrs3_rtype),
    .io_iss_uop_rflag(RegisterReadDecode_2_io_iss_uop_rflag),
    .io_iss_uop_wflag(RegisterReadDecode_2_io_iss_uop_wflag),
    .io_iss_uop_prflag(RegisterReadDecode_2_io_iss_uop_prflag),
    .io_iss_uop_pwflag(RegisterReadDecode_2_io_iss_uop_pwflag),
    .io_iss_uop_pflag_busy(RegisterReadDecode_2_io_iss_uop_pflag_busy),
    .io_iss_uop_stale_pflag(RegisterReadDecode_2_io_iss_uop_stale_pflag),
    .io_iss_uop_op1_sel(RegisterReadDecode_2_io_iss_uop_op1_sel),
    .io_iss_uop_op2_sel(RegisterReadDecode_2_io_iss_uop_op2_sel),
    .io_iss_uop_split_num(RegisterReadDecode_2_io_iss_uop_split_num),
    .io_iss_uop_self_index(RegisterReadDecode_2_io_iss_uop_self_index),
    .io_iss_uop_rob_inst_idx(RegisterReadDecode_2_io_iss_uop_rob_inst_idx),
    .io_iss_uop_address_num(RegisterReadDecode_2_io_iss_uop_address_num),
    .io_iss_uop_uopc(RegisterReadDecode_2_io_iss_uop_uopc),
    .io_iss_uop_inst(RegisterReadDecode_2_io_iss_uop_inst),
    .io_iss_uop_debug_inst(RegisterReadDecode_2_io_iss_uop_debug_inst),
    .io_iss_uop_is_rvc(RegisterReadDecode_2_io_iss_uop_is_rvc),
    .io_iss_uop_debug_pc(RegisterReadDecode_2_io_iss_uop_debug_pc),
    .io_iss_uop_iq_type(RegisterReadDecode_2_io_iss_uop_iq_type),
    .io_iss_uop_fu_code(RegisterReadDecode_2_io_iss_uop_fu_code),
    .io_iss_uop_ctrl_br_type(RegisterReadDecode_2_io_iss_uop_ctrl_br_type),
    .io_iss_uop_ctrl_op1_sel(RegisterReadDecode_2_io_iss_uop_ctrl_op1_sel),
    .io_iss_uop_ctrl_op2_sel(RegisterReadDecode_2_io_iss_uop_ctrl_op2_sel),
    .io_iss_uop_ctrl_imm_sel(RegisterReadDecode_2_io_iss_uop_ctrl_imm_sel),
    .io_iss_uop_ctrl_op_fcn(RegisterReadDecode_2_io_iss_uop_ctrl_op_fcn),
    .io_iss_uop_ctrl_fcn_dw(RegisterReadDecode_2_io_iss_uop_ctrl_fcn_dw),
    .io_iss_uop_ctrl_csr_cmd(RegisterReadDecode_2_io_iss_uop_ctrl_csr_cmd),
    .io_iss_uop_ctrl_is_load(RegisterReadDecode_2_io_iss_uop_ctrl_is_load),
    .io_iss_uop_ctrl_is_sta(RegisterReadDecode_2_io_iss_uop_ctrl_is_sta),
    .io_iss_uop_ctrl_is_std(RegisterReadDecode_2_io_iss_uop_ctrl_is_std),
    .io_iss_uop_ctrl_op3_sel(RegisterReadDecode_2_io_iss_uop_ctrl_op3_sel),
    .io_iss_uop_iw_state(RegisterReadDecode_2_io_iss_uop_iw_state),
    .io_iss_uop_iw_p1_poisoned(RegisterReadDecode_2_io_iss_uop_iw_p1_poisoned),
    .io_iss_uop_iw_p2_poisoned(RegisterReadDecode_2_io_iss_uop_iw_p2_poisoned),
    .io_iss_uop_is_br(RegisterReadDecode_2_io_iss_uop_is_br),
    .io_iss_uop_is_jalr(RegisterReadDecode_2_io_iss_uop_is_jalr),
    .io_iss_uop_is_jal(RegisterReadDecode_2_io_iss_uop_is_jal),
    .io_iss_uop_is_sfb(RegisterReadDecode_2_io_iss_uop_is_sfb),
    .io_iss_uop_br_mask(RegisterReadDecode_2_io_iss_uop_br_mask),
    .io_iss_uop_br_tag(RegisterReadDecode_2_io_iss_uop_br_tag),
    .io_iss_uop_ftq_idx(RegisterReadDecode_2_io_iss_uop_ftq_idx),
    .io_iss_uop_edge_inst(RegisterReadDecode_2_io_iss_uop_edge_inst),
    .io_iss_uop_pc_lob(RegisterReadDecode_2_io_iss_uop_pc_lob),
    .io_iss_uop_taken(RegisterReadDecode_2_io_iss_uop_taken),
    .io_iss_uop_imm_packed(RegisterReadDecode_2_io_iss_uop_imm_packed),
    .io_iss_uop_csr_addr(RegisterReadDecode_2_io_iss_uop_csr_addr),
    .io_iss_uop_rob_idx(RegisterReadDecode_2_io_iss_uop_rob_idx),
    .io_iss_uop_ldq_idx(RegisterReadDecode_2_io_iss_uop_ldq_idx),
    .io_iss_uop_stq_idx(RegisterReadDecode_2_io_iss_uop_stq_idx),
    .io_iss_uop_rxq_idx(RegisterReadDecode_2_io_iss_uop_rxq_idx),
    .io_iss_uop_pdst(RegisterReadDecode_2_io_iss_uop_pdst),
    .io_iss_uop_prs1(RegisterReadDecode_2_io_iss_uop_prs1),
    .io_iss_uop_prs2(RegisterReadDecode_2_io_iss_uop_prs2),
    .io_iss_uop_prs3(RegisterReadDecode_2_io_iss_uop_prs3),
    .io_iss_uop_ppred(RegisterReadDecode_2_io_iss_uop_ppred),
    .io_iss_uop_prs1_busy(RegisterReadDecode_2_io_iss_uop_prs1_busy),
    .io_iss_uop_prs2_busy(RegisterReadDecode_2_io_iss_uop_prs2_busy),
    .io_iss_uop_prs3_busy(RegisterReadDecode_2_io_iss_uop_prs3_busy),
    .io_iss_uop_ppred_busy(RegisterReadDecode_2_io_iss_uop_ppred_busy),
    .io_iss_uop_stale_pdst(RegisterReadDecode_2_io_iss_uop_stale_pdst),
    .io_iss_uop_exception(RegisterReadDecode_2_io_iss_uop_exception),
    .io_iss_uop_exc_cause(RegisterReadDecode_2_io_iss_uop_exc_cause),
    .io_iss_uop_bypassable(RegisterReadDecode_2_io_iss_uop_bypassable),
    .io_iss_uop_mem_cmd(RegisterReadDecode_2_io_iss_uop_mem_cmd),
    .io_iss_uop_mem_size(RegisterReadDecode_2_io_iss_uop_mem_size),
    .io_iss_uop_mem_signed(RegisterReadDecode_2_io_iss_uop_mem_signed),
    .io_iss_uop_is_fence(RegisterReadDecode_2_io_iss_uop_is_fence),
    .io_iss_uop_is_fencei(RegisterReadDecode_2_io_iss_uop_is_fencei),
    .io_iss_uop_is_amo(RegisterReadDecode_2_io_iss_uop_is_amo),
    .io_iss_uop_uses_ldq(RegisterReadDecode_2_io_iss_uop_uses_ldq),
    .io_iss_uop_uses_stq(RegisterReadDecode_2_io_iss_uop_uses_stq),
    .io_iss_uop_is_sys_pc2epc(RegisterReadDecode_2_io_iss_uop_is_sys_pc2epc),
    .io_iss_uop_is_unique(RegisterReadDecode_2_io_iss_uop_is_unique),
    .io_iss_uop_flush_on_commit(RegisterReadDecode_2_io_iss_uop_flush_on_commit),
    .io_iss_uop_ldst_is_rs1(RegisterReadDecode_2_io_iss_uop_ldst_is_rs1),
    .io_iss_uop_ldst(RegisterReadDecode_2_io_iss_uop_ldst),
    .io_iss_uop_lrs1(RegisterReadDecode_2_io_iss_uop_lrs1),
    .io_iss_uop_lrs2(RegisterReadDecode_2_io_iss_uop_lrs2),
    .io_iss_uop_lrs3(RegisterReadDecode_2_io_iss_uop_lrs3),
    .io_iss_uop_ldst_val(RegisterReadDecode_2_io_iss_uop_ldst_val),
    .io_iss_uop_dst_rtype(RegisterReadDecode_2_io_iss_uop_dst_rtype),
    .io_iss_uop_lrs1_rtype(RegisterReadDecode_2_io_iss_uop_lrs1_rtype),
    .io_iss_uop_lrs2_rtype(RegisterReadDecode_2_io_iss_uop_lrs2_rtype),
    .io_iss_uop_frs3_en(RegisterReadDecode_2_io_iss_uop_frs3_en),
    .io_iss_uop_fp_val(RegisterReadDecode_2_io_iss_uop_fp_val),
    .io_iss_uop_fp_single(RegisterReadDecode_2_io_iss_uop_fp_single),
    .io_iss_uop_xcpt_pf_if(RegisterReadDecode_2_io_iss_uop_xcpt_pf_if),
    .io_iss_uop_xcpt_ae_if(RegisterReadDecode_2_io_iss_uop_xcpt_ae_if),
    .io_iss_uop_xcpt_ma_if(RegisterReadDecode_2_io_iss_uop_xcpt_ma_if),
    .io_iss_uop_bp_debug_if(RegisterReadDecode_2_io_iss_uop_bp_debug_if),
    .io_iss_uop_bp_xcpt_if(RegisterReadDecode_2_io_iss_uop_bp_xcpt_if),
    .io_iss_uop_debug_fsrc(RegisterReadDecode_2_io_iss_uop_debug_fsrc),
    .io_iss_uop_debug_tsrc(RegisterReadDecode_2_io_iss_uop_debug_tsrc),
    .io_rrd_valid(RegisterReadDecode_2_io_rrd_valid),
    .io_rrd_uop_switch(RegisterReadDecode_2_io_rrd_uop_switch),
    .io_rrd_uop_switch_off(RegisterReadDecode_2_io_rrd_uop_switch_off),
    .io_rrd_uop_is_unicore(RegisterReadDecode_2_io_rrd_uop_is_unicore),
    .io_rrd_uop_shift(RegisterReadDecode_2_io_rrd_uop_shift),
    .io_rrd_uop_lrs3_rtype(RegisterReadDecode_2_io_rrd_uop_lrs3_rtype),
    .io_rrd_uop_rflag(RegisterReadDecode_2_io_rrd_uop_rflag),
    .io_rrd_uop_wflag(RegisterReadDecode_2_io_rrd_uop_wflag),
    .io_rrd_uop_prflag(RegisterReadDecode_2_io_rrd_uop_prflag),
    .io_rrd_uop_pwflag(RegisterReadDecode_2_io_rrd_uop_pwflag),
    .io_rrd_uop_pflag_busy(RegisterReadDecode_2_io_rrd_uop_pflag_busy),
    .io_rrd_uop_stale_pflag(RegisterReadDecode_2_io_rrd_uop_stale_pflag),
    .io_rrd_uop_op1_sel(RegisterReadDecode_2_io_rrd_uop_op1_sel),
    .io_rrd_uop_op2_sel(RegisterReadDecode_2_io_rrd_uop_op2_sel),
    .io_rrd_uop_split_num(RegisterReadDecode_2_io_rrd_uop_split_num),
    .io_rrd_uop_self_index(RegisterReadDecode_2_io_rrd_uop_self_index),
    .io_rrd_uop_rob_inst_idx(RegisterReadDecode_2_io_rrd_uop_rob_inst_idx),
    .io_rrd_uop_address_num(RegisterReadDecode_2_io_rrd_uop_address_num),
    .io_rrd_uop_uopc(RegisterReadDecode_2_io_rrd_uop_uopc),
    .io_rrd_uop_inst(RegisterReadDecode_2_io_rrd_uop_inst),
    .io_rrd_uop_debug_inst(RegisterReadDecode_2_io_rrd_uop_debug_inst),
    .io_rrd_uop_is_rvc(RegisterReadDecode_2_io_rrd_uop_is_rvc),
    .io_rrd_uop_debug_pc(RegisterReadDecode_2_io_rrd_uop_debug_pc),
    .io_rrd_uop_iq_type(RegisterReadDecode_2_io_rrd_uop_iq_type),
    .io_rrd_uop_fu_code(RegisterReadDecode_2_io_rrd_uop_fu_code),
    .io_rrd_uop_ctrl_br_type(RegisterReadDecode_2_io_rrd_uop_ctrl_br_type),
    .io_rrd_uop_ctrl_op1_sel(RegisterReadDecode_2_io_rrd_uop_ctrl_op1_sel),
    .io_rrd_uop_ctrl_op2_sel(RegisterReadDecode_2_io_rrd_uop_ctrl_op2_sel),
    .io_rrd_uop_ctrl_imm_sel(RegisterReadDecode_2_io_rrd_uop_ctrl_imm_sel),
    .io_rrd_uop_ctrl_op_fcn(RegisterReadDecode_2_io_rrd_uop_ctrl_op_fcn),
    .io_rrd_uop_ctrl_fcn_dw(RegisterReadDecode_2_io_rrd_uop_ctrl_fcn_dw),
    .io_rrd_uop_ctrl_csr_cmd(RegisterReadDecode_2_io_rrd_uop_ctrl_csr_cmd),
    .io_rrd_uop_ctrl_is_load(RegisterReadDecode_2_io_rrd_uop_ctrl_is_load),
    .io_rrd_uop_ctrl_is_sta(RegisterReadDecode_2_io_rrd_uop_ctrl_is_sta),
    .io_rrd_uop_ctrl_is_std(RegisterReadDecode_2_io_rrd_uop_ctrl_is_std),
    .io_rrd_uop_ctrl_op3_sel(RegisterReadDecode_2_io_rrd_uop_ctrl_op3_sel),
    .io_rrd_uop_iw_state(RegisterReadDecode_2_io_rrd_uop_iw_state),
    .io_rrd_uop_iw_p1_poisoned(RegisterReadDecode_2_io_rrd_uop_iw_p1_poisoned),
    .io_rrd_uop_iw_p2_poisoned(RegisterReadDecode_2_io_rrd_uop_iw_p2_poisoned),
    .io_rrd_uop_is_br(RegisterReadDecode_2_io_rrd_uop_is_br),
    .io_rrd_uop_is_jalr(RegisterReadDecode_2_io_rrd_uop_is_jalr),
    .io_rrd_uop_is_jal(RegisterReadDecode_2_io_rrd_uop_is_jal),
    .io_rrd_uop_is_sfb(RegisterReadDecode_2_io_rrd_uop_is_sfb),
    .io_rrd_uop_br_mask(RegisterReadDecode_2_io_rrd_uop_br_mask),
    .io_rrd_uop_br_tag(RegisterReadDecode_2_io_rrd_uop_br_tag),
    .io_rrd_uop_ftq_idx(RegisterReadDecode_2_io_rrd_uop_ftq_idx),
    .io_rrd_uop_edge_inst(RegisterReadDecode_2_io_rrd_uop_edge_inst),
    .io_rrd_uop_pc_lob(RegisterReadDecode_2_io_rrd_uop_pc_lob),
    .io_rrd_uop_taken(RegisterReadDecode_2_io_rrd_uop_taken),
    .io_rrd_uop_imm_packed(RegisterReadDecode_2_io_rrd_uop_imm_packed),
    .io_rrd_uop_csr_addr(RegisterReadDecode_2_io_rrd_uop_csr_addr),
    .io_rrd_uop_rob_idx(RegisterReadDecode_2_io_rrd_uop_rob_idx),
    .io_rrd_uop_ldq_idx(RegisterReadDecode_2_io_rrd_uop_ldq_idx),
    .io_rrd_uop_stq_idx(RegisterReadDecode_2_io_rrd_uop_stq_idx),
    .io_rrd_uop_rxq_idx(RegisterReadDecode_2_io_rrd_uop_rxq_idx),
    .io_rrd_uop_pdst(RegisterReadDecode_2_io_rrd_uop_pdst),
    .io_rrd_uop_prs1(RegisterReadDecode_2_io_rrd_uop_prs1),
    .io_rrd_uop_prs2(RegisterReadDecode_2_io_rrd_uop_prs2),
    .io_rrd_uop_prs3(RegisterReadDecode_2_io_rrd_uop_prs3),
    .io_rrd_uop_ppred(RegisterReadDecode_2_io_rrd_uop_ppred),
    .io_rrd_uop_prs1_busy(RegisterReadDecode_2_io_rrd_uop_prs1_busy),
    .io_rrd_uop_prs2_busy(RegisterReadDecode_2_io_rrd_uop_prs2_busy),
    .io_rrd_uop_prs3_busy(RegisterReadDecode_2_io_rrd_uop_prs3_busy),
    .io_rrd_uop_ppred_busy(RegisterReadDecode_2_io_rrd_uop_ppred_busy),
    .io_rrd_uop_stale_pdst(RegisterReadDecode_2_io_rrd_uop_stale_pdst),
    .io_rrd_uop_exception(RegisterReadDecode_2_io_rrd_uop_exception),
    .io_rrd_uop_exc_cause(RegisterReadDecode_2_io_rrd_uop_exc_cause),
    .io_rrd_uop_bypassable(RegisterReadDecode_2_io_rrd_uop_bypassable),
    .io_rrd_uop_mem_cmd(RegisterReadDecode_2_io_rrd_uop_mem_cmd),
    .io_rrd_uop_mem_size(RegisterReadDecode_2_io_rrd_uop_mem_size),
    .io_rrd_uop_mem_signed(RegisterReadDecode_2_io_rrd_uop_mem_signed),
    .io_rrd_uop_is_fence(RegisterReadDecode_2_io_rrd_uop_is_fence),
    .io_rrd_uop_is_fencei(RegisterReadDecode_2_io_rrd_uop_is_fencei),
    .io_rrd_uop_is_amo(RegisterReadDecode_2_io_rrd_uop_is_amo),
    .io_rrd_uop_uses_ldq(RegisterReadDecode_2_io_rrd_uop_uses_ldq),
    .io_rrd_uop_uses_stq(RegisterReadDecode_2_io_rrd_uop_uses_stq),
    .io_rrd_uop_is_sys_pc2epc(RegisterReadDecode_2_io_rrd_uop_is_sys_pc2epc),
    .io_rrd_uop_is_unique(RegisterReadDecode_2_io_rrd_uop_is_unique),
    .io_rrd_uop_flush_on_commit(RegisterReadDecode_2_io_rrd_uop_flush_on_commit),
    .io_rrd_uop_ldst_is_rs1(RegisterReadDecode_2_io_rrd_uop_ldst_is_rs1),
    .io_rrd_uop_ldst(RegisterReadDecode_2_io_rrd_uop_ldst),
    .io_rrd_uop_lrs1(RegisterReadDecode_2_io_rrd_uop_lrs1),
    .io_rrd_uop_lrs2(RegisterReadDecode_2_io_rrd_uop_lrs2),
    .io_rrd_uop_lrs3(RegisterReadDecode_2_io_rrd_uop_lrs3),
    .io_rrd_uop_ldst_val(RegisterReadDecode_2_io_rrd_uop_ldst_val),
    .io_rrd_uop_dst_rtype(RegisterReadDecode_2_io_rrd_uop_dst_rtype),
    .io_rrd_uop_lrs1_rtype(RegisterReadDecode_2_io_rrd_uop_lrs1_rtype),
    .io_rrd_uop_lrs2_rtype(RegisterReadDecode_2_io_rrd_uop_lrs2_rtype),
    .io_rrd_uop_frs3_en(RegisterReadDecode_2_io_rrd_uop_frs3_en),
    .io_rrd_uop_fp_val(RegisterReadDecode_2_io_rrd_uop_fp_val),
    .io_rrd_uop_fp_single(RegisterReadDecode_2_io_rrd_uop_fp_single),
    .io_rrd_uop_xcpt_pf_if(RegisterReadDecode_2_io_rrd_uop_xcpt_pf_if),
    .io_rrd_uop_xcpt_ae_if(RegisterReadDecode_2_io_rrd_uop_xcpt_ae_if),
    .io_rrd_uop_xcpt_ma_if(RegisterReadDecode_2_io_rrd_uop_xcpt_ma_if),
    .io_rrd_uop_bp_debug_if(RegisterReadDecode_2_io_rrd_uop_bp_debug_if),
    .io_rrd_uop_bp_xcpt_if(RegisterReadDecode_2_io_rrd_uop_bp_xcpt_if),
    .io_rrd_uop_debug_fsrc(RegisterReadDecode_2_io_rrd_uop_debug_fsrc),
    .io_rrd_uop_debug_tsrc(RegisterReadDecode_2_io_rrd_uop_debug_tsrc)
  );
  assign io_rf_read_ports_0_addr = io_iss_uops_0_prs1; // @[register-read.scala 127:56]
  assign io_rf_read_ports_1_addr = io_iss_uops_0_prs2; // @[register-read.scala 128:56]
  assign io_rf_read_ports_2_addr = io_iss_uops_0_prs3; // @[register-read.scala 129:56]
  assign io_rf_read_ports_3_addr = io_iss_uops_1_prs1; // @[register-read.scala 127:56]
  assign io_rf_read_ports_4_addr = io_iss_uops_1_prs2; // @[register-read.scala 128:56]
  assign io_rf_read_ports_5_addr = io_iss_uops_1_prs3; // @[register-read.scala 129:56]
  assign io_rf_read_ports_6_addr = io_iss_uops_2_prs1; // @[register-read.scala 127:56]
  assign io_rf_read_ports_7_addr = io_iss_uops_2_prs2; // @[register-read.scala 128:56]
  assign io_rf_read_ports_8_addr = io_iss_uops_2_prs3; // @[register-read.scala 129:56]
  assign io_prf_read_ports_0_addr = 5'h0;
  assign io_prf_read_ports_1_addr = 5'h0;
  assign io_prf_read_ports_2_addr = 5'h0;
  assign io_flag_rf_read_ports_0_addr = {{3'd0}, io_iss_uops_0_prflag}; // @[register-read.scala 142:35]
  assign io_flag_rf_read_ports_1_addr = {{3'd0}, io_iss_uops_1_prflag}; // @[register-read.scala 142:35]
  assign io_flag_rf_read_ports_2_addr = {{3'd0}, io_iss_uops_2_prflag}; // @[register-read.scala 142:35]
  assign io_exe_reqs_0_valid = exe_reg_valids_0; // @[register-read.scala 254:29]
  assign io_exe_reqs_0_bits_uop_switch = exe_reg_uops_0_switch; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_switch_off = exe_reg_uops_0_switch_off; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_is_unicore = exe_reg_uops_0_is_unicore; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_shift = exe_reg_uops_0_shift; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_lrs3_rtype = exe_reg_uops_0_lrs3_rtype; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_rflag = exe_reg_uops_0_rflag; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_wflag = exe_reg_uops_0_wflag; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_prflag = exe_reg_uops_0_prflag; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_pwflag = exe_reg_uops_0_pwflag; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_pflag_busy = exe_reg_uops_0_pflag_busy; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_stale_pflag = exe_reg_uops_0_stale_pflag; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_op1_sel = exe_reg_uops_0_op1_sel; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_op2_sel = exe_reg_uops_0_op2_sel; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_split_num = exe_reg_uops_0_split_num; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_self_index = exe_reg_uops_0_self_index; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_rob_inst_idx = exe_reg_uops_0_rob_inst_idx; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_address_num = exe_reg_uops_0_address_num; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_uopc = exe_reg_uops_0_uopc; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_inst = exe_reg_uops_0_inst; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_debug_inst = exe_reg_uops_0_debug_inst; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_is_rvc = exe_reg_uops_0_is_rvc; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_debug_pc = exe_reg_uops_0_debug_pc; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_iq_type = exe_reg_uops_0_iq_type; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_fu_code = exe_reg_uops_0_fu_code; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_ctrl_br_type = exe_reg_uops_0_ctrl_br_type; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_ctrl_op1_sel = exe_reg_uops_0_ctrl_op1_sel; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_ctrl_op2_sel = exe_reg_uops_0_ctrl_op2_sel; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_ctrl_imm_sel = exe_reg_uops_0_ctrl_imm_sel; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_ctrl_op_fcn = exe_reg_uops_0_ctrl_op_fcn; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_ctrl_fcn_dw = exe_reg_uops_0_ctrl_fcn_dw; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_ctrl_csr_cmd = exe_reg_uops_0_ctrl_csr_cmd; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_ctrl_is_load = exe_reg_uops_0_ctrl_is_load; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_ctrl_is_sta = exe_reg_uops_0_ctrl_is_sta; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_ctrl_is_std = exe_reg_uops_0_ctrl_is_std; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_ctrl_op3_sel = exe_reg_uops_0_ctrl_op3_sel; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_iw_state = exe_reg_uops_0_iw_state; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_iw_p1_poisoned = exe_reg_uops_0_iw_p1_poisoned; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_iw_p2_poisoned = exe_reg_uops_0_iw_p2_poisoned; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_is_br = exe_reg_uops_0_is_br; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_is_jalr = exe_reg_uops_0_is_jalr; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_is_jal = exe_reg_uops_0_is_jal; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_is_sfb = exe_reg_uops_0_is_sfb; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_br_mask = exe_reg_uops_0_br_mask; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_br_tag = exe_reg_uops_0_br_tag; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_ftq_idx = exe_reg_uops_0_ftq_idx; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_edge_inst = exe_reg_uops_0_edge_inst; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_pc_lob = exe_reg_uops_0_pc_lob; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_taken = exe_reg_uops_0_taken; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_imm_packed = exe_reg_uops_0_imm_packed; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_csr_addr = exe_reg_uops_0_csr_addr; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_rob_idx = exe_reg_uops_0_rob_idx; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_ldq_idx = exe_reg_uops_0_ldq_idx; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_stq_idx = exe_reg_uops_0_stq_idx; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_rxq_idx = exe_reg_uops_0_rxq_idx; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_pdst = exe_reg_uops_0_pdst; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_prs1 = exe_reg_uops_0_prs1; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_prs2 = exe_reg_uops_0_prs2; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_prs3 = exe_reg_uops_0_prs3; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_ppred = exe_reg_uops_0_ppred; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_prs1_busy = exe_reg_uops_0_prs1_busy; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_prs2_busy = exe_reg_uops_0_prs2_busy; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_prs3_busy = exe_reg_uops_0_prs3_busy; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_ppred_busy = exe_reg_uops_0_ppred_busy; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_stale_pdst = exe_reg_uops_0_stale_pdst; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_exception = exe_reg_uops_0_exception; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_exc_cause = exe_reg_uops_0_exc_cause; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_bypassable = exe_reg_uops_0_bypassable; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_mem_cmd = exe_reg_uops_0_mem_cmd; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_mem_size = exe_reg_uops_0_mem_size; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_mem_signed = exe_reg_uops_0_mem_signed; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_is_fence = exe_reg_uops_0_is_fence; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_is_fencei = exe_reg_uops_0_is_fencei; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_is_amo = exe_reg_uops_0_is_amo; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_uses_ldq = exe_reg_uops_0_uses_ldq; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_uses_stq = exe_reg_uops_0_uses_stq; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_is_sys_pc2epc = exe_reg_uops_0_is_sys_pc2epc; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_is_unique = exe_reg_uops_0_is_unique; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_flush_on_commit = exe_reg_uops_0_flush_on_commit; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_ldst_is_rs1 = exe_reg_uops_0_ldst_is_rs1; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_ldst = exe_reg_uops_0_ldst; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_lrs1 = exe_reg_uops_0_lrs1; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_lrs2 = exe_reg_uops_0_lrs2; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_lrs3 = exe_reg_uops_0_lrs3; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_ldst_val = exe_reg_uops_0_ldst_val; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_dst_rtype = exe_reg_uops_0_dst_rtype; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_lrs1_rtype = exe_reg_uops_0_lrs1_rtype; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_lrs2_rtype = exe_reg_uops_0_lrs2_rtype; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_frs3_en = exe_reg_uops_0_frs3_en; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_fp_val = exe_reg_uops_0_fp_val; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_fp_single = exe_reg_uops_0_fp_single; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_xcpt_pf_if = exe_reg_uops_0_xcpt_pf_if; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_xcpt_ae_if = exe_reg_uops_0_xcpt_ae_if; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_xcpt_ma_if = exe_reg_uops_0_xcpt_ma_if; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_bp_debug_if = exe_reg_uops_0_bp_debug_if; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_bp_xcpt_if = exe_reg_uops_0_bp_xcpt_if; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_debug_fsrc = exe_reg_uops_0_debug_fsrc; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_uop_debug_tsrc = exe_reg_uops_0_debug_tsrc; // @[register-read.scala 255:29]
  assign io_exe_reqs_0_bits_rs1_data = exe_reg_rs1_data_0; // @[register-read.scala 256:56]
  assign io_exe_reqs_0_bits_rs2_data = exe_reg_rs2_data_0; // @[register-read.scala 257:56]
  assign io_exe_reqs_0_bits_rs3_data = exe_reg_rs3_data_0; // @[register-read.scala 258:56]
  assign io_exe_reqs_0_bits_pred_data = 1'h0;
  assign io_exe_reqs_0_bits_flagdata = exe_reg_flag_data_0; // @[register-read.scala 261:34]
  assign io_exe_reqs_0_bits_fflagdata = 32'h0;
  assign io_exe_reqs_0_bits_kill = 1'h0;
  assign io_exe_reqs_1_valid = exe_reg_valids_1; // @[register-read.scala 254:29]
  assign io_exe_reqs_1_bits_uop_switch = exe_reg_uops_1_switch; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_switch_off = exe_reg_uops_1_switch_off; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_is_unicore = exe_reg_uops_1_is_unicore; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_shift = exe_reg_uops_1_shift; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_lrs3_rtype = exe_reg_uops_1_lrs3_rtype; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_rflag = exe_reg_uops_1_rflag; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_wflag = exe_reg_uops_1_wflag; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_prflag = exe_reg_uops_1_prflag; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_pwflag = exe_reg_uops_1_pwflag; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_pflag_busy = exe_reg_uops_1_pflag_busy; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_stale_pflag = exe_reg_uops_1_stale_pflag; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_op1_sel = exe_reg_uops_1_op1_sel; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_op2_sel = exe_reg_uops_1_op2_sel; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_split_num = exe_reg_uops_1_split_num; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_self_index = exe_reg_uops_1_self_index; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_rob_inst_idx = exe_reg_uops_1_rob_inst_idx; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_address_num = exe_reg_uops_1_address_num; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_uopc = exe_reg_uops_1_uopc; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_inst = exe_reg_uops_1_inst; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_debug_inst = exe_reg_uops_1_debug_inst; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_is_rvc = exe_reg_uops_1_is_rvc; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_debug_pc = exe_reg_uops_1_debug_pc; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_iq_type = exe_reg_uops_1_iq_type; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_fu_code = exe_reg_uops_1_fu_code; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_ctrl_br_type = exe_reg_uops_1_ctrl_br_type; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_ctrl_op1_sel = exe_reg_uops_1_ctrl_op1_sel; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_ctrl_op2_sel = exe_reg_uops_1_ctrl_op2_sel; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_ctrl_imm_sel = exe_reg_uops_1_ctrl_imm_sel; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_ctrl_op_fcn = exe_reg_uops_1_ctrl_op_fcn; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_ctrl_fcn_dw = exe_reg_uops_1_ctrl_fcn_dw; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_ctrl_csr_cmd = exe_reg_uops_1_ctrl_csr_cmd; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_ctrl_is_load = exe_reg_uops_1_ctrl_is_load; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_ctrl_is_sta = exe_reg_uops_1_ctrl_is_sta; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_ctrl_is_std = exe_reg_uops_1_ctrl_is_std; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_ctrl_op3_sel = exe_reg_uops_1_ctrl_op3_sel; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_iw_state = exe_reg_uops_1_iw_state; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_iw_p1_poisoned = exe_reg_uops_1_iw_p1_poisoned; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_iw_p2_poisoned = exe_reg_uops_1_iw_p2_poisoned; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_is_br = exe_reg_uops_1_is_br; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_is_jalr = exe_reg_uops_1_is_jalr; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_is_jal = exe_reg_uops_1_is_jal; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_is_sfb = exe_reg_uops_1_is_sfb; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_br_mask = exe_reg_uops_1_br_mask; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_br_tag = exe_reg_uops_1_br_tag; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_ftq_idx = exe_reg_uops_1_ftq_idx; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_edge_inst = exe_reg_uops_1_edge_inst; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_pc_lob = exe_reg_uops_1_pc_lob; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_taken = exe_reg_uops_1_taken; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_imm_packed = exe_reg_uops_1_imm_packed; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_csr_addr = exe_reg_uops_1_csr_addr; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_rob_idx = exe_reg_uops_1_rob_idx; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_ldq_idx = exe_reg_uops_1_ldq_idx; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_stq_idx = exe_reg_uops_1_stq_idx; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_rxq_idx = exe_reg_uops_1_rxq_idx; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_pdst = exe_reg_uops_1_pdst; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_prs1 = exe_reg_uops_1_prs1; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_prs2 = exe_reg_uops_1_prs2; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_prs3 = exe_reg_uops_1_prs3; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_ppred = exe_reg_uops_1_ppred; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_prs1_busy = exe_reg_uops_1_prs1_busy; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_prs2_busy = exe_reg_uops_1_prs2_busy; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_prs3_busy = exe_reg_uops_1_prs3_busy; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_ppred_busy = exe_reg_uops_1_ppred_busy; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_stale_pdst = exe_reg_uops_1_stale_pdst; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_exception = exe_reg_uops_1_exception; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_exc_cause = exe_reg_uops_1_exc_cause; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_bypassable = exe_reg_uops_1_bypassable; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_mem_cmd = exe_reg_uops_1_mem_cmd; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_mem_size = exe_reg_uops_1_mem_size; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_mem_signed = exe_reg_uops_1_mem_signed; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_is_fence = exe_reg_uops_1_is_fence; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_is_fencei = exe_reg_uops_1_is_fencei; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_is_amo = exe_reg_uops_1_is_amo; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_uses_ldq = exe_reg_uops_1_uses_ldq; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_uses_stq = exe_reg_uops_1_uses_stq; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_is_sys_pc2epc = exe_reg_uops_1_is_sys_pc2epc; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_is_unique = exe_reg_uops_1_is_unique; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_flush_on_commit = exe_reg_uops_1_flush_on_commit; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_ldst_is_rs1 = exe_reg_uops_1_ldst_is_rs1; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_ldst = exe_reg_uops_1_ldst; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_lrs1 = exe_reg_uops_1_lrs1; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_lrs2 = exe_reg_uops_1_lrs2; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_lrs3 = exe_reg_uops_1_lrs3; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_ldst_val = exe_reg_uops_1_ldst_val; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_dst_rtype = exe_reg_uops_1_dst_rtype; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_lrs1_rtype = exe_reg_uops_1_lrs1_rtype; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_lrs2_rtype = exe_reg_uops_1_lrs2_rtype; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_frs3_en = exe_reg_uops_1_frs3_en; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_fp_val = exe_reg_uops_1_fp_val; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_fp_single = exe_reg_uops_1_fp_single; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_xcpt_pf_if = exe_reg_uops_1_xcpt_pf_if; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_xcpt_ae_if = exe_reg_uops_1_xcpt_ae_if; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_xcpt_ma_if = exe_reg_uops_1_xcpt_ma_if; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_bp_debug_if = exe_reg_uops_1_bp_debug_if; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_bp_xcpt_if = exe_reg_uops_1_bp_xcpt_if; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_debug_fsrc = exe_reg_uops_1_debug_fsrc; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_uop_debug_tsrc = exe_reg_uops_1_debug_tsrc; // @[register-read.scala 255:29]
  assign io_exe_reqs_1_bits_rs1_data = exe_reg_rs1_data_1; // @[register-read.scala 256:56]
  assign io_exe_reqs_1_bits_rs2_data = exe_reg_rs2_data_1; // @[register-read.scala 257:56]
  assign io_exe_reqs_1_bits_rs3_data = exe_reg_rs3_data_1; // @[register-read.scala 258:56]
  assign io_exe_reqs_1_bits_pred_data = 1'h0;
  assign io_exe_reqs_1_bits_flagdata = exe_reg_flag_data_1; // @[register-read.scala 261:34]
  assign io_exe_reqs_1_bits_fflagdata = 32'h0;
  assign io_exe_reqs_1_bits_kill = 1'h0;
  assign io_exe_reqs_2_valid = exe_reg_valids_2; // @[register-read.scala 254:29]
  assign io_exe_reqs_2_bits_uop_switch = exe_reg_uops_2_switch; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_switch_off = exe_reg_uops_2_switch_off; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_is_unicore = exe_reg_uops_2_is_unicore; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_shift = exe_reg_uops_2_shift; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_lrs3_rtype = exe_reg_uops_2_lrs3_rtype; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_rflag = exe_reg_uops_2_rflag; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_wflag = exe_reg_uops_2_wflag; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_prflag = exe_reg_uops_2_prflag; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_pwflag = exe_reg_uops_2_pwflag; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_pflag_busy = exe_reg_uops_2_pflag_busy; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_stale_pflag = exe_reg_uops_2_stale_pflag; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_op1_sel = exe_reg_uops_2_op1_sel; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_op2_sel = exe_reg_uops_2_op2_sel; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_split_num = exe_reg_uops_2_split_num; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_self_index = exe_reg_uops_2_self_index; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_rob_inst_idx = exe_reg_uops_2_rob_inst_idx; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_address_num = exe_reg_uops_2_address_num; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_uopc = exe_reg_uops_2_uopc; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_inst = exe_reg_uops_2_inst; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_debug_inst = exe_reg_uops_2_debug_inst; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_is_rvc = exe_reg_uops_2_is_rvc; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_debug_pc = exe_reg_uops_2_debug_pc; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_iq_type = exe_reg_uops_2_iq_type; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_fu_code = exe_reg_uops_2_fu_code; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_ctrl_br_type = exe_reg_uops_2_ctrl_br_type; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_ctrl_op1_sel = exe_reg_uops_2_ctrl_op1_sel; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_ctrl_op2_sel = exe_reg_uops_2_ctrl_op2_sel; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_ctrl_imm_sel = exe_reg_uops_2_ctrl_imm_sel; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_ctrl_op_fcn = exe_reg_uops_2_ctrl_op_fcn; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_ctrl_fcn_dw = exe_reg_uops_2_ctrl_fcn_dw; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_ctrl_csr_cmd = exe_reg_uops_2_ctrl_csr_cmd; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_ctrl_is_load = exe_reg_uops_2_ctrl_is_load; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_ctrl_is_sta = exe_reg_uops_2_ctrl_is_sta; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_ctrl_is_std = exe_reg_uops_2_ctrl_is_std; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_ctrl_op3_sel = exe_reg_uops_2_ctrl_op3_sel; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_iw_state = exe_reg_uops_2_iw_state; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_iw_p1_poisoned = exe_reg_uops_2_iw_p1_poisoned; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_iw_p2_poisoned = exe_reg_uops_2_iw_p2_poisoned; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_is_br = exe_reg_uops_2_is_br; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_is_jalr = exe_reg_uops_2_is_jalr; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_is_jal = exe_reg_uops_2_is_jal; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_is_sfb = exe_reg_uops_2_is_sfb; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_br_mask = exe_reg_uops_2_br_mask; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_br_tag = exe_reg_uops_2_br_tag; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_ftq_idx = exe_reg_uops_2_ftq_idx; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_edge_inst = exe_reg_uops_2_edge_inst; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_pc_lob = exe_reg_uops_2_pc_lob; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_taken = exe_reg_uops_2_taken; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_imm_packed = exe_reg_uops_2_imm_packed; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_csr_addr = exe_reg_uops_2_csr_addr; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_rob_idx = exe_reg_uops_2_rob_idx; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_ldq_idx = exe_reg_uops_2_ldq_idx; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_stq_idx = exe_reg_uops_2_stq_idx; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_rxq_idx = exe_reg_uops_2_rxq_idx; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_pdst = exe_reg_uops_2_pdst; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_prs1 = exe_reg_uops_2_prs1; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_prs2 = exe_reg_uops_2_prs2; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_prs3 = exe_reg_uops_2_prs3; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_ppred = exe_reg_uops_2_ppred; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_prs1_busy = exe_reg_uops_2_prs1_busy; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_prs2_busy = exe_reg_uops_2_prs2_busy; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_prs3_busy = exe_reg_uops_2_prs3_busy; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_ppred_busy = exe_reg_uops_2_ppred_busy; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_stale_pdst = exe_reg_uops_2_stale_pdst; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_exception = exe_reg_uops_2_exception; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_exc_cause = exe_reg_uops_2_exc_cause; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_bypassable = exe_reg_uops_2_bypassable; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_mem_cmd = exe_reg_uops_2_mem_cmd; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_mem_size = exe_reg_uops_2_mem_size; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_mem_signed = exe_reg_uops_2_mem_signed; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_is_fence = exe_reg_uops_2_is_fence; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_is_fencei = exe_reg_uops_2_is_fencei; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_is_amo = exe_reg_uops_2_is_amo; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_uses_ldq = exe_reg_uops_2_uses_ldq; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_uses_stq = exe_reg_uops_2_uses_stq; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_is_sys_pc2epc = exe_reg_uops_2_is_sys_pc2epc; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_is_unique = exe_reg_uops_2_is_unique; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_flush_on_commit = exe_reg_uops_2_flush_on_commit; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_ldst_is_rs1 = exe_reg_uops_2_ldst_is_rs1; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_ldst = exe_reg_uops_2_ldst; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_lrs1 = exe_reg_uops_2_lrs1; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_lrs2 = exe_reg_uops_2_lrs2; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_lrs3 = exe_reg_uops_2_lrs3; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_ldst_val = exe_reg_uops_2_ldst_val; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_dst_rtype = exe_reg_uops_2_dst_rtype; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_lrs1_rtype = exe_reg_uops_2_lrs1_rtype; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_lrs2_rtype = exe_reg_uops_2_lrs2_rtype; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_frs3_en = exe_reg_uops_2_frs3_en; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_fp_val = exe_reg_uops_2_fp_val; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_fp_single = exe_reg_uops_2_fp_single; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_xcpt_pf_if = exe_reg_uops_2_xcpt_pf_if; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_xcpt_ae_if = exe_reg_uops_2_xcpt_ae_if; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_xcpt_ma_if = exe_reg_uops_2_xcpt_ma_if; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_bp_debug_if = exe_reg_uops_2_bp_debug_if; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_bp_xcpt_if = exe_reg_uops_2_bp_xcpt_if; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_debug_fsrc = exe_reg_uops_2_debug_fsrc; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_uop_debug_tsrc = exe_reg_uops_2_debug_tsrc; // @[register-read.scala 255:29]
  assign io_exe_reqs_2_bits_rs1_data = exe_reg_rs1_data_2; // @[register-read.scala 256:56]
  assign io_exe_reqs_2_bits_rs2_data = exe_reg_rs2_data_2; // @[register-read.scala 257:56]
  assign io_exe_reqs_2_bits_rs3_data = exe_reg_rs3_data_2; // @[register-read.scala 258:56]
  assign io_exe_reqs_2_bits_pred_data = 1'h0;
  assign io_exe_reqs_2_bits_flagdata = exe_reg_flag_data_2; // @[register-read.scala 261:34]
  assign io_exe_reqs_2_bits_fflagdata = 32'h0;
  assign io_exe_reqs_2_bits_kill = 1'h0;
  assign RegisterReadDecode_clock = clock;
  assign RegisterReadDecode_reset = reset;
  assign RegisterReadDecode_io_iss_valid = io_iss_valids_0; // @[register-read.scala 87:34]
  assign RegisterReadDecode_io_iss_uop_switch = io_iss_uops_0_switch; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_switch_off = io_iss_uops_0_switch_off; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_is_unicore = io_iss_uops_0_is_unicore; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_shift = io_iss_uops_0_shift; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_lrs3_rtype = io_iss_uops_0_lrs3_rtype; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_rflag = io_iss_uops_0_rflag; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_wflag = io_iss_uops_0_wflag; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_prflag = io_iss_uops_0_prflag; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_pwflag = io_iss_uops_0_pwflag; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_pflag_busy = io_iss_uops_0_pflag_busy; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_stale_pflag = io_iss_uops_0_stale_pflag; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_op1_sel = io_iss_uops_0_op1_sel; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_op2_sel = io_iss_uops_0_op2_sel; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_split_num = io_iss_uops_0_split_num; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_self_index = io_iss_uops_0_self_index; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_rob_inst_idx = io_iss_uops_0_rob_inst_idx; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_address_num = io_iss_uops_0_address_num; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_uopc = io_iss_uops_0_uopc; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_inst = io_iss_uops_0_inst; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_debug_inst = io_iss_uops_0_debug_inst; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_is_rvc = io_iss_uops_0_is_rvc; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_debug_pc = io_iss_uops_0_debug_pc; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_iq_type = io_iss_uops_0_iq_type; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_fu_code = io_iss_uops_0_fu_code; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_ctrl_br_type = io_iss_uops_0_ctrl_br_type; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_ctrl_op1_sel = io_iss_uops_0_ctrl_op1_sel; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_ctrl_op2_sel = io_iss_uops_0_ctrl_op2_sel; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_ctrl_imm_sel = io_iss_uops_0_ctrl_imm_sel; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_ctrl_op_fcn = io_iss_uops_0_ctrl_op_fcn; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_ctrl_fcn_dw = io_iss_uops_0_ctrl_fcn_dw; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_ctrl_csr_cmd = io_iss_uops_0_ctrl_csr_cmd; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_ctrl_is_load = io_iss_uops_0_ctrl_is_load; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_ctrl_is_sta = io_iss_uops_0_ctrl_is_sta; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_ctrl_is_std = io_iss_uops_0_ctrl_is_std; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_ctrl_op3_sel = io_iss_uops_0_ctrl_op3_sel; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_iw_state = io_iss_uops_0_iw_state; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_iw_p1_poisoned = io_iss_uops_0_iw_p1_poisoned; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_iw_p2_poisoned = io_iss_uops_0_iw_p2_poisoned; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_is_br = io_iss_uops_0_is_br; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_is_jalr = io_iss_uops_0_is_jalr; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_is_jal = io_iss_uops_0_is_jal; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_is_sfb = io_iss_uops_0_is_sfb; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_br_mask = io_iss_uops_0_br_mask; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_br_tag = io_iss_uops_0_br_tag; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_ftq_idx = io_iss_uops_0_ftq_idx; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_edge_inst = io_iss_uops_0_edge_inst; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_pc_lob = io_iss_uops_0_pc_lob; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_taken = io_iss_uops_0_taken; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_imm_packed = io_iss_uops_0_imm_packed; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_csr_addr = io_iss_uops_0_csr_addr; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_rob_idx = io_iss_uops_0_rob_idx; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_ldq_idx = io_iss_uops_0_ldq_idx; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_stq_idx = io_iss_uops_0_stq_idx; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_rxq_idx = io_iss_uops_0_rxq_idx; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_pdst = io_iss_uops_0_pdst; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_prs1 = io_iss_uops_0_prs1; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_prs2 = io_iss_uops_0_prs2; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_prs3 = io_iss_uops_0_prs3; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_ppred = io_iss_uops_0_ppred; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_prs1_busy = io_iss_uops_0_prs1_busy; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_prs2_busy = io_iss_uops_0_prs2_busy; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_prs3_busy = io_iss_uops_0_prs3_busy; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_ppred_busy = io_iss_uops_0_ppred_busy; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_stale_pdst = io_iss_uops_0_stale_pdst; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_exception = io_iss_uops_0_exception; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_exc_cause = io_iss_uops_0_exc_cause; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_bypassable = io_iss_uops_0_bypassable; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_mem_cmd = io_iss_uops_0_mem_cmd; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_mem_size = io_iss_uops_0_mem_size; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_mem_signed = io_iss_uops_0_mem_signed; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_is_fence = io_iss_uops_0_is_fence; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_is_fencei = io_iss_uops_0_is_fencei; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_is_amo = io_iss_uops_0_is_amo; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_uses_ldq = io_iss_uops_0_uses_ldq; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_uses_stq = io_iss_uops_0_uses_stq; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_is_sys_pc2epc = io_iss_uops_0_is_sys_pc2epc; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_is_unique = io_iss_uops_0_is_unique; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_flush_on_commit = io_iss_uops_0_flush_on_commit; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_ldst_is_rs1 = io_iss_uops_0_ldst_is_rs1; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_ldst = io_iss_uops_0_ldst; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_lrs1 = io_iss_uops_0_lrs1; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_lrs2 = io_iss_uops_0_lrs2; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_lrs3 = io_iss_uops_0_lrs3; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_ldst_val = io_iss_uops_0_ldst_val; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_dst_rtype = io_iss_uops_0_dst_rtype; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_lrs1_rtype = io_iss_uops_0_lrs1_rtype; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_lrs2_rtype = io_iss_uops_0_lrs2_rtype; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_frs3_en = io_iss_uops_0_frs3_en; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_fp_val = io_iss_uops_0_fp_val; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_fp_single = io_iss_uops_0_fp_single; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_xcpt_pf_if = io_iss_uops_0_xcpt_pf_if; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_xcpt_ae_if = io_iss_uops_0_xcpt_ae_if; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_xcpt_ma_if = io_iss_uops_0_xcpt_ma_if; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_bp_debug_if = io_iss_uops_0_bp_debug_if; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_bp_xcpt_if = io_iss_uops_0_bp_xcpt_if; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_debug_fsrc = io_iss_uops_0_debug_fsrc; // @[register-read.scala 88:34]
  assign RegisterReadDecode_io_iss_uop_debug_tsrc = io_iss_uops_0_debug_tsrc; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_clock = clock;
  assign RegisterReadDecode_1_reset = reset;
  assign RegisterReadDecode_1_io_iss_valid = io_iss_valids_1; // @[register-read.scala 87:34]
  assign RegisterReadDecode_1_io_iss_uop_switch = io_iss_uops_1_switch; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_switch_off = io_iss_uops_1_switch_off; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_is_unicore = io_iss_uops_1_is_unicore; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_shift = io_iss_uops_1_shift; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_lrs3_rtype = io_iss_uops_1_lrs3_rtype; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_rflag = io_iss_uops_1_rflag; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_wflag = io_iss_uops_1_wflag; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_prflag = io_iss_uops_1_prflag; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_pwflag = io_iss_uops_1_pwflag; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_pflag_busy = io_iss_uops_1_pflag_busy; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_stale_pflag = io_iss_uops_1_stale_pflag; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_op1_sel = io_iss_uops_1_op1_sel; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_op2_sel = io_iss_uops_1_op2_sel; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_split_num = io_iss_uops_1_split_num; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_self_index = io_iss_uops_1_self_index; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_rob_inst_idx = io_iss_uops_1_rob_inst_idx; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_address_num = io_iss_uops_1_address_num; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_uopc = io_iss_uops_1_uopc; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_inst = io_iss_uops_1_inst; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_debug_inst = io_iss_uops_1_debug_inst; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_is_rvc = io_iss_uops_1_is_rvc; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_debug_pc = io_iss_uops_1_debug_pc; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_iq_type = io_iss_uops_1_iq_type; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_fu_code = io_iss_uops_1_fu_code; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_ctrl_br_type = io_iss_uops_1_ctrl_br_type; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_ctrl_op1_sel = io_iss_uops_1_ctrl_op1_sel; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_ctrl_op2_sel = io_iss_uops_1_ctrl_op2_sel; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_ctrl_imm_sel = io_iss_uops_1_ctrl_imm_sel; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_ctrl_op_fcn = io_iss_uops_1_ctrl_op_fcn; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_ctrl_fcn_dw = io_iss_uops_1_ctrl_fcn_dw; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_ctrl_csr_cmd = io_iss_uops_1_ctrl_csr_cmd; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_ctrl_is_load = io_iss_uops_1_ctrl_is_load; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_ctrl_is_sta = io_iss_uops_1_ctrl_is_sta; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_ctrl_is_std = io_iss_uops_1_ctrl_is_std; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_ctrl_op3_sel = io_iss_uops_1_ctrl_op3_sel; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_iw_state = io_iss_uops_1_iw_state; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_iw_p1_poisoned = io_iss_uops_1_iw_p1_poisoned; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_iw_p2_poisoned = io_iss_uops_1_iw_p2_poisoned; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_is_br = io_iss_uops_1_is_br; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_is_jalr = io_iss_uops_1_is_jalr; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_is_jal = io_iss_uops_1_is_jal; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_is_sfb = io_iss_uops_1_is_sfb; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_br_mask = io_iss_uops_1_br_mask; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_br_tag = io_iss_uops_1_br_tag; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_ftq_idx = io_iss_uops_1_ftq_idx; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_edge_inst = io_iss_uops_1_edge_inst; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_pc_lob = io_iss_uops_1_pc_lob; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_taken = io_iss_uops_1_taken; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_imm_packed = io_iss_uops_1_imm_packed; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_csr_addr = io_iss_uops_1_csr_addr; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_rob_idx = io_iss_uops_1_rob_idx; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_ldq_idx = io_iss_uops_1_ldq_idx; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_stq_idx = io_iss_uops_1_stq_idx; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_rxq_idx = io_iss_uops_1_rxq_idx; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_pdst = io_iss_uops_1_pdst; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_prs1 = io_iss_uops_1_prs1; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_prs2 = io_iss_uops_1_prs2; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_prs3 = io_iss_uops_1_prs3; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_ppred = io_iss_uops_1_ppred; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_prs1_busy = io_iss_uops_1_prs1_busy; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_prs2_busy = io_iss_uops_1_prs2_busy; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_prs3_busy = io_iss_uops_1_prs3_busy; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_ppred_busy = io_iss_uops_1_ppred_busy; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_stale_pdst = io_iss_uops_1_stale_pdst; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_exception = io_iss_uops_1_exception; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_exc_cause = io_iss_uops_1_exc_cause; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_bypassable = io_iss_uops_1_bypassable; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_mem_cmd = io_iss_uops_1_mem_cmd; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_mem_size = io_iss_uops_1_mem_size; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_mem_signed = io_iss_uops_1_mem_signed; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_is_fence = io_iss_uops_1_is_fence; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_is_fencei = io_iss_uops_1_is_fencei; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_is_amo = io_iss_uops_1_is_amo; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_uses_ldq = io_iss_uops_1_uses_ldq; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_uses_stq = io_iss_uops_1_uses_stq; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_is_sys_pc2epc = io_iss_uops_1_is_sys_pc2epc; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_is_unique = io_iss_uops_1_is_unique; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_flush_on_commit = io_iss_uops_1_flush_on_commit; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_ldst_is_rs1 = io_iss_uops_1_ldst_is_rs1; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_ldst = io_iss_uops_1_ldst; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_lrs1 = io_iss_uops_1_lrs1; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_lrs2 = io_iss_uops_1_lrs2; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_lrs3 = io_iss_uops_1_lrs3; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_ldst_val = io_iss_uops_1_ldst_val; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_dst_rtype = io_iss_uops_1_dst_rtype; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_lrs1_rtype = io_iss_uops_1_lrs1_rtype; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_lrs2_rtype = io_iss_uops_1_lrs2_rtype; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_frs3_en = io_iss_uops_1_frs3_en; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_fp_val = io_iss_uops_1_fp_val; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_fp_single = io_iss_uops_1_fp_single; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_xcpt_pf_if = io_iss_uops_1_xcpt_pf_if; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_xcpt_ae_if = io_iss_uops_1_xcpt_ae_if; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_xcpt_ma_if = io_iss_uops_1_xcpt_ma_if; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_bp_debug_if = io_iss_uops_1_bp_debug_if; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_bp_xcpt_if = io_iss_uops_1_bp_xcpt_if; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_debug_fsrc = io_iss_uops_1_debug_fsrc; // @[register-read.scala 88:34]
  assign RegisterReadDecode_1_io_iss_uop_debug_tsrc = io_iss_uops_1_debug_tsrc; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_clock = clock;
  assign RegisterReadDecode_2_reset = reset;
  assign RegisterReadDecode_2_io_iss_valid = io_iss_valids_2; // @[register-read.scala 87:34]
  assign RegisterReadDecode_2_io_iss_uop_switch = io_iss_uops_2_switch; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_switch_off = io_iss_uops_2_switch_off; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_is_unicore = io_iss_uops_2_is_unicore; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_shift = io_iss_uops_2_shift; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_lrs3_rtype = io_iss_uops_2_lrs3_rtype; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_rflag = io_iss_uops_2_rflag; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_wflag = io_iss_uops_2_wflag; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_prflag = io_iss_uops_2_prflag; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_pwflag = io_iss_uops_2_pwflag; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_pflag_busy = io_iss_uops_2_pflag_busy; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_stale_pflag = io_iss_uops_2_stale_pflag; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_op1_sel = io_iss_uops_2_op1_sel; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_op2_sel = io_iss_uops_2_op2_sel; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_split_num = io_iss_uops_2_split_num; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_self_index = io_iss_uops_2_self_index; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_rob_inst_idx = io_iss_uops_2_rob_inst_idx; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_address_num = io_iss_uops_2_address_num; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_uopc = io_iss_uops_2_uopc; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_inst = io_iss_uops_2_inst; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_debug_inst = io_iss_uops_2_debug_inst; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_is_rvc = io_iss_uops_2_is_rvc; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_debug_pc = io_iss_uops_2_debug_pc; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_iq_type = io_iss_uops_2_iq_type; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_fu_code = io_iss_uops_2_fu_code; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_ctrl_br_type = io_iss_uops_2_ctrl_br_type; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_ctrl_op1_sel = io_iss_uops_2_ctrl_op1_sel; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_ctrl_op2_sel = io_iss_uops_2_ctrl_op2_sel; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_ctrl_imm_sel = io_iss_uops_2_ctrl_imm_sel; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_ctrl_op_fcn = io_iss_uops_2_ctrl_op_fcn; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_ctrl_fcn_dw = io_iss_uops_2_ctrl_fcn_dw; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_ctrl_csr_cmd = io_iss_uops_2_ctrl_csr_cmd; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_ctrl_is_load = io_iss_uops_2_ctrl_is_load; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_ctrl_is_sta = io_iss_uops_2_ctrl_is_sta; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_ctrl_is_std = io_iss_uops_2_ctrl_is_std; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_ctrl_op3_sel = io_iss_uops_2_ctrl_op3_sel; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_iw_state = io_iss_uops_2_iw_state; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_iw_p1_poisoned = io_iss_uops_2_iw_p1_poisoned; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_iw_p2_poisoned = io_iss_uops_2_iw_p2_poisoned; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_is_br = io_iss_uops_2_is_br; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_is_jalr = io_iss_uops_2_is_jalr; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_is_jal = io_iss_uops_2_is_jal; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_is_sfb = io_iss_uops_2_is_sfb; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_br_mask = io_iss_uops_2_br_mask; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_br_tag = io_iss_uops_2_br_tag; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_ftq_idx = io_iss_uops_2_ftq_idx; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_edge_inst = io_iss_uops_2_edge_inst; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_pc_lob = io_iss_uops_2_pc_lob; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_taken = io_iss_uops_2_taken; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_imm_packed = io_iss_uops_2_imm_packed; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_csr_addr = io_iss_uops_2_csr_addr; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_rob_idx = io_iss_uops_2_rob_idx; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_ldq_idx = io_iss_uops_2_ldq_idx; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_stq_idx = io_iss_uops_2_stq_idx; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_rxq_idx = io_iss_uops_2_rxq_idx; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_pdst = io_iss_uops_2_pdst; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_prs1 = io_iss_uops_2_prs1; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_prs2 = io_iss_uops_2_prs2; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_prs3 = io_iss_uops_2_prs3; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_ppred = io_iss_uops_2_ppred; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_prs1_busy = io_iss_uops_2_prs1_busy; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_prs2_busy = io_iss_uops_2_prs2_busy; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_prs3_busy = io_iss_uops_2_prs3_busy; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_ppred_busy = io_iss_uops_2_ppred_busy; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_stale_pdst = io_iss_uops_2_stale_pdst; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_exception = io_iss_uops_2_exception; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_exc_cause = io_iss_uops_2_exc_cause; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_bypassable = io_iss_uops_2_bypassable; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_mem_cmd = io_iss_uops_2_mem_cmd; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_mem_size = io_iss_uops_2_mem_size; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_mem_signed = io_iss_uops_2_mem_signed; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_is_fence = io_iss_uops_2_is_fence; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_is_fencei = io_iss_uops_2_is_fencei; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_is_amo = io_iss_uops_2_is_amo; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_uses_ldq = io_iss_uops_2_uses_ldq; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_uses_stq = io_iss_uops_2_uses_stq; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_is_sys_pc2epc = io_iss_uops_2_is_sys_pc2epc; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_is_unique = io_iss_uops_2_is_unique; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_flush_on_commit = io_iss_uops_2_flush_on_commit; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_ldst_is_rs1 = io_iss_uops_2_ldst_is_rs1; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_ldst = io_iss_uops_2_ldst; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_lrs1 = io_iss_uops_2_lrs1; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_lrs2 = io_iss_uops_2_lrs2; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_lrs3 = io_iss_uops_2_lrs3; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_ldst_val = io_iss_uops_2_ldst_val; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_dst_rtype = io_iss_uops_2_dst_rtype; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_lrs1_rtype = io_iss_uops_2_lrs1_rtype; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_lrs2_rtype = io_iss_uops_2_lrs2_rtype; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_frs3_en = io_iss_uops_2_frs3_en; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_fp_val = io_iss_uops_2_fp_val; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_fp_single = io_iss_uops_2_fp_single; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_xcpt_pf_if = io_iss_uops_2_xcpt_pf_if; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_xcpt_ae_if = io_iss_uops_2_xcpt_ae_if; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_xcpt_ma_if = io_iss_uops_2_xcpt_ma_if; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_bp_debug_if = io_iss_uops_2_bp_debug_if; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_bp_xcpt_if = io_iss_uops_2_bp_xcpt_if; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_debug_fsrc = io_iss_uops_2_debug_fsrc; // @[register-read.scala 88:34]
  assign RegisterReadDecode_2_io_iss_uop_debug_tsrc = io_iss_uops_2_debug_tsrc; // @[register-read.scala 88:34]
  always @(posedge clock) begin
    if (reset) begin // @[register-read.scala 72:33]
      exe_reg_valids_0 <= 1'h0; // @[register-read.scala 72:33]
    end else if (_T_34) begin // @[register-read.scala 147:29]
      exe_reg_valids_0 <= 1'h0;
    end else begin
      exe_reg_valids_0 <= REG;
    end
    if (reset) begin // @[register-read.scala 72:33]
      exe_reg_valids_1 <= 1'h0; // @[register-read.scala 72:33]
    end else if (_T_55) begin // @[register-read.scala 147:29]
      exe_reg_valids_1 <= 1'h0;
    end else begin
      exe_reg_valids_1 <= REG_2;
    end
    if (reset) begin // @[register-read.scala 72:33]
      exe_reg_valids_2 <= 1'h0; // @[register-read.scala 72:33]
    end else if (_T_76) begin // @[register-read.scala 147:29]
      exe_reg_valids_2 <= 1'h0;
    end else begin
      exe_reg_valids_2 <= REG_4;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_switch <= 1'h0;
    end else begin
      exe_reg_uops_0_switch <= REG_1_switch;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_switch_off <= 1'h0;
    end else begin
      exe_reg_uops_0_switch_off <= REG_1_switch_off;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_is_unicore <= 1'h0;
    end else begin
      exe_reg_uops_0_is_unicore <= REG_1_is_unicore;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_shift <= 3'h0;
    end else begin
      exe_reg_uops_0_shift <= REG_1_shift;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_lrs3_rtype <= 2'h0;
    end else begin
      exe_reg_uops_0_lrs3_rtype <= REG_1_lrs3_rtype;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_rflag <= 1'h0;
    end else begin
      exe_reg_uops_0_rflag <= REG_1_rflag;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_wflag <= 1'h0;
    end else begin
      exe_reg_uops_0_wflag <= REG_1_wflag;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_prflag <= 4'h0;
    end else begin
      exe_reg_uops_0_prflag <= REG_1_prflag;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_pwflag <= 4'h0;
    end else begin
      exe_reg_uops_0_pwflag <= REG_1_pwflag;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_pflag_busy <= 1'h0;
    end else begin
      exe_reg_uops_0_pflag_busy <= REG_1_pflag_busy;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_stale_pflag <= 4'h0;
    end else begin
      exe_reg_uops_0_stale_pflag <= REG_1_stale_pflag;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_op1_sel <= 4'h0;
    end else begin
      exe_reg_uops_0_op1_sel <= REG_1_op1_sel;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_op2_sel <= 4'h0;
    end else begin
      exe_reg_uops_0_op2_sel <= REG_1_op2_sel;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_split_num <= 6'h0;
    end else begin
      exe_reg_uops_0_split_num <= REG_1_split_num;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_self_index <= 6'h0;
    end else begin
      exe_reg_uops_0_self_index <= REG_1_self_index;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_rob_inst_idx <= 6'h0;
    end else begin
      exe_reg_uops_0_rob_inst_idx <= REG_1_rob_inst_idx;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_address_num <= 6'h0;
    end else begin
      exe_reg_uops_0_address_num <= REG_1_address_num;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_uopc <= 7'h0;
    end else begin
      exe_reg_uops_0_uopc <= REG_1_uopc;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_inst <= 32'h0;
    end else begin
      exe_reg_uops_0_inst <= REG_1_inst;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_debug_inst <= 32'h0;
    end else begin
      exe_reg_uops_0_debug_inst <= REG_1_debug_inst;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_is_rvc <= 1'h0;
    end else begin
      exe_reg_uops_0_is_rvc <= REG_1_is_rvc;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_debug_pc <= 40'h0;
    end else begin
      exe_reg_uops_0_debug_pc <= REG_1_debug_pc;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_iq_type <= 3'h0;
    end else begin
      exe_reg_uops_0_iq_type <= REG_1_iq_type;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_fu_code <= 10'h0;
    end else begin
      exe_reg_uops_0_fu_code <= REG_1_fu_code;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_ctrl_br_type <= 4'h0;
    end else begin
      exe_reg_uops_0_ctrl_br_type <= REG_1_ctrl_br_type;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_ctrl_op1_sel <= 2'h0;
    end else begin
      exe_reg_uops_0_ctrl_op1_sel <= REG_1_ctrl_op1_sel;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_ctrl_op2_sel <= 3'h0;
    end else begin
      exe_reg_uops_0_ctrl_op2_sel <= REG_1_ctrl_op2_sel;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_ctrl_imm_sel <= 3'h0;
    end else begin
      exe_reg_uops_0_ctrl_imm_sel <= REG_1_ctrl_imm_sel;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_ctrl_op_fcn <= 4'h0;
    end else begin
      exe_reg_uops_0_ctrl_op_fcn <= REG_1_ctrl_op_fcn;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_ctrl_fcn_dw <= 1'h0;
    end else begin
      exe_reg_uops_0_ctrl_fcn_dw <= REG_1_ctrl_fcn_dw;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_ctrl_csr_cmd <= 3'h0;
    end else begin
      exe_reg_uops_0_ctrl_csr_cmd <= REG_1_ctrl_csr_cmd;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_ctrl_is_load <= 1'h0;
    end else begin
      exe_reg_uops_0_ctrl_is_load <= REG_1_ctrl_is_load;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_ctrl_is_sta <= 1'h0;
    end else begin
      exe_reg_uops_0_ctrl_is_sta <= REG_1_ctrl_is_sta;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_ctrl_is_std <= 1'h0;
    end else begin
      exe_reg_uops_0_ctrl_is_std <= REG_1_ctrl_is_std;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_ctrl_op3_sel <= 2'h0;
    end else begin
      exe_reg_uops_0_ctrl_op3_sel <= REG_1_ctrl_op3_sel;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_iw_state <= 2'h0;
    end else begin
      exe_reg_uops_0_iw_state <= REG_1_iw_state;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_iw_p1_poisoned <= 1'h0;
    end else begin
      exe_reg_uops_0_iw_p1_poisoned <= REG_1_iw_p1_poisoned;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_iw_p2_poisoned <= 1'h0;
    end else begin
      exe_reg_uops_0_iw_p2_poisoned <= REG_1_iw_p2_poisoned;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_is_br <= 1'h0;
    end else begin
      exe_reg_uops_0_is_br <= REG_1_is_br;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_is_jalr <= 1'h0;
    end else begin
      exe_reg_uops_0_is_jalr <= REG_1_is_jalr;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_is_jal <= 1'h0;
    end else begin
      exe_reg_uops_0_is_jal <= REG_1_is_jal;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_is_sfb <= 1'h0;
    end else begin
      exe_reg_uops_0_is_sfb <= REG_1_is_sfb;
    end
    exe_reg_uops_0_br_mask <= REG_1_br_mask & _T_4; // @[util.scala 142:25]
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_br_tag <= 4'h0;
    end else begin
      exe_reg_uops_0_br_tag <= REG_1_br_tag;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_ftq_idx <= 5'h0;
    end else begin
      exe_reg_uops_0_ftq_idx <= REG_1_ftq_idx;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_edge_inst <= 1'h0;
    end else begin
      exe_reg_uops_0_edge_inst <= REG_1_edge_inst;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_pc_lob <= 6'h0;
    end else begin
      exe_reg_uops_0_pc_lob <= REG_1_pc_lob;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_taken <= 1'h0;
    end else begin
      exe_reg_uops_0_taken <= REG_1_taken;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_imm_packed <= 20'h0;
    end else begin
      exe_reg_uops_0_imm_packed <= REG_1_imm_packed;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_csr_addr <= 12'h0;
    end else begin
      exe_reg_uops_0_csr_addr <= REG_1_csr_addr;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_rob_idx <= 6'h0;
    end else begin
      exe_reg_uops_0_rob_idx <= REG_1_rob_idx;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_ldq_idx <= 5'h0;
    end else begin
      exe_reg_uops_0_ldq_idx <= REG_1_ldq_idx;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_stq_idx <= 5'h0;
    end else begin
      exe_reg_uops_0_stq_idx <= REG_1_stq_idx;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_rxq_idx <= 2'h0;
    end else begin
      exe_reg_uops_0_rxq_idx <= REG_1_rxq_idx;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_pdst <= 7'h0;
    end else begin
      exe_reg_uops_0_pdst <= REG_1_pdst;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_prs1 <= 7'h0;
    end else begin
      exe_reg_uops_0_prs1 <= REG_1_prs1;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_prs2 <= 7'h0;
    end else begin
      exe_reg_uops_0_prs2 <= REG_1_prs2;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_prs3 <= 7'h0;
    end else begin
      exe_reg_uops_0_prs3 <= REG_1_prs3;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_ppred <= 5'h0;
    end else begin
      exe_reg_uops_0_ppred <= REG_1_ppred;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_prs1_busy <= 1'h0;
    end else begin
      exe_reg_uops_0_prs1_busy <= REG_1_prs1_busy;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_prs2_busy <= 1'h0;
    end else begin
      exe_reg_uops_0_prs2_busy <= REG_1_prs2_busy;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_prs3_busy <= 1'h0;
    end else begin
      exe_reg_uops_0_prs3_busy <= REG_1_prs3_busy;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_ppred_busy <= 1'h0;
    end else begin
      exe_reg_uops_0_ppred_busy <= REG_1_ppred_busy;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_stale_pdst <= 7'h0;
    end else begin
      exe_reg_uops_0_stale_pdst <= REG_1_stale_pdst;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_exception <= 1'h0;
    end else begin
      exe_reg_uops_0_exception <= REG_1_exception;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_exc_cause <= 64'h0;
    end else begin
      exe_reg_uops_0_exc_cause <= REG_1_exc_cause;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_bypassable <= 1'h0;
    end else begin
      exe_reg_uops_0_bypassable <= REG_1_bypassable;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_mem_cmd <= 5'h0;
    end else begin
      exe_reg_uops_0_mem_cmd <= REG_1_mem_cmd;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_mem_size <= 2'h0;
    end else begin
      exe_reg_uops_0_mem_size <= REG_1_mem_size;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_mem_signed <= 1'h0;
    end else begin
      exe_reg_uops_0_mem_signed <= REG_1_mem_signed;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_is_fence <= 1'h0;
    end else begin
      exe_reg_uops_0_is_fence <= REG_1_is_fence;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_is_fencei <= 1'h0;
    end else begin
      exe_reg_uops_0_is_fencei <= REG_1_is_fencei;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_is_amo <= 1'h0;
    end else begin
      exe_reg_uops_0_is_amo <= REG_1_is_amo;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_uses_ldq <= 1'h0;
    end else begin
      exe_reg_uops_0_uses_ldq <= REG_1_uses_ldq;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_uses_stq <= 1'h0;
    end else begin
      exe_reg_uops_0_uses_stq <= REG_1_uses_stq;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_is_sys_pc2epc <= 1'h0;
    end else begin
      exe_reg_uops_0_is_sys_pc2epc <= REG_1_is_sys_pc2epc;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_is_unique <= 1'h0;
    end else begin
      exe_reg_uops_0_is_unique <= REG_1_is_unique;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_flush_on_commit <= 1'h0;
    end else begin
      exe_reg_uops_0_flush_on_commit <= REG_1_flush_on_commit;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_ldst_is_rs1 <= 1'h0;
    end else begin
      exe_reg_uops_0_ldst_is_rs1 <= REG_1_ldst_is_rs1;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_ldst <= 6'h0;
    end else begin
      exe_reg_uops_0_ldst <= REG_1_ldst;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_lrs1 <= 6'h0;
    end else begin
      exe_reg_uops_0_lrs1 <= REG_1_lrs1;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_lrs2 <= 6'h0;
    end else begin
      exe_reg_uops_0_lrs2 <= REG_1_lrs2;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_lrs3 <= 6'h0;
    end else begin
      exe_reg_uops_0_lrs3 <= REG_1_lrs3;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_ldst_val <= 1'h0;
    end else begin
      exe_reg_uops_0_ldst_val <= REG_1_ldst_val;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_dst_rtype <= 2'h2;
    end else begin
      exe_reg_uops_0_dst_rtype <= REG_1_dst_rtype;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_lrs1_rtype <= 2'h0;
    end else begin
      exe_reg_uops_0_lrs1_rtype <= REG_1_lrs1_rtype;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_lrs2_rtype <= 2'h0;
    end else begin
      exe_reg_uops_0_lrs2_rtype <= REG_1_lrs2_rtype;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_frs3_en <= 1'h0;
    end else begin
      exe_reg_uops_0_frs3_en <= REG_1_frs3_en;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_fp_val <= 1'h0;
    end else begin
      exe_reg_uops_0_fp_val <= REG_1_fp_val;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_fp_single <= 1'h0;
    end else begin
      exe_reg_uops_0_fp_single <= REG_1_fp_single;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_xcpt_pf_if <= 1'h0;
    end else begin
      exe_reg_uops_0_xcpt_pf_if <= REG_1_xcpt_pf_if;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_xcpt_ae_if <= 1'h0;
    end else begin
      exe_reg_uops_0_xcpt_ae_if <= REG_1_xcpt_ae_if;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_xcpt_ma_if <= 1'h0;
    end else begin
      exe_reg_uops_0_xcpt_ma_if <= REG_1_xcpt_ma_if;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_bp_debug_if <= 1'h0;
    end else begin
      exe_reg_uops_0_bp_debug_if <= REG_1_bp_debug_if;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_bp_xcpt_if <= 1'h0;
    end else begin
      exe_reg_uops_0_bp_xcpt_if <= REG_1_bp_xcpt_if;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_debug_fsrc <= 2'h0;
    end else begin
      exe_reg_uops_0_debug_fsrc <= REG_1_debug_fsrc;
    end
    if (_T_34) begin // @[register-read.scala 149:29]
      exe_reg_uops_0_debug_tsrc <= 2'h0;
    end else begin
      exe_reg_uops_0_debug_tsrc <= REG_1_debug_tsrc;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_switch <= 1'h0;
    end else begin
      exe_reg_uops_1_switch <= REG_3_switch;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_switch_off <= 1'h0;
    end else begin
      exe_reg_uops_1_switch_off <= REG_3_switch_off;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_is_unicore <= 1'h0;
    end else begin
      exe_reg_uops_1_is_unicore <= REG_3_is_unicore;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_shift <= 3'h0;
    end else begin
      exe_reg_uops_1_shift <= REG_3_shift;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_lrs3_rtype <= 2'h0;
    end else begin
      exe_reg_uops_1_lrs3_rtype <= REG_3_lrs3_rtype;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_rflag <= 1'h0;
    end else begin
      exe_reg_uops_1_rflag <= REG_3_rflag;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_wflag <= 1'h0;
    end else begin
      exe_reg_uops_1_wflag <= REG_3_wflag;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_prflag <= 4'h0;
    end else begin
      exe_reg_uops_1_prflag <= REG_3_prflag;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_pwflag <= 4'h0;
    end else begin
      exe_reg_uops_1_pwflag <= REG_3_pwflag;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_pflag_busy <= 1'h0;
    end else begin
      exe_reg_uops_1_pflag_busy <= REG_3_pflag_busy;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_stale_pflag <= 4'h0;
    end else begin
      exe_reg_uops_1_stale_pflag <= REG_3_stale_pflag;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_op1_sel <= 4'h0;
    end else begin
      exe_reg_uops_1_op1_sel <= REG_3_op1_sel;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_op2_sel <= 4'h0;
    end else begin
      exe_reg_uops_1_op2_sel <= REG_3_op2_sel;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_split_num <= 6'h0;
    end else begin
      exe_reg_uops_1_split_num <= REG_3_split_num;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_self_index <= 6'h0;
    end else begin
      exe_reg_uops_1_self_index <= REG_3_self_index;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_rob_inst_idx <= 6'h0;
    end else begin
      exe_reg_uops_1_rob_inst_idx <= REG_3_rob_inst_idx;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_address_num <= 6'h0;
    end else begin
      exe_reg_uops_1_address_num <= REG_3_address_num;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_uopc <= 7'h0;
    end else begin
      exe_reg_uops_1_uopc <= REG_3_uopc;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_inst <= 32'h0;
    end else begin
      exe_reg_uops_1_inst <= REG_3_inst;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_debug_inst <= 32'h0;
    end else begin
      exe_reg_uops_1_debug_inst <= REG_3_debug_inst;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_is_rvc <= 1'h0;
    end else begin
      exe_reg_uops_1_is_rvc <= REG_3_is_rvc;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_debug_pc <= 40'h0;
    end else begin
      exe_reg_uops_1_debug_pc <= REG_3_debug_pc;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_iq_type <= 3'h0;
    end else begin
      exe_reg_uops_1_iq_type <= REG_3_iq_type;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_fu_code <= 10'h0;
    end else begin
      exe_reg_uops_1_fu_code <= REG_3_fu_code;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_ctrl_br_type <= 4'h0;
    end else begin
      exe_reg_uops_1_ctrl_br_type <= REG_3_ctrl_br_type;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_ctrl_op1_sel <= 2'h0;
    end else begin
      exe_reg_uops_1_ctrl_op1_sel <= REG_3_ctrl_op1_sel;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_ctrl_op2_sel <= 3'h0;
    end else begin
      exe_reg_uops_1_ctrl_op2_sel <= REG_3_ctrl_op2_sel;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_ctrl_imm_sel <= 3'h0;
    end else begin
      exe_reg_uops_1_ctrl_imm_sel <= REG_3_ctrl_imm_sel;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_ctrl_op_fcn <= 4'h0;
    end else begin
      exe_reg_uops_1_ctrl_op_fcn <= REG_3_ctrl_op_fcn;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_ctrl_fcn_dw <= 1'h0;
    end else begin
      exe_reg_uops_1_ctrl_fcn_dw <= REG_3_ctrl_fcn_dw;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_ctrl_csr_cmd <= 3'h0;
    end else begin
      exe_reg_uops_1_ctrl_csr_cmd <= REG_3_ctrl_csr_cmd;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_ctrl_is_load <= 1'h0;
    end else begin
      exe_reg_uops_1_ctrl_is_load <= REG_3_ctrl_is_load;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_ctrl_is_sta <= 1'h0;
    end else begin
      exe_reg_uops_1_ctrl_is_sta <= REG_3_ctrl_is_sta;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_ctrl_is_std <= 1'h0;
    end else begin
      exe_reg_uops_1_ctrl_is_std <= REG_3_ctrl_is_std;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_ctrl_op3_sel <= 2'h0;
    end else begin
      exe_reg_uops_1_ctrl_op3_sel <= REG_3_ctrl_op3_sel;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_iw_state <= 2'h0;
    end else begin
      exe_reg_uops_1_iw_state <= REG_3_iw_state;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_iw_p1_poisoned <= 1'h0;
    end else begin
      exe_reg_uops_1_iw_p1_poisoned <= REG_3_iw_p1_poisoned;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_iw_p2_poisoned <= 1'h0;
    end else begin
      exe_reg_uops_1_iw_p2_poisoned <= REG_3_iw_p2_poisoned;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_is_br <= 1'h0;
    end else begin
      exe_reg_uops_1_is_br <= REG_3_is_br;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_is_jalr <= 1'h0;
    end else begin
      exe_reg_uops_1_is_jalr <= REG_3_is_jalr;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_is_jal <= 1'h0;
    end else begin
      exe_reg_uops_1_is_jal <= REG_3_is_jal;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_is_sfb <= 1'h0;
    end else begin
      exe_reg_uops_1_is_sfb <= REG_3_is_sfb;
    end
    exe_reg_uops_1_br_mask <= REG_3_br_mask & _T_4; // @[util.scala 142:25]
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_br_tag <= 4'h0;
    end else begin
      exe_reg_uops_1_br_tag <= REG_3_br_tag;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_ftq_idx <= 5'h0;
    end else begin
      exe_reg_uops_1_ftq_idx <= REG_3_ftq_idx;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_edge_inst <= 1'h0;
    end else begin
      exe_reg_uops_1_edge_inst <= REG_3_edge_inst;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_pc_lob <= 6'h0;
    end else begin
      exe_reg_uops_1_pc_lob <= REG_3_pc_lob;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_taken <= 1'h0;
    end else begin
      exe_reg_uops_1_taken <= REG_3_taken;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_imm_packed <= 20'h0;
    end else begin
      exe_reg_uops_1_imm_packed <= REG_3_imm_packed;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_csr_addr <= 12'h0;
    end else begin
      exe_reg_uops_1_csr_addr <= REG_3_csr_addr;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_rob_idx <= 6'h0;
    end else begin
      exe_reg_uops_1_rob_idx <= REG_3_rob_idx;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_ldq_idx <= 5'h0;
    end else begin
      exe_reg_uops_1_ldq_idx <= REG_3_ldq_idx;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_stq_idx <= 5'h0;
    end else begin
      exe_reg_uops_1_stq_idx <= REG_3_stq_idx;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_rxq_idx <= 2'h0;
    end else begin
      exe_reg_uops_1_rxq_idx <= REG_3_rxq_idx;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_pdst <= 7'h0;
    end else begin
      exe_reg_uops_1_pdst <= REG_3_pdst;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_prs1 <= 7'h0;
    end else begin
      exe_reg_uops_1_prs1 <= REG_3_prs1;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_prs2 <= 7'h0;
    end else begin
      exe_reg_uops_1_prs2 <= REG_3_prs2;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_prs3 <= 7'h0;
    end else begin
      exe_reg_uops_1_prs3 <= REG_3_prs3;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_ppred <= 5'h0;
    end else begin
      exe_reg_uops_1_ppred <= REG_3_ppred;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_prs1_busy <= 1'h0;
    end else begin
      exe_reg_uops_1_prs1_busy <= REG_3_prs1_busy;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_prs2_busy <= 1'h0;
    end else begin
      exe_reg_uops_1_prs2_busy <= REG_3_prs2_busy;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_prs3_busy <= 1'h0;
    end else begin
      exe_reg_uops_1_prs3_busy <= REG_3_prs3_busy;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_ppred_busy <= 1'h0;
    end else begin
      exe_reg_uops_1_ppred_busy <= REG_3_ppred_busy;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_stale_pdst <= 7'h0;
    end else begin
      exe_reg_uops_1_stale_pdst <= REG_3_stale_pdst;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_exception <= 1'h0;
    end else begin
      exe_reg_uops_1_exception <= REG_3_exception;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_exc_cause <= 64'h0;
    end else begin
      exe_reg_uops_1_exc_cause <= REG_3_exc_cause;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_bypassable <= 1'h0;
    end else begin
      exe_reg_uops_1_bypassable <= REG_3_bypassable;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_mem_cmd <= 5'h0;
    end else begin
      exe_reg_uops_1_mem_cmd <= REG_3_mem_cmd;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_mem_size <= 2'h0;
    end else begin
      exe_reg_uops_1_mem_size <= REG_3_mem_size;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_mem_signed <= 1'h0;
    end else begin
      exe_reg_uops_1_mem_signed <= REG_3_mem_signed;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_is_fence <= 1'h0;
    end else begin
      exe_reg_uops_1_is_fence <= REG_3_is_fence;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_is_fencei <= 1'h0;
    end else begin
      exe_reg_uops_1_is_fencei <= REG_3_is_fencei;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_is_amo <= 1'h0;
    end else begin
      exe_reg_uops_1_is_amo <= REG_3_is_amo;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_uses_ldq <= 1'h0;
    end else begin
      exe_reg_uops_1_uses_ldq <= REG_3_uses_ldq;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_uses_stq <= 1'h0;
    end else begin
      exe_reg_uops_1_uses_stq <= REG_3_uses_stq;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_is_sys_pc2epc <= 1'h0;
    end else begin
      exe_reg_uops_1_is_sys_pc2epc <= REG_3_is_sys_pc2epc;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_is_unique <= 1'h0;
    end else begin
      exe_reg_uops_1_is_unique <= REG_3_is_unique;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_flush_on_commit <= 1'h0;
    end else begin
      exe_reg_uops_1_flush_on_commit <= REG_3_flush_on_commit;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_ldst_is_rs1 <= 1'h0;
    end else begin
      exe_reg_uops_1_ldst_is_rs1 <= REG_3_ldst_is_rs1;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_ldst <= 6'h0;
    end else begin
      exe_reg_uops_1_ldst <= REG_3_ldst;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_lrs1 <= 6'h0;
    end else begin
      exe_reg_uops_1_lrs1 <= REG_3_lrs1;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_lrs2 <= 6'h0;
    end else begin
      exe_reg_uops_1_lrs2 <= REG_3_lrs2;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_lrs3 <= 6'h0;
    end else begin
      exe_reg_uops_1_lrs3 <= REG_3_lrs3;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_ldst_val <= 1'h0;
    end else begin
      exe_reg_uops_1_ldst_val <= REG_3_ldst_val;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_dst_rtype <= 2'h2;
    end else begin
      exe_reg_uops_1_dst_rtype <= REG_3_dst_rtype;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_lrs1_rtype <= 2'h0;
    end else begin
      exe_reg_uops_1_lrs1_rtype <= REG_3_lrs1_rtype;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_lrs2_rtype <= 2'h0;
    end else begin
      exe_reg_uops_1_lrs2_rtype <= REG_3_lrs2_rtype;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_frs3_en <= 1'h0;
    end else begin
      exe_reg_uops_1_frs3_en <= REG_3_frs3_en;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_fp_val <= 1'h0;
    end else begin
      exe_reg_uops_1_fp_val <= REG_3_fp_val;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_fp_single <= 1'h0;
    end else begin
      exe_reg_uops_1_fp_single <= REG_3_fp_single;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_xcpt_pf_if <= 1'h0;
    end else begin
      exe_reg_uops_1_xcpt_pf_if <= REG_3_xcpt_pf_if;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_xcpt_ae_if <= 1'h0;
    end else begin
      exe_reg_uops_1_xcpt_ae_if <= REG_3_xcpt_ae_if;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_xcpt_ma_if <= 1'h0;
    end else begin
      exe_reg_uops_1_xcpt_ma_if <= REG_3_xcpt_ma_if;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_bp_debug_if <= 1'h0;
    end else begin
      exe_reg_uops_1_bp_debug_if <= REG_3_bp_debug_if;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_bp_xcpt_if <= 1'h0;
    end else begin
      exe_reg_uops_1_bp_xcpt_if <= REG_3_bp_xcpt_if;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_debug_fsrc <= 2'h0;
    end else begin
      exe_reg_uops_1_debug_fsrc <= REG_3_debug_fsrc;
    end
    if (_T_55) begin // @[register-read.scala 149:29]
      exe_reg_uops_1_debug_tsrc <= 2'h0;
    end else begin
      exe_reg_uops_1_debug_tsrc <= REG_3_debug_tsrc;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_switch <= 1'h0;
    end else begin
      exe_reg_uops_2_switch <= REG_5_switch;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_switch_off <= 1'h0;
    end else begin
      exe_reg_uops_2_switch_off <= REG_5_switch_off;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_is_unicore <= 1'h0;
    end else begin
      exe_reg_uops_2_is_unicore <= REG_5_is_unicore;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_shift <= 3'h0;
    end else begin
      exe_reg_uops_2_shift <= REG_5_shift;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_lrs3_rtype <= 2'h0;
    end else begin
      exe_reg_uops_2_lrs3_rtype <= REG_5_lrs3_rtype;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_rflag <= 1'h0;
    end else begin
      exe_reg_uops_2_rflag <= REG_5_rflag;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_wflag <= 1'h0;
    end else begin
      exe_reg_uops_2_wflag <= REG_5_wflag;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_prflag <= 4'h0;
    end else begin
      exe_reg_uops_2_prflag <= REG_5_prflag;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_pwflag <= 4'h0;
    end else begin
      exe_reg_uops_2_pwflag <= REG_5_pwflag;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_pflag_busy <= 1'h0;
    end else begin
      exe_reg_uops_2_pflag_busy <= REG_5_pflag_busy;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_stale_pflag <= 4'h0;
    end else begin
      exe_reg_uops_2_stale_pflag <= REG_5_stale_pflag;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_op1_sel <= 4'h0;
    end else begin
      exe_reg_uops_2_op1_sel <= REG_5_op1_sel;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_op2_sel <= 4'h0;
    end else begin
      exe_reg_uops_2_op2_sel <= REG_5_op2_sel;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_split_num <= 6'h0;
    end else begin
      exe_reg_uops_2_split_num <= REG_5_split_num;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_self_index <= 6'h0;
    end else begin
      exe_reg_uops_2_self_index <= REG_5_self_index;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_rob_inst_idx <= 6'h0;
    end else begin
      exe_reg_uops_2_rob_inst_idx <= REG_5_rob_inst_idx;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_address_num <= 6'h0;
    end else begin
      exe_reg_uops_2_address_num <= REG_5_address_num;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_uopc <= 7'h0;
    end else begin
      exe_reg_uops_2_uopc <= REG_5_uopc;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_inst <= 32'h0;
    end else begin
      exe_reg_uops_2_inst <= REG_5_inst;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_debug_inst <= 32'h0;
    end else begin
      exe_reg_uops_2_debug_inst <= REG_5_debug_inst;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_is_rvc <= 1'h0;
    end else begin
      exe_reg_uops_2_is_rvc <= REG_5_is_rvc;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_debug_pc <= 40'h0;
    end else begin
      exe_reg_uops_2_debug_pc <= REG_5_debug_pc;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_iq_type <= 3'h0;
    end else begin
      exe_reg_uops_2_iq_type <= REG_5_iq_type;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_fu_code <= 10'h0;
    end else begin
      exe_reg_uops_2_fu_code <= REG_5_fu_code;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_ctrl_br_type <= 4'h0;
    end else begin
      exe_reg_uops_2_ctrl_br_type <= REG_5_ctrl_br_type;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_ctrl_op1_sel <= 2'h0;
    end else begin
      exe_reg_uops_2_ctrl_op1_sel <= REG_5_ctrl_op1_sel;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_ctrl_op2_sel <= 3'h0;
    end else begin
      exe_reg_uops_2_ctrl_op2_sel <= REG_5_ctrl_op2_sel;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_ctrl_imm_sel <= 3'h0;
    end else begin
      exe_reg_uops_2_ctrl_imm_sel <= REG_5_ctrl_imm_sel;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_ctrl_op_fcn <= 4'h0;
    end else begin
      exe_reg_uops_2_ctrl_op_fcn <= REG_5_ctrl_op_fcn;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_ctrl_fcn_dw <= 1'h0;
    end else begin
      exe_reg_uops_2_ctrl_fcn_dw <= REG_5_ctrl_fcn_dw;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_ctrl_csr_cmd <= 3'h0;
    end else begin
      exe_reg_uops_2_ctrl_csr_cmd <= REG_5_ctrl_csr_cmd;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_ctrl_is_load <= 1'h0;
    end else begin
      exe_reg_uops_2_ctrl_is_load <= REG_5_ctrl_is_load;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_ctrl_is_sta <= 1'h0;
    end else begin
      exe_reg_uops_2_ctrl_is_sta <= REG_5_ctrl_is_sta;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_ctrl_is_std <= 1'h0;
    end else begin
      exe_reg_uops_2_ctrl_is_std <= REG_5_ctrl_is_std;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_ctrl_op3_sel <= 2'h0;
    end else begin
      exe_reg_uops_2_ctrl_op3_sel <= REG_5_ctrl_op3_sel;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_iw_state <= 2'h0;
    end else begin
      exe_reg_uops_2_iw_state <= REG_5_iw_state;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_iw_p1_poisoned <= 1'h0;
    end else begin
      exe_reg_uops_2_iw_p1_poisoned <= REG_5_iw_p1_poisoned;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_iw_p2_poisoned <= 1'h0;
    end else begin
      exe_reg_uops_2_iw_p2_poisoned <= REG_5_iw_p2_poisoned;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_is_br <= 1'h0;
    end else begin
      exe_reg_uops_2_is_br <= REG_5_is_br;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_is_jalr <= 1'h0;
    end else begin
      exe_reg_uops_2_is_jalr <= REG_5_is_jalr;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_is_jal <= 1'h0;
    end else begin
      exe_reg_uops_2_is_jal <= REG_5_is_jal;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_is_sfb <= 1'h0;
    end else begin
      exe_reg_uops_2_is_sfb <= REG_5_is_sfb;
    end
    exe_reg_uops_2_br_mask <= REG_5_br_mask & _T_4; // @[util.scala 142:25]
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_br_tag <= 4'h0;
    end else begin
      exe_reg_uops_2_br_tag <= REG_5_br_tag;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_ftq_idx <= 5'h0;
    end else begin
      exe_reg_uops_2_ftq_idx <= REG_5_ftq_idx;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_edge_inst <= 1'h0;
    end else begin
      exe_reg_uops_2_edge_inst <= REG_5_edge_inst;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_pc_lob <= 6'h0;
    end else begin
      exe_reg_uops_2_pc_lob <= REG_5_pc_lob;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_taken <= 1'h0;
    end else begin
      exe_reg_uops_2_taken <= REG_5_taken;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_imm_packed <= 20'h0;
    end else begin
      exe_reg_uops_2_imm_packed <= REG_5_imm_packed;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_csr_addr <= 12'h0;
    end else begin
      exe_reg_uops_2_csr_addr <= REG_5_csr_addr;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_rob_idx <= 6'h0;
    end else begin
      exe_reg_uops_2_rob_idx <= REG_5_rob_idx;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_ldq_idx <= 5'h0;
    end else begin
      exe_reg_uops_2_ldq_idx <= REG_5_ldq_idx;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_stq_idx <= 5'h0;
    end else begin
      exe_reg_uops_2_stq_idx <= REG_5_stq_idx;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_rxq_idx <= 2'h0;
    end else begin
      exe_reg_uops_2_rxq_idx <= REG_5_rxq_idx;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_pdst <= 7'h0;
    end else begin
      exe_reg_uops_2_pdst <= REG_5_pdst;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_prs1 <= 7'h0;
    end else begin
      exe_reg_uops_2_prs1 <= REG_5_prs1;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_prs2 <= 7'h0;
    end else begin
      exe_reg_uops_2_prs2 <= REG_5_prs2;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_prs3 <= 7'h0;
    end else begin
      exe_reg_uops_2_prs3 <= REG_5_prs3;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_ppred <= 5'h0;
    end else begin
      exe_reg_uops_2_ppred <= REG_5_ppred;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_prs1_busy <= 1'h0;
    end else begin
      exe_reg_uops_2_prs1_busy <= REG_5_prs1_busy;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_prs2_busy <= 1'h0;
    end else begin
      exe_reg_uops_2_prs2_busy <= REG_5_prs2_busy;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_prs3_busy <= 1'h0;
    end else begin
      exe_reg_uops_2_prs3_busy <= REG_5_prs3_busy;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_ppred_busy <= 1'h0;
    end else begin
      exe_reg_uops_2_ppred_busy <= REG_5_ppred_busy;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_stale_pdst <= 7'h0;
    end else begin
      exe_reg_uops_2_stale_pdst <= REG_5_stale_pdst;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_exception <= 1'h0;
    end else begin
      exe_reg_uops_2_exception <= REG_5_exception;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_exc_cause <= 64'h0;
    end else begin
      exe_reg_uops_2_exc_cause <= REG_5_exc_cause;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_bypassable <= 1'h0;
    end else begin
      exe_reg_uops_2_bypassable <= REG_5_bypassable;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_mem_cmd <= 5'h0;
    end else begin
      exe_reg_uops_2_mem_cmd <= REG_5_mem_cmd;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_mem_size <= 2'h0;
    end else begin
      exe_reg_uops_2_mem_size <= REG_5_mem_size;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_mem_signed <= 1'h0;
    end else begin
      exe_reg_uops_2_mem_signed <= REG_5_mem_signed;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_is_fence <= 1'h0;
    end else begin
      exe_reg_uops_2_is_fence <= REG_5_is_fence;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_is_fencei <= 1'h0;
    end else begin
      exe_reg_uops_2_is_fencei <= REG_5_is_fencei;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_is_amo <= 1'h0;
    end else begin
      exe_reg_uops_2_is_amo <= REG_5_is_amo;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_uses_ldq <= 1'h0;
    end else begin
      exe_reg_uops_2_uses_ldq <= REG_5_uses_ldq;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_uses_stq <= 1'h0;
    end else begin
      exe_reg_uops_2_uses_stq <= REG_5_uses_stq;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_is_sys_pc2epc <= 1'h0;
    end else begin
      exe_reg_uops_2_is_sys_pc2epc <= REG_5_is_sys_pc2epc;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_is_unique <= 1'h0;
    end else begin
      exe_reg_uops_2_is_unique <= REG_5_is_unique;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_flush_on_commit <= 1'h0;
    end else begin
      exe_reg_uops_2_flush_on_commit <= REG_5_flush_on_commit;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_ldst_is_rs1 <= 1'h0;
    end else begin
      exe_reg_uops_2_ldst_is_rs1 <= REG_5_ldst_is_rs1;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_ldst <= 6'h0;
    end else begin
      exe_reg_uops_2_ldst <= REG_5_ldst;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_lrs1 <= 6'h0;
    end else begin
      exe_reg_uops_2_lrs1 <= REG_5_lrs1;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_lrs2 <= 6'h0;
    end else begin
      exe_reg_uops_2_lrs2 <= REG_5_lrs2;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_lrs3 <= 6'h0;
    end else begin
      exe_reg_uops_2_lrs3 <= REG_5_lrs3;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_ldst_val <= 1'h0;
    end else begin
      exe_reg_uops_2_ldst_val <= REG_5_ldst_val;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_dst_rtype <= 2'h2;
    end else begin
      exe_reg_uops_2_dst_rtype <= REG_5_dst_rtype;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_lrs1_rtype <= 2'h0;
    end else begin
      exe_reg_uops_2_lrs1_rtype <= REG_5_lrs1_rtype;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_lrs2_rtype <= 2'h0;
    end else begin
      exe_reg_uops_2_lrs2_rtype <= REG_5_lrs2_rtype;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_frs3_en <= 1'h0;
    end else begin
      exe_reg_uops_2_frs3_en <= REG_5_frs3_en;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_fp_val <= 1'h0;
    end else begin
      exe_reg_uops_2_fp_val <= REG_5_fp_val;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_fp_single <= 1'h0;
    end else begin
      exe_reg_uops_2_fp_single <= REG_5_fp_single;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_xcpt_pf_if <= 1'h0;
    end else begin
      exe_reg_uops_2_xcpt_pf_if <= REG_5_xcpt_pf_if;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_xcpt_ae_if <= 1'h0;
    end else begin
      exe_reg_uops_2_xcpt_ae_if <= REG_5_xcpt_ae_if;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_xcpt_ma_if <= 1'h0;
    end else begin
      exe_reg_uops_2_xcpt_ma_if <= REG_5_xcpt_ma_if;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_bp_debug_if <= 1'h0;
    end else begin
      exe_reg_uops_2_bp_debug_if <= REG_5_bp_debug_if;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_bp_xcpt_if <= 1'h0;
    end else begin
      exe_reg_uops_2_bp_xcpt_if <= REG_5_bp_xcpt_if;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_debug_fsrc <= 2'h0;
    end else begin
      exe_reg_uops_2_debug_fsrc <= REG_5_debug_fsrc;
    end
    if (_T_76) begin // @[register-read.scala 149:29]
      exe_reg_uops_2_debug_tsrc <= 2'h0;
    end else begin
      exe_reg_uops_2_debug_tsrc <= REG_5_debug_tsrc;
    end
    if (_T_90) begin // @[Mux.scala 98:16]
      exe_reg_rs1_data_0 <= io_bypass_0_bits_data;
    end else if (_T_126) begin // @[Mux.scala 98:16]
      exe_reg_rs1_data_0 <= io_bypass_1_bits_data;
    end else if (_T_162) begin // @[Mux.scala 98:16]
      exe_reg_rs1_data_0 <= io_bypass_2_bits_data;
    end else if (_T_198) begin // @[Mux.scala 98:16]
      exe_reg_rs1_data_0 <= io_bypass_3_bits_data;
    end else begin
      exe_reg_rs1_data_0 <= rrd_rs1_data_0;
    end
    if (_T_269) begin // @[Mux.scala 98:16]
      exe_reg_rs1_data_1 <= io_bypass_0_bits_data;
    end else if (_T_305) begin // @[Mux.scala 98:16]
      exe_reg_rs1_data_1 <= io_bypass_1_bits_data;
    end else if (_T_341) begin // @[Mux.scala 98:16]
      exe_reg_rs1_data_1 <= io_bypass_2_bits_data;
    end else if (_T_377) begin // @[Mux.scala 98:16]
      exe_reg_rs1_data_1 <= io_bypass_3_bits_data;
    end else begin
      exe_reg_rs1_data_1 <= rrd_rs1_data_1;
    end
    if (_T_448) begin // @[Mux.scala 98:16]
      exe_reg_rs1_data_2 <= io_bypass_0_bits_data;
    end else if (_T_484) begin // @[Mux.scala 98:16]
      exe_reg_rs1_data_2 <= io_bypass_1_bits_data;
    end else if (_T_520) begin // @[Mux.scala 98:16]
      exe_reg_rs1_data_2 <= io_bypass_2_bits_data;
    end else if (_T_556) begin // @[Mux.scala 98:16]
      exe_reg_rs1_data_2 <= io_bypass_3_bits_data;
    end else begin
      exe_reg_rs1_data_2 <= rrd_rs1_data_2;
    end
    if (_T_100) begin // @[Mux.scala 98:16]
      exe_reg_rs2_data_0 <= io_bypass_0_bits_data;
    end else if (_T_136) begin // @[Mux.scala 98:16]
      exe_reg_rs2_data_0 <= io_bypass_1_bits_data;
    end else if (_T_172) begin // @[Mux.scala 98:16]
      exe_reg_rs2_data_0 <= io_bypass_2_bits_data;
    end else if (_T_208) begin // @[Mux.scala 98:16]
      exe_reg_rs2_data_0 <= io_bypass_3_bits_data;
    end else begin
      exe_reg_rs2_data_0 <= rrd_rs2_data_0;
    end
    if (_T_279) begin // @[Mux.scala 98:16]
      exe_reg_rs2_data_1 <= io_bypass_0_bits_data;
    end else if (_T_315) begin // @[Mux.scala 98:16]
      exe_reg_rs2_data_1 <= io_bypass_1_bits_data;
    end else if (_T_351) begin // @[Mux.scala 98:16]
      exe_reg_rs2_data_1 <= io_bypass_2_bits_data;
    end else if (_T_387) begin // @[Mux.scala 98:16]
      exe_reg_rs2_data_1 <= io_bypass_3_bits_data;
    end else begin
      exe_reg_rs2_data_1 <= rrd_rs2_data_1;
    end
    if (_T_458) begin // @[Mux.scala 98:16]
      exe_reg_rs2_data_2 <= io_bypass_0_bits_data;
    end else if (_T_494) begin // @[Mux.scala 98:16]
      exe_reg_rs2_data_2 <= io_bypass_1_bits_data;
    end else if (_T_530) begin // @[Mux.scala 98:16]
      exe_reg_rs2_data_2 <= io_bypass_2_bits_data;
    end else if (_T_566) begin // @[Mux.scala 98:16]
      exe_reg_rs2_data_2 <= io_bypass_3_bits_data;
    end else begin
      exe_reg_rs2_data_2 <= rrd_rs2_data_2;
    end
    if (_T_110) begin // @[Mux.scala 98:16]
      exe_reg_rs3_data_0 <= io_bypass_0_bits_data;
    end else if (_T_146) begin // @[Mux.scala 98:16]
      exe_reg_rs3_data_0 <= io_bypass_1_bits_data;
    end else if (_T_182) begin // @[Mux.scala 98:16]
      exe_reg_rs3_data_0 <= io_bypass_2_bits_data;
    end else if (_T_218) begin // @[Mux.scala 98:16]
      exe_reg_rs3_data_0 <= io_bypass_3_bits_data;
    end else begin
      exe_reg_rs3_data_0 <= rrd_rs3_data_0;
    end
    if (_T_289) begin // @[Mux.scala 98:16]
      exe_reg_rs3_data_1 <= io_bypass_0_bits_data;
    end else if (_T_325) begin // @[Mux.scala 98:16]
      exe_reg_rs3_data_1 <= io_bypass_1_bits_data;
    end else if (_T_361) begin // @[Mux.scala 98:16]
      exe_reg_rs3_data_1 <= io_bypass_2_bits_data;
    end else if (_T_397) begin // @[Mux.scala 98:16]
      exe_reg_rs3_data_1 <= io_bypass_3_bits_data;
    end else begin
      exe_reg_rs3_data_1 <= rrd_rs3_data_1;
    end
    if (_T_468) begin // @[Mux.scala 98:16]
      exe_reg_rs3_data_2 <= io_bypass_0_bits_data;
    end else if (_T_504) begin // @[Mux.scala 98:16]
      exe_reg_rs3_data_2 <= io_bypass_1_bits_data;
    end else if (_T_540) begin // @[Mux.scala 98:16]
      exe_reg_rs3_data_2 <= io_bypass_2_bits_data;
    end else if (_T_576) begin // @[Mux.scala 98:16]
      exe_reg_rs3_data_2 <= io_bypass_3_bits_data;
    end else begin
      exe_reg_rs3_data_2 <= rrd_rs3_data_2;
    end
    if (_T_116) begin // @[Mux.scala 98:16]
      exe_reg_flag_data_0 <= io_bypass_0_bits_flagdata;
    end else if (_T_152) begin // @[Mux.scala 98:16]
      exe_reg_flag_data_0 <= io_bypass_1_bits_flagdata;
    end else if (_T_188) begin // @[Mux.scala 98:16]
      exe_reg_flag_data_0 <= io_bypass_2_bits_flagdata;
    end else if (_T_224) begin // @[Mux.scala 98:16]
      exe_reg_flag_data_0 <= io_bypass_3_bits_flagdata;
    end else begin
      exe_reg_flag_data_0 <= rrd_flag_data_0;
    end
    if (_T_295) begin // @[Mux.scala 98:16]
      exe_reg_flag_data_1 <= io_bypass_0_bits_flagdata;
    end else if (_T_331) begin // @[Mux.scala 98:16]
      exe_reg_flag_data_1 <= io_bypass_1_bits_flagdata;
    end else if (_T_367) begin // @[Mux.scala 98:16]
      exe_reg_flag_data_1 <= io_bypass_2_bits_flagdata;
    end else if (_T_403) begin // @[Mux.scala 98:16]
      exe_reg_flag_data_1 <= io_bypass_3_bits_flagdata;
    end else begin
      exe_reg_flag_data_1 <= rrd_flag_data_1;
    end
    if (_T_474) begin // @[Mux.scala 98:16]
      exe_reg_flag_data_2 <= io_bypass_0_bits_flagdata;
    end else if (_T_510) begin // @[Mux.scala 98:16]
      exe_reg_flag_data_2 <= io_bypass_1_bits_flagdata;
    end else if (_T_546) begin // @[Mux.scala 98:16]
      exe_reg_flag_data_2 <= io_bypass_2_bits_flagdata;
    end else if (_T_582) begin // @[Mux.scala 98:16]
      exe_reg_flag_data_2 <= io_bypass_3_bits_flagdata;
    end else begin
      exe_reg_flag_data_2 <= rrd_flag_data_2;
    end
    REG <= RegisterReadDecode_io_rrd_valid & _T_2; // @[register-read.scala 90:59]
    REG_1_switch <= RegisterReadDecode_io_rrd_uop_switch; // @[register-read.scala 92:29]
    REG_1_switch_off <= RegisterReadDecode_io_rrd_uop_switch_off; // @[register-read.scala 92:29]
    REG_1_is_unicore <= RegisterReadDecode_io_rrd_uop_is_unicore; // @[register-read.scala 92:29]
    REG_1_shift <= RegisterReadDecode_io_rrd_uop_shift; // @[register-read.scala 92:29]
    REG_1_lrs3_rtype <= RegisterReadDecode_io_rrd_uop_lrs3_rtype; // @[register-read.scala 92:29]
    REG_1_rflag <= RegisterReadDecode_io_rrd_uop_rflag; // @[register-read.scala 92:29]
    REG_1_wflag <= RegisterReadDecode_io_rrd_uop_wflag; // @[register-read.scala 92:29]
    REG_1_prflag <= RegisterReadDecode_io_rrd_uop_prflag; // @[register-read.scala 92:29]
    REG_1_pwflag <= RegisterReadDecode_io_rrd_uop_pwflag; // @[register-read.scala 92:29]
    REG_1_pflag_busy <= RegisterReadDecode_io_rrd_uop_pflag_busy; // @[register-read.scala 92:29]
    REG_1_stale_pflag <= RegisterReadDecode_io_rrd_uop_stale_pflag; // @[register-read.scala 92:29]
    REG_1_op1_sel <= RegisterReadDecode_io_rrd_uop_op1_sel; // @[register-read.scala 92:29]
    REG_1_op2_sel <= RegisterReadDecode_io_rrd_uop_op2_sel; // @[register-read.scala 92:29]
    REG_1_split_num <= RegisterReadDecode_io_rrd_uop_split_num; // @[register-read.scala 92:29]
    REG_1_self_index <= RegisterReadDecode_io_rrd_uop_self_index; // @[register-read.scala 92:29]
    REG_1_rob_inst_idx <= RegisterReadDecode_io_rrd_uop_rob_inst_idx; // @[register-read.scala 92:29]
    REG_1_address_num <= RegisterReadDecode_io_rrd_uop_address_num; // @[register-read.scala 92:29]
    REG_1_uopc <= RegisterReadDecode_io_rrd_uop_uopc; // @[register-read.scala 92:29]
    REG_1_inst <= RegisterReadDecode_io_rrd_uop_inst; // @[register-read.scala 92:29]
    REG_1_debug_inst <= RegisterReadDecode_io_rrd_uop_debug_inst; // @[register-read.scala 92:29]
    REG_1_is_rvc <= RegisterReadDecode_io_rrd_uop_is_rvc; // @[register-read.scala 92:29]
    REG_1_debug_pc <= RegisterReadDecode_io_rrd_uop_debug_pc; // @[register-read.scala 92:29]
    REG_1_iq_type <= RegisterReadDecode_io_rrd_uop_iq_type; // @[register-read.scala 92:29]
    REG_1_fu_code <= RegisterReadDecode_io_rrd_uop_fu_code; // @[register-read.scala 92:29]
    REG_1_ctrl_br_type <= RegisterReadDecode_io_rrd_uop_ctrl_br_type; // @[register-read.scala 92:29]
    REG_1_ctrl_op1_sel <= RegisterReadDecode_io_rrd_uop_ctrl_op1_sel; // @[register-read.scala 92:29]
    REG_1_ctrl_op2_sel <= RegisterReadDecode_io_rrd_uop_ctrl_op2_sel; // @[register-read.scala 92:29]
    REG_1_ctrl_imm_sel <= RegisterReadDecode_io_rrd_uop_ctrl_imm_sel; // @[register-read.scala 92:29]
    REG_1_ctrl_op_fcn <= RegisterReadDecode_io_rrd_uop_ctrl_op_fcn; // @[register-read.scala 92:29]
    REG_1_ctrl_fcn_dw <= RegisterReadDecode_io_rrd_uop_ctrl_fcn_dw; // @[register-read.scala 92:29]
    REG_1_ctrl_csr_cmd <= RegisterReadDecode_io_rrd_uop_ctrl_csr_cmd; // @[register-read.scala 92:29]
    REG_1_ctrl_is_load <= RegisterReadDecode_io_rrd_uop_ctrl_is_load; // @[register-read.scala 92:29]
    REG_1_ctrl_is_sta <= RegisterReadDecode_io_rrd_uop_ctrl_is_sta; // @[register-read.scala 92:29]
    REG_1_ctrl_is_std <= RegisterReadDecode_io_rrd_uop_ctrl_is_std; // @[register-read.scala 92:29]
    REG_1_ctrl_op3_sel <= RegisterReadDecode_io_rrd_uop_ctrl_op3_sel; // @[register-read.scala 92:29]
    REG_1_iw_state <= RegisterReadDecode_io_rrd_uop_iw_state; // @[register-read.scala 92:29]
    REG_1_iw_p1_poisoned <= RegisterReadDecode_io_rrd_uop_iw_p1_poisoned; // @[register-read.scala 92:29]
    REG_1_iw_p2_poisoned <= RegisterReadDecode_io_rrd_uop_iw_p2_poisoned; // @[register-read.scala 92:29]
    REG_1_is_br <= RegisterReadDecode_io_rrd_uop_is_br; // @[register-read.scala 92:29]
    REG_1_is_jalr <= RegisterReadDecode_io_rrd_uop_is_jalr; // @[register-read.scala 92:29]
    REG_1_is_jal <= RegisterReadDecode_io_rrd_uop_is_jal; // @[register-read.scala 92:29]
    REG_1_is_sfb <= RegisterReadDecode_io_rrd_uop_is_sfb; // @[register-read.scala 92:29]
    REG_1_br_mask <= RegisterReadDecode_io_rrd_uop_br_mask & _T_4; // @[util.scala 131:35]
    REG_1_br_tag <= RegisterReadDecode_io_rrd_uop_br_tag; // @[register-read.scala 92:29]
    REG_1_ftq_idx <= RegisterReadDecode_io_rrd_uop_ftq_idx; // @[register-read.scala 92:29]
    REG_1_edge_inst <= RegisterReadDecode_io_rrd_uop_edge_inst; // @[register-read.scala 92:29]
    REG_1_pc_lob <= RegisterReadDecode_io_rrd_uop_pc_lob; // @[register-read.scala 92:29]
    REG_1_taken <= RegisterReadDecode_io_rrd_uop_taken; // @[register-read.scala 92:29]
    REG_1_imm_packed <= RegisterReadDecode_io_rrd_uop_imm_packed; // @[register-read.scala 92:29]
    REG_1_csr_addr <= RegisterReadDecode_io_rrd_uop_csr_addr; // @[register-read.scala 92:29]
    REG_1_rob_idx <= RegisterReadDecode_io_rrd_uop_rob_idx; // @[register-read.scala 92:29]
    REG_1_ldq_idx <= RegisterReadDecode_io_rrd_uop_ldq_idx; // @[register-read.scala 92:29]
    REG_1_stq_idx <= RegisterReadDecode_io_rrd_uop_stq_idx; // @[register-read.scala 92:29]
    REG_1_rxq_idx <= RegisterReadDecode_io_rrd_uop_rxq_idx; // @[register-read.scala 92:29]
    REG_1_pdst <= RegisterReadDecode_io_rrd_uop_pdst; // @[register-read.scala 92:29]
    REG_1_prs1 <= RegisterReadDecode_io_rrd_uop_prs1; // @[register-read.scala 92:29]
    REG_1_prs2 <= RegisterReadDecode_io_rrd_uop_prs2; // @[register-read.scala 92:29]
    REG_1_prs3 <= RegisterReadDecode_io_rrd_uop_prs3; // @[register-read.scala 92:29]
    REG_1_ppred <= RegisterReadDecode_io_rrd_uop_ppred; // @[register-read.scala 92:29]
    REG_1_prs1_busy <= RegisterReadDecode_io_rrd_uop_prs1_busy; // @[register-read.scala 92:29]
    REG_1_prs2_busy <= RegisterReadDecode_io_rrd_uop_prs2_busy; // @[register-read.scala 92:29]
    REG_1_prs3_busy <= RegisterReadDecode_io_rrd_uop_prs3_busy; // @[register-read.scala 92:29]
    REG_1_ppred_busy <= RegisterReadDecode_io_rrd_uop_ppred_busy; // @[register-read.scala 92:29]
    REG_1_stale_pdst <= RegisterReadDecode_io_rrd_uop_stale_pdst; // @[register-read.scala 92:29]
    REG_1_exception <= RegisterReadDecode_io_rrd_uop_exception; // @[register-read.scala 92:29]
    REG_1_exc_cause <= RegisterReadDecode_io_rrd_uop_exc_cause; // @[register-read.scala 92:29]
    REG_1_bypassable <= RegisterReadDecode_io_rrd_uop_bypassable; // @[register-read.scala 92:29]
    REG_1_mem_cmd <= RegisterReadDecode_io_rrd_uop_mem_cmd; // @[register-read.scala 92:29]
    REG_1_mem_size <= RegisterReadDecode_io_rrd_uop_mem_size; // @[register-read.scala 92:29]
    REG_1_mem_signed <= RegisterReadDecode_io_rrd_uop_mem_signed; // @[register-read.scala 92:29]
    REG_1_is_fence <= RegisterReadDecode_io_rrd_uop_is_fence; // @[register-read.scala 92:29]
    REG_1_is_fencei <= RegisterReadDecode_io_rrd_uop_is_fencei; // @[register-read.scala 92:29]
    REG_1_is_amo <= RegisterReadDecode_io_rrd_uop_is_amo; // @[register-read.scala 92:29]
    REG_1_uses_ldq <= RegisterReadDecode_io_rrd_uop_uses_ldq; // @[register-read.scala 92:29]
    REG_1_uses_stq <= RegisterReadDecode_io_rrd_uop_uses_stq; // @[register-read.scala 92:29]
    REG_1_is_sys_pc2epc <= RegisterReadDecode_io_rrd_uop_is_sys_pc2epc; // @[register-read.scala 92:29]
    REG_1_is_unique <= RegisterReadDecode_io_rrd_uop_is_unique; // @[register-read.scala 92:29]
    REG_1_flush_on_commit <= RegisterReadDecode_io_rrd_uop_flush_on_commit; // @[register-read.scala 92:29]
    REG_1_ldst_is_rs1 <= RegisterReadDecode_io_rrd_uop_ldst_is_rs1; // @[register-read.scala 92:29]
    REG_1_ldst <= RegisterReadDecode_io_rrd_uop_ldst; // @[register-read.scala 92:29]
    REG_1_lrs1 <= RegisterReadDecode_io_rrd_uop_lrs1; // @[register-read.scala 92:29]
    REG_1_lrs2 <= RegisterReadDecode_io_rrd_uop_lrs2; // @[register-read.scala 92:29]
    REG_1_lrs3 <= RegisterReadDecode_io_rrd_uop_lrs3; // @[register-read.scala 92:29]
    REG_1_ldst_val <= RegisterReadDecode_io_rrd_uop_ldst_val; // @[register-read.scala 92:29]
    REG_1_dst_rtype <= RegisterReadDecode_io_rrd_uop_dst_rtype; // @[register-read.scala 92:29]
    REG_1_lrs1_rtype <= RegisterReadDecode_io_rrd_uop_lrs1_rtype; // @[register-read.scala 92:29]
    REG_1_lrs2_rtype <= RegisterReadDecode_io_rrd_uop_lrs2_rtype; // @[register-read.scala 92:29]
    REG_1_frs3_en <= RegisterReadDecode_io_rrd_uop_frs3_en; // @[register-read.scala 92:29]
    REG_1_fp_val <= RegisterReadDecode_io_rrd_uop_fp_val; // @[register-read.scala 92:29]
    REG_1_fp_single <= RegisterReadDecode_io_rrd_uop_fp_single; // @[register-read.scala 92:29]
    REG_1_xcpt_pf_if <= RegisterReadDecode_io_rrd_uop_xcpt_pf_if; // @[register-read.scala 92:29]
    REG_1_xcpt_ae_if <= RegisterReadDecode_io_rrd_uop_xcpt_ae_if; // @[register-read.scala 92:29]
    REG_1_xcpt_ma_if <= RegisterReadDecode_io_rrd_uop_xcpt_ma_if; // @[register-read.scala 92:29]
    REG_1_bp_debug_if <= RegisterReadDecode_io_rrd_uop_bp_debug_if; // @[register-read.scala 92:29]
    REG_1_bp_xcpt_if <= RegisterReadDecode_io_rrd_uop_bp_xcpt_if; // @[register-read.scala 92:29]
    REG_1_debug_fsrc <= RegisterReadDecode_io_rrd_uop_debug_fsrc; // @[register-read.scala 92:29]
    REG_1_debug_tsrc <= RegisterReadDecode_io_rrd_uop_debug_tsrc; // @[register-read.scala 92:29]
    REG_2 <= RegisterReadDecode_1_io_rrd_valid & _T_8; // @[register-read.scala 90:59]
    REG_3_switch <= RegisterReadDecode_1_io_rrd_uop_switch; // @[register-read.scala 92:29]
    REG_3_switch_off <= RegisterReadDecode_1_io_rrd_uop_switch_off; // @[register-read.scala 92:29]
    REG_3_is_unicore <= RegisterReadDecode_1_io_rrd_uop_is_unicore; // @[register-read.scala 92:29]
    REG_3_shift <= RegisterReadDecode_1_io_rrd_uop_shift; // @[register-read.scala 92:29]
    REG_3_lrs3_rtype <= RegisterReadDecode_1_io_rrd_uop_lrs3_rtype; // @[register-read.scala 92:29]
    REG_3_rflag <= RegisterReadDecode_1_io_rrd_uop_rflag; // @[register-read.scala 92:29]
    REG_3_wflag <= RegisterReadDecode_1_io_rrd_uop_wflag; // @[register-read.scala 92:29]
    REG_3_prflag <= RegisterReadDecode_1_io_rrd_uop_prflag; // @[register-read.scala 92:29]
    REG_3_pwflag <= RegisterReadDecode_1_io_rrd_uop_pwflag; // @[register-read.scala 92:29]
    REG_3_pflag_busy <= RegisterReadDecode_1_io_rrd_uop_pflag_busy; // @[register-read.scala 92:29]
    REG_3_stale_pflag <= RegisterReadDecode_1_io_rrd_uop_stale_pflag; // @[register-read.scala 92:29]
    REG_3_op1_sel <= RegisterReadDecode_1_io_rrd_uop_op1_sel; // @[register-read.scala 92:29]
    REG_3_op2_sel <= RegisterReadDecode_1_io_rrd_uop_op2_sel; // @[register-read.scala 92:29]
    REG_3_split_num <= RegisterReadDecode_1_io_rrd_uop_split_num; // @[register-read.scala 92:29]
    REG_3_self_index <= RegisterReadDecode_1_io_rrd_uop_self_index; // @[register-read.scala 92:29]
    REG_3_rob_inst_idx <= RegisterReadDecode_1_io_rrd_uop_rob_inst_idx; // @[register-read.scala 92:29]
    REG_3_address_num <= RegisterReadDecode_1_io_rrd_uop_address_num; // @[register-read.scala 92:29]
    REG_3_uopc <= RegisterReadDecode_1_io_rrd_uop_uopc; // @[register-read.scala 92:29]
    REG_3_inst <= RegisterReadDecode_1_io_rrd_uop_inst; // @[register-read.scala 92:29]
    REG_3_debug_inst <= RegisterReadDecode_1_io_rrd_uop_debug_inst; // @[register-read.scala 92:29]
    REG_3_is_rvc <= RegisterReadDecode_1_io_rrd_uop_is_rvc; // @[register-read.scala 92:29]
    REG_3_debug_pc <= RegisterReadDecode_1_io_rrd_uop_debug_pc; // @[register-read.scala 92:29]
    REG_3_iq_type <= RegisterReadDecode_1_io_rrd_uop_iq_type; // @[register-read.scala 92:29]
    REG_3_fu_code <= RegisterReadDecode_1_io_rrd_uop_fu_code; // @[register-read.scala 92:29]
    REG_3_ctrl_br_type <= RegisterReadDecode_1_io_rrd_uop_ctrl_br_type; // @[register-read.scala 92:29]
    REG_3_ctrl_op1_sel <= RegisterReadDecode_1_io_rrd_uop_ctrl_op1_sel; // @[register-read.scala 92:29]
    REG_3_ctrl_op2_sel <= RegisterReadDecode_1_io_rrd_uop_ctrl_op2_sel; // @[register-read.scala 92:29]
    REG_3_ctrl_imm_sel <= RegisterReadDecode_1_io_rrd_uop_ctrl_imm_sel; // @[register-read.scala 92:29]
    REG_3_ctrl_op_fcn <= RegisterReadDecode_1_io_rrd_uop_ctrl_op_fcn; // @[register-read.scala 92:29]
    REG_3_ctrl_fcn_dw <= RegisterReadDecode_1_io_rrd_uop_ctrl_fcn_dw; // @[register-read.scala 92:29]
    REG_3_ctrl_csr_cmd <= RegisterReadDecode_1_io_rrd_uop_ctrl_csr_cmd; // @[register-read.scala 92:29]
    REG_3_ctrl_is_load <= RegisterReadDecode_1_io_rrd_uop_ctrl_is_load; // @[register-read.scala 92:29]
    REG_3_ctrl_is_sta <= RegisterReadDecode_1_io_rrd_uop_ctrl_is_sta; // @[register-read.scala 92:29]
    REG_3_ctrl_is_std <= RegisterReadDecode_1_io_rrd_uop_ctrl_is_std; // @[register-read.scala 92:29]
    REG_3_ctrl_op3_sel <= RegisterReadDecode_1_io_rrd_uop_ctrl_op3_sel; // @[register-read.scala 92:29]
    REG_3_iw_state <= RegisterReadDecode_1_io_rrd_uop_iw_state; // @[register-read.scala 92:29]
    REG_3_iw_p1_poisoned <= RegisterReadDecode_1_io_rrd_uop_iw_p1_poisoned; // @[register-read.scala 92:29]
    REG_3_iw_p2_poisoned <= RegisterReadDecode_1_io_rrd_uop_iw_p2_poisoned; // @[register-read.scala 92:29]
    REG_3_is_br <= RegisterReadDecode_1_io_rrd_uop_is_br; // @[register-read.scala 92:29]
    REG_3_is_jalr <= RegisterReadDecode_1_io_rrd_uop_is_jalr; // @[register-read.scala 92:29]
    REG_3_is_jal <= RegisterReadDecode_1_io_rrd_uop_is_jal; // @[register-read.scala 92:29]
    REG_3_is_sfb <= RegisterReadDecode_1_io_rrd_uop_is_sfb; // @[register-read.scala 92:29]
    REG_3_br_mask <= RegisterReadDecode_1_io_rrd_uop_br_mask & _T_4; // @[util.scala 131:35]
    REG_3_br_tag <= RegisterReadDecode_1_io_rrd_uop_br_tag; // @[register-read.scala 92:29]
    REG_3_ftq_idx <= RegisterReadDecode_1_io_rrd_uop_ftq_idx; // @[register-read.scala 92:29]
    REG_3_edge_inst <= RegisterReadDecode_1_io_rrd_uop_edge_inst; // @[register-read.scala 92:29]
    REG_3_pc_lob <= RegisterReadDecode_1_io_rrd_uop_pc_lob; // @[register-read.scala 92:29]
    REG_3_taken <= RegisterReadDecode_1_io_rrd_uop_taken; // @[register-read.scala 92:29]
    REG_3_imm_packed <= RegisterReadDecode_1_io_rrd_uop_imm_packed; // @[register-read.scala 92:29]
    REG_3_csr_addr <= RegisterReadDecode_1_io_rrd_uop_csr_addr; // @[register-read.scala 92:29]
    REG_3_rob_idx <= RegisterReadDecode_1_io_rrd_uop_rob_idx; // @[register-read.scala 92:29]
    REG_3_ldq_idx <= RegisterReadDecode_1_io_rrd_uop_ldq_idx; // @[register-read.scala 92:29]
    REG_3_stq_idx <= RegisterReadDecode_1_io_rrd_uop_stq_idx; // @[register-read.scala 92:29]
    REG_3_rxq_idx <= RegisterReadDecode_1_io_rrd_uop_rxq_idx; // @[register-read.scala 92:29]
    REG_3_pdst <= RegisterReadDecode_1_io_rrd_uop_pdst; // @[register-read.scala 92:29]
    REG_3_prs1 <= RegisterReadDecode_1_io_rrd_uop_prs1; // @[register-read.scala 92:29]
    REG_3_prs2 <= RegisterReadDecode_1_io_rrd_uop_prs2; // @[register-read.scala 92:29]
    REG_3_prs3 <= RegisterReadDecode_1_io_rrd_uop_prs3; // @[register-read.scala 92:29]
    REG_3_ppred <= RegisterReadDecode_1_io_rrd_uop_ppred; // @[register-read.scala 92:29]
    REG_3_prs1_busy <= RegisterReadDecode_1_io_rrd_uop_prs1_busy; // @[register-read.scala 92:29]
    REG_3_prs2_busy <= RegisterReadDecode_1_io_rrd_uop_prs2_busy; // @[register-read.scala 92:29]
    REG_3_prs3_busy <= RegisterReadDecode_1_io_rrd_uop_prs3_busy; // @[register-read.scala 92:29]
    REG_3_ppred_busy <= RegisterReadDecode_1_io_rrd_uop_ppred_busy; // @[register-read.scala 92:29]
    REG_3_stale_pdst <= RegisterReadDecode_1_io_rrd_uop_stale_pdst; // @[register-read.scala 92:29]
    REG_3_exception <= RegisterReadDecode_1_io_rrd_uop_exception; // @[register-read.scala 92:29]
    REG_3_exc_cause <= RegisterReadDecode_1_io_rrd_uop_exc_cause; // @[register-read.scala 92:29]
    REG_3_bypassable <= RegisterReadDecode_1_io_rrd_uop_bypassable; // @[register-read.scala 92:29]
    REG_3_mem_cmd <= RegisterReadDecode_1_io_rrd_uop_mem_cmd; // @[register-read.scala 92:29]
    REG_3_mem_size <= RegisterReadDecode_1_io_rrd_uop_mem_size; // @[register-read.scala 92:29]
    REG_3_mem_signed <= RegisterReadDecode_1_io_rrd_uop_mem_signed; // @[register-read.scala 92:29]
    REG_3_is_fence <= RegisterReadDecode_1_io_rrd_uop_is_fence; // @[register-read.scala 92:29]
    REG_3_is_fencei <= RegisterReadDecode_1_io_rrd_uop_is_fencei; // @[register-read.scala 92:29]
    REG_3_is_amo <= RegisterReadDecode_1_io_rrd_uop_is_amo; // @[register-read.scala 92:29]
    REG_3_uses_ldq <= RegisterReadDecode_1_io_rrd_uop_uses_ldq; // @[register-read.scala 92:29]
    REG_3_uses_stq <= RegisterReadDecode_1_io_rrd_uop_uses_stq; // @[register-read.scala 92:29]
    REG_3_is_sys_pc2epc <= RegisterReadDecode_1_io_rrd_uop_is_sys_pc2epc; // @[register-read.scala 92:29]
    REG_3_is_unique <= RegisterReadDecode_1_io_rrd_uop_is_unique; // @[register-read.scala 92:29]
    REG_3_flush_on_commit <= RegisterReadDecode_1_io_rrd_uop_flush_on_commit; // @[register-read.scala 92:29]
    REG_3_ldst_is_rs1 <= RegisterReadDecode_1_io_rrd_uop_ldst_is_rs1; // @[register-read.scala 92:29]
    REG_3_ldst <= RegisterReadDecode_1_io_rrd_uop_ldst; // @[register-read.scala 92:29]
    REG_3_lrs1 <= RegisterReadDecode_1_io_rrd_uop_lrs1; // @[register-read.scala 92:29]
    REG_3_lrs2 <= RegisterReadDecode_1_io_rrd_uop_lrs2; // @[register-read.scala 92:29]
    REG_3_lrs3 <= RegisterReadDecode_1_io_rrd_uop_lrs3; // @[register-read.scala 92:29]
    REG_3_ldst_val <= RegisterReadDecode_1_io_rrd_uop_ldst_val; // @[register-read.scala 92:29]
    REG_3_dst_rtype <= RegisterReadDecode_1_io_rrd_uop_dst_rtype; // @[register-read.scala 92:29]
    REG_3_lrs1_rtype <= RegisterReadDecode_1_io_rrd_uop_lrs1_rtype; // @[register-read.scala 92:29]
    REG_3_lrs2_rtype <= RegisterReadDecode_1_io_rrd_uop_lrs2_rtype; // @[register-read.scala 92:29]
    REG_3_frs3_en <= RegisterReadDecode_1_io_rrd_uop_frs3_en; // @[register-read.scala 92:29]
    REG_3_fp_val <= RegisterReadDecode_1_io_rrd_uop_fp_val; // @[register-read.scala 92:29]
    REG_3_fp_single <= RegisterReadDecode_1_io_rrd_uop_fp_single; // @[register-read.scala 92:29]
    REG_3_xcpt_pf_if <= RegisterReadDecode_1_io_rrd_uop_xcpt_pf_if; // @[register-read.scala 92:29]
    REG_3_xcpt_ae_if <= RegisterReadDecode_1_io_rrd_uop_xcpt_ae_if; // @[register-read.scala 92:29]
    REG_3_xcpt_ma_if <= RegisterReadDecode_1_io_rrd_uop_xcpt_ma_if; // @[register-read.scala 92:29]
    REG_3_bp_debug_if <= RegisterReadDecode_1_io_rrd_uop_bp_debug_if; // @[register-read.scala 92:29]
    REG_3_bp_xcpt_if <= RegisterReadDecode_1_io_rrd_uop_bp_xcpt_if; // @[register-read.scala 92:29]
    REG_3_debug_fsrc <= RegisterReadDecode_1_io_rrd_uop_debug_fsrc; // @[register-read.scala 92:29]
    REG_3_debug_tsrc <= RegisterReadDecode_1_io_rrd_uop_debug_tsrc; // @[register-read.scala 92:29]
    REG_4 <= RegisterReadDecode_2_io_rrd_valid & _T_14; // @[register-read.scala 90:59]
    REG_5_switch <= RegisterReadDecode_2_io_rrd_uop_switch; // @[register-read.scala 92:29]
    REG_5_switch_off <= RegisterReadDecode_2_io_rrd_uop_switch_off; // @[register-read.scala 92:29]
    REG_5_is_unicore <= RegisterReadDecode_2_io_rrd_uop_is_unicore; // @[register-read.scala 92:29]
    REG_5_shift <= RegisterReadDecode_2_io_rrd_uop_shift; // @[register-read.scala 92:29]
    REG_5_lrs3_rtype <= RegisterReadDecode_2_io_rrd_uop_lrs3_rtype; // @[register-read.scala 92:29]
    REG_5_rflag <= RegisterReadDecode_2_io_rrd_uop_rflag; // @[register-read.scala 92:29]
    REG_5_wflag <= RegisterReadDecode_2_io_rrd_uop_wflag; // @[register-read.scala 92:29]
    REG_5_prflag <= RegisterReadDecode_2_io_rrd_uop_prflag; // @[register-read.scala 92:29]
    REG_5_pwflag <= RegisterReadDecode_2_io_rrd_uop_pwflag; // @[register-read.scala 92:29]
    REG_5_pflag_busy <= RegisterReadDecode_2_io_rrd_uop_pflag_busy; // @[register-read.scala 92:29]
    REG_5_stale_pflag <= RegisterReadDecode_2_io_rrd_uop_stale_pflag; // @[register-read.scala 92:29]
    REG_5_op1_sel <= RegisterReadDecode_2_io_rrd_uop_op1_sel; // @[register-read.scala 92:29]
    REG_5_op2_sel <= RegisterReadDecode_2_io_rrd_uop_op2_sel; // @[register-read.scala 92:29]
    REG_5_split_num <= RegisterReadDecode_2_io_rrd_uop_split_num; // @[register-read.scala 92:29]
    REG_5_self_index <= RegisterReadDecode_2_io_rrd_uop_self_index; // @[register-read.scala 92:29]
    REG_5_rob_inst_idx <= RegisterReadDecode_2_io_rrd_uop_rob_inst_idx; // @[register-read.scala 92:29]
    REG_5_address_num <= RegisterReadDecode_2_io_rrd_uop_address_num; // @[register-read.scala 92:29]
    REG_5_uopc <= RegisterReadDecode_2_io_rrd_uop_uopc; // @[register-read.scala 92:29]
    REG_5_inst <= RegisterReadDecode_2_io_rrd_uop_inst; // @[register-read.scala 92:29]
    REG_5_debug_inst <= RegisterReadDecode_2_io_rrd_uop_debug_inst; // @[register-read.scala 92:29]
    REG_5_is_rvc <= RegisterReadDecode_2_io_rrd_uop_is_rvc; // @[register-read.scala 92:29]
    REG_5_debug_pc <= RegisterReadDecode_2_io_rrd_uop_debug_pc; // @[register-read.scala 92:29]
    REG_5_iq_type <= RegisterReadDecode_2_io_rrd_uop_iq_type; // @[register-read.scala 92:29]
    REG_5_fu_code <= RegisterReadDecode_2_io_rrd_uop_fu_code; // @[register-read.scala 92:29]
    REG_5_ctrl_br_type <= RegisterReadDecode_2_io_rrd_uop_ctrl_br_type; // @[register-read.scala 92:29]
    REG_5_ctrl_op1_sel <= RegisterReadDecode_2_io_rrd_uop_ctrl_op1_sel; // @[register-read.scala 92:29]
    REG_5_ctrl_op2_sel <= RegisterReadDecode_2_io_rrd_uop_ctrl_op2_sel; // @[register-read.scala 92:29]
    REG_5_ctrl_imm_sel <= RegisterReadDecode_2_io_rrd_uop_ctrl_imm_sel; // @[register-read.scala 92:29]
    REG_5_ctrl_op_fcn <= RegisterReadDecode_2_io_rrd_uop_ctrl_op_fcn; // @[register-read.scala 92:29]
    REG_5_ctrl_fcn_dw <= RegisterReadDecode_2_io_rrd_uop_ctrl_fcn_dw; // @[register-read.scala 92:29]
    REG_5_ctrl_csr_cmd <= RegisterReadDecode_2_io_rrd_uop_ctrl_csr_cmd; // @[register-read.scala 92:29]
    REG_5_ctrl_is_load <= RegisterReadDecode_2_io_rrd_uop_ctrl_is_load; // @[register-read.scala 92:29]
    REG_5_ctrl_is_sta <= RegisterReadDecode_2_io_rrd_uop_ctrl_is_sta; // @[register-read.scala 92:29]
    REG_5_ctrl_is_std <= RegisterReadDecode_2_io_rrd_uop_ctrl_is_std; // @[register-read.scala 92:29]
    REG_5_ctrl_op3_sel <= RegisterReadDecode_2_io_rrd_uop_ctrl_op3_sel; // @[register-read.scala 92:29]
    REG_5_iw_state <= RegisterReadDecode_2_io_rrd_uop_iw_state; // @[register-read.scala 92:29]
    REG_5_iw_p1_poisoned <= RegisterReadDecode_2_io_rrd_uop_iw_p1_poisoned; // @[register-read.scala 92:29]
    REG_5_iw_p2_poisoned <= RegisterReadDecode_2_io_rrd_uop_iw_p2_poisoned; // @[register-read.scala 92:29]
    REG_5_is_br <= RegisterReadDecode_2_io_rrd_uop_is_br; // @[register-read.scala 92:29]
    REG_5_is_jalr <= RegisterReadDecode_2_io_rrd_uop_is_jalr; // @[register-read.scala 92:29]
    REG_5_is_jal <= RegisterReadDecode_2_io_rrd_uop_is_jal; // @[register-read.scala 92:29]
    REG_5_is_sfb <= RegisterReadDecode_2_io_rrd_uop_is_sfb; // @[register-read.scala 92:29]
    REG_5_br_mask <= RegisterReadDecode_2_io_rrd_uop_br_mask & _T_4; // @[util.scala 131:35]
    REG_5_br_tag <= RegisterReadDecode_2_io_rrd_uop_br_tag; // @[register-read.scala 92:29]
    REG_5_ftq_idx <= RegisterReadDecode_2_io_rrd_uop_ftq_idx; // @[register-read.scala 92:29]
    REG_5_edge_inst <= RegisterReadDecode_2_io_rrd_uop_edge_inst; // @[register-read.scala 92:29]
    REG_5_pc_lob <= RegisterReadDecode_2_io_rrd_uop_pc_lob; // @[register-read.scala 92:29]
    REG_5_taken <= RegisterReadDecode_2_io_rrd_uop_taken; // @[register-read.scala 92:29]
    REG_5_imm_packed <= RegisterReadDecode_2_io_rrd_uop_imm_packed; // @[register-read.scala 92:29]
    REG_5_csr_addr <= RegisterReadDecode_2_io_rrd_uop_csr_addr; // @[register-read.scala 92:29]
    REG_5_rob_idx <= RegisterReadDecode_2_io_rrd_uop_rob_idx; // @[register-read.scala 92:29]
    REG_5_ldq_idx <= RegisterReadDecode_2_io_rrd_uop_ldq_idx; // @[register-read.scala 92:29]
    REG_5_stq_idx <= RegisterReadDecode_2_io_rrd_uop_stq_idx; // @[register-read.scala 92:29]
    REG_5_rxq_idx <= RegisterReadDecode_2_io_rrd_uop_rxq_idx; // @[register-read.scala 92:29]
    REG_5_pdst <= RegisterReadDecode_2_io_rrd_uop_pdst; // @[register-read.scala 92:29]
    REG_5_prs1 <= RegisterReadDecode_2_io_rrd_uop_prs1; // @[register-read.scala 92:29]
    REG_5_prs2 <= RegisterReadDecode_2_io_rrd_uop_prs2; // @[register-read.scala 92:29]
    REG_5_prs3 <= RegisterReadDecode_2_io_rrd_uop_prs3; // @[register-read.scala 92:29]
    REG_5_ppred <= RegisterReadDecode_2_io_rrd_uop_ppred; // @[register-read.scala 92:29]
    REG_5_prs1_busy <= RegisterReadDecode_2_io_rrd_uop_prs1_busy; // @[register-read.scala 92:29]
    REG_5_prs2_busy <= RegisterReadDecode_2_io_rrd_uop_prs2_busy; // @[register-read.scala 92:29]
    REG_5_prs3_busy <= RegisterReadDecode_2_io_rrd_uop_prs3_busy; // @[register-read.scala 92:29]
    REG_5_ppred_busy <= RegisterReadDecode_2_io_rrd_uop_ppred_busy; // @[register-read.scala 92:29]
    REG_5_stale_pdst <= RegisterReadDecode_2_io_rrd_uop_stale_pdst; // @[register-read.scala 92:29]
    REG_5_exception <= RegisterReadDecode_2_io_rrd_uop_exception; // @[register-read.scala 92:29]
    REG_5_exc_cause <= RegisterReadDecode_2_io_rrd_uop_exc_cause; // @[register-read.scala 92:29]
    REG_5_bypassable <= RegisterReadDecode_2_io_rrd_uop_bypassable; // @[register-read.scala 92:29]
    REG_5_mem_cmd <= RegisterReadDecode_2_io_rrd_uop_mem_cmd; // @[register-read.scala 92:29]
    REG_5_mem_size <= RegisterReadDecode_2_io_rrd_uop_mem_size; // @[register-read.scala 92:29]
    REG_5_mem_signed <= RegisterReadDecode_2_io_rrd_uop_mem_signed; // @[register-read.scala 92:29]
    REG_5_is_fence <= RegisterReadDecode_2_io_rrd_uop_is_fence; // @[register-read.scala 92:29]
    REG_5_is_fencei <= RegisterReadDecode_2_io_rrd_uop_is_fencei; // @[register-read.scala 92:29]
    REG_5_is_amo <= RegisterReadDecode_2_io_rrd_uop_is_amo; // @[register-read.scala 92:29]
    REG_5_uses_ldq <= RegisterReadDecode_2_io_rrd_uop_uses_ldq; // @[register-read.scala 92:29]
    REG_5_uses_stq <= RegisterReadDecode_2_io_rrd_uop_uses_stq; // @[register-read.scala 92:29]
    REG_5_is_sys_pc2epc <= RegisterReadDecode_2_io_rrd_uop_is_sys_pc2epc; // @[register-read.scala 92:29]
    REG_5_is_unique <= RegisterReadDecode_2_io_rrd_uop_is_unique; // @[register-read.scala 92:29]
    REG_5_flush_on_commit <= RegisterReadDecode_2_io_rrd_uop_flush_on_commit; // @[register-read.scala 92:29]
    REG_5_ldst_is_rs1 <= RegisterReadDecode_2_io_rrd_uop_ldst_is_rs1; // @[register-read.scala 92:29]
    REG_5_ldst <= RegisterReadDecode_2_io_rrd_uop_ldst; // @[register-read.scala 92:29]
    REG_5_lrs1 <= RegisterReadDecode_2_io_rrd_uop_lrs1; // @[register-read.scala 92:29]
    REG_5_lrs2 <= RegisterReadDecode_2_io_rrd_uop_lrs2; // @[register-read.scala 92:29]
    REG_5_lrs3 <= RegisterReadDecode_2_io_rrd_uop_lrs3; // @[register-read.scala 92:29]
    REG_5_ldst_val <= RegisterReadDecode_2_io_rrd_uop_ldst_val; // @[register-read.scala 92:29]
    REG_5_dst_rtype <= RegisterReadDecode_2_io_rrd_uop_dst_rtype; // @[register-read.scala 92:29]
    REG_5_lrs1_rtype <= RegisterReadDecode_2_io_rrd_uop_lrs1_rtype; // @[register-read.scala 92:29]
    REG_5_lrs2_rtype <= RegisterReadDecode_2_io_rrd_uop_lrs2_rtype; // @[register-read.scala 92:29]
    REG_5_frs3_en <= RegisterReadDecode_2_io_rrd_uop_frs3_en; // @[register-read.scala 92:29]
    REG_5_fp_val <= RegisterReadDecode_2_io_rrd_uop_fp_val; // @[register-read.scala 92:29]
    REG_5_fp_single <= RegisterReadDecode_2_io_rrd_uop_fp_single; // @[register-read.scala 92:29]
    REG_5_xcpt_pf_if <= RegisterReadDecode_2_io_rrd_uop_xcpt_pf_if; // @[register-read.scala 92:29]
    REG_5_xcpt_ae_if <= RegisterReadDecode_2_io_rrd_uop_xcpt_ae_if; // @[register-read.scala 92:29]
    REG_5_xcpt_ma_if <= RegisterReadDecode_2_io_rrd_uop_xcpt_ma_if; // @[register-read.scala 92:29]
    REG_5_bp_debug_if <= RegisterReadDecode_2_io_rrd_uop_bp_debug_if; // @[register-read.scala 92:29]
    REG_5_bp_xcpt_if <= RegisterReadDecode_2_io_rrd_uop_bp_xcpt_if; // @[register-read.scala 92:29]
    REG_5_debug_fsrc <= RegisterReadDecode_2_io_rrd_uop_debug_fsrc; // @[register-read.scala 92:29]
    REG_5_debug_tsrc <= RegisterReadDecode_2_io_rrd_uop_debug_tsrc; // @[register-read.scala 92:29]
    REG_6 <= io_iss_uops_0_prs1 == 7'h0 & ~io_iss_uops_0_is_unicore; // @[register-read.scala 134:75]
    REG_7 <= io_iss_uops_0_prs2 == 7'h0 & _T_19; // @[register-read.scala 135:75]
    REG_8 <= io_iss_uops_0_prs3 == 7'h0 & _T_19; // @[register-read.scala 136:75]
    REG_9 <= io_iss_uops_0_rflag & io_iss_uops_0_is_unicore; // @[register-read.scala 143:58]
    REG_10 <= io_iss_uops_1_prs1 == 7'h0 & ~io_iss_uops_1_is_unicore; // @[register-read.scala 134:75]
    REG_11 <= io_iss_uops_1_prs2 == 7'h0 & _T_40; // @[register-read.scala 135:75]
    REG_12 <= io_iss_uops_1_prs3 == 7'h0 & _T_40; // @[register-read.scala 136:75]
    REG_13 <= io_iss_uops_1_rflag & io_iss_uops_1_is_unicore; // @[register-read.scala 143:58]
    REG_14 <= io_iss_uops_2_prs1 == 7'h0 & ~io_iss_uops_2_is_unicore; // @[register-read.scala 134:75]
    REG_15 <= io_iss_uops_2_prs2 == 7'h0 & _T_61; // @[register-read.scala 135:75]
    REG_16 <= io_iss_uops_2_prs3 == 7'h0 & _T_61; // @[register-read.scala 136:75]
    REG_17 <= io_iss_uops_2_rflag & io_iss_uops_2_is_unicore; // @[register-read.scala 143:58]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  exe_reg_valids_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  exe_reg_valids_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  exe_reg_valids_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  exe_reg_uops_0_switch = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  exe_reg_uops_0_switch_off = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  exe_reg_uops_0_is_unicore = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  exe_reg_uops_0_shift = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  exe_reg_uops_0_lrs3_rtype = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  exe_reg_uops_0_rflag = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  exe_reg_uops_0_wflag = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  exe_reg_uops_0_prflag = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  exe_reg_uops_0_pwflag = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  exe_reg_uops_0_pflag_busy = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  exe_reg_uops_0_stale_pflag = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  exe_reg_uops_0_op1_sel = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  exe_reg_uops_0_op2_sel = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  exe_reg_uops_0_split_num = _RAND_16[5:0];
  _RAND_17 = {1{`RANDOM}};
  exe_reg_uops_0_self_index = _RAND_17[5:0];
  _RAND_18 = {1{`RANDOM}};
  exe_reg_uops_0_rob_inst_idx = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
  exe_reg_uops_0_address_num = _RAND_19[5:0];
  _RAND_20 = {1{`RANDOM}};
  exe_reg_uops_0_uopc = _RAND_20[6:0];
  _RAND_21 = {1{`RANDOM}};
  exe_reg_uops_0_inst = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  exe_reg_uops_0_debug_inst = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  exe_reg_uops_0_is_rvc = _RAND_23[0:0];
  _RAND_24 = {2{`RANDOM}};
  exe_reg_uops_0_debug_pc = _RAND_24[39:0];
  _RAND_25 = {1{`RANDOM}};
  exe_reg_uops_0_iq_type = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  exe_reg_uops_0_fu_code = _RAND_26[9:0];
  _RAND_27 = {1{`RANDOM}};
  exe_reg_uops_0_ctrl_br_type = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  exe_reg_uops_0_ctrl_op1_sel = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  exe_reg_uops_0_ctrl_op2_sel = _RAND_29[2:0];
  _RAND_30 = {1{`RANDOM}};
  exe_reg_uops_0_ctrl_imm_sel = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  exe_reg_uops_0_ctrl_op_fcn = _RAND_31[3:0];
  _RAND_32 = {1{`RANDOM}};
  exe_reg_uops_0_ctrl_fcn_dw = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  exe_reg_uops_0_ctrl_csr_cmd = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  exe_reg_uops_0_ctrl_is_load = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  exe_reg_uops_0_ctrl_is_sta = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  exe_reg_uops_0_ctrl_is_std = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  exe_reg_uops_0_ctrl_op3_sel = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  exe_reg_uops_0_iw_state = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  exe_reg_uops_0_iw_p1_poisoned = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  exe_reg_uops_0_iw_p2_poisoned = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  exe_reg_uops_0_is_br = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  exe_reg_uops_0_is_jalr = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  exe_reg_uops_0_is_jal = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  exe_reg_uops_0_is_sfb = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  exe_reg_uops_0_br_mask = _RAND_45[11:0];
  _RAND_46 = {1{`RANDOM}};
  exe_reg_uops_0_br_tag = _RAND_46[3:0];
  _RAND_47 = {1{`RANDOM}};
  exe_reg_uops_0_ftq_idx = _RAND_47[4:0];
  _RAND_48 = {1{`RANDOM}};
  exe_reg_uops_0_edge_inst = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  exe_reg_uops_0_pc_lob = _RAND_49[5:0];
  _RAND_50 = {1{`RANDOM}};
  exe_reg_uops_0_taken = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  exe_reg_uops_0_imm_packed = _RAND_51[19:0];
  _RAND_52 = {1{`RANDOM}};
  exe_reg_uops_0_csr_addr = _RAND_52[11:0];
  _RAND_53 = {1{`RANDOM}};
  exe_reg_uops_0_rob_idx = _RAND_53[5:0];
  _RAND_54 = {1{`RANDOM}};
  exe_reg_uops_0_ldq_idx = _RAND_54[4:0];
  _RAND_55 = {1{`RANDOM}};
  exe_reg_uops_0_stq_idx = _RAND_55[4:0];
  _RAND_56 = {1{`RANDOM}};
  exe_reg_uops_0_rxq_idx = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  exe_reg_uops_0_pdst = _RAND_57[6:0];
  _RAND_58 = {1{`RANDOM}};
  exe_reg_uops_0_prs1 = _RAND_58[6:0];
  _RAND_59 = {1{`RANDOM}};
  exe_reg_uops_0_prs2 = _RAND_59[6:0];
  _RAND_60 = {1{`RANDOM}};
  exe_reg_uops_0_prs3 = _RAND_60[6:0];
  _RAND_61 = {1{`RANDOM}};
  exe_reg_uops_0_ppred = _RAND_61[4:0];
  _RAND_62 = {1{`RANDOM}};
  exe_reg_uops_0_prs1_busy = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  exe_reg_uops_0_prs2_busy = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  exe_reg_uops_0_prs3_busy = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  exe_reg_uops_0_ppred_busy = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  exe_reg_uops_0_stale_pdst = _RAND_66[6:0];
  _RAND_67 = {1{`RANDOM}};
  exe_reg_uops_0_exception = _RAND_67[0:0];
  _RAND_68 = {2{`RANDOM}};
  exe_reg_uops_0_exc_cause = _RAND_68[63:0];
  _RAND_69 = {1{`RANDOM}};
  exe_reg_uops_0_bypassable = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  exe_reg_uops_0_mem_cmd = _RAND_70[4:0];
  _RAND_71 = {1{`RANDOM}};
  exe_reg_uops_0_mem_size = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  exe_reg_uops_0_mem_signed = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  exe_reg_uops_0_is_fence = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  exe_reg_uops_0_is_fencei = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  exe_reg_uops_0_is_amo = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  exe_reg_uops_0_uses_ldq = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  exe_reg_uops_0_uses_stq = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  exe_reg_uops_0_is_sys_pc2epc = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  exe_reg_uops_0_is_unique = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  exe_reg_uops_0_flush_on_commit = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  exe_reg_uops_0_ldst_is_rs1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  exe_reg_uops_0_ldst = _RAND_82[5:0];
  _RAND_83 = {1{`RANDOM}};
  exe_reg_uops_0_lrs1 = _RAND_83[5:0];
  _RAND_84 = {1{`RANDOM}};
  exe_reg_uops_0_lrs2 = _RAND_84[5:0];
  _RAND_85 = {1{`RANDOM}};
  exe_reg_uops_0_lrs3 = _RAND_85[5:0];
  _RAND_86 = {1{`RANDOM}};
  exe_reg_uops_0_ldst_val = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  exe_reg_uops_0_dst_rtype = _RAND_87[1:0];
  _RAND_88 = {1{`RANDOM}};
  exe_reg_uops_0_lrs1_rtype = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  exe_reg_uops_0_lrs2_rtype = _RAND_89[1:0];
  _RAND_90 = {1{`RANDOM}};
  exe_reg_uops_0_frs3_en = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  exe_reg_uops_0_fp_val = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  exe_reg_uops_0_fp_single = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  exe_reg_uops_0_xcpt_pf_if = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  exe_reg_uops_0_xcpt_ae_if = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  exe_reg_uops_0_xcpt_ma_if = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  exe_reg_uops_0_bp_debug_if = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  exe_reg_uops_0_bp_xcpt_if = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  exe_reg_uops_0_debug_fsrc = _RAND_98[1:0];
  _RAND_99 = {1{`RANDOM}};
  exe_reg_uops_0_debug_tsrc = _RAND_99[1:0];
  _RAND_100 = {1{`RANDOM}};
  exe_reg_uops_1_switch = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  exe_reg_uops_1_switch_off = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  exe_reg_uops_1_is_unicore = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  exe_reg_uops_1_shift = _RAND_103[2:0];
  _RAND_104 = {1{`RANDOM}};
  exe_reg_uops_1_lrs3_rtype = _RAND_104[1:0];
  _RAND_105 = {1{`RANDOM}};
  exe_reg_uops_1_rflag = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  exe_reg_uops_1_wflag = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  exe_reg_uops_1_prflag = _RAND_107[3:0];
  _RAND_108 = {1{`RANDOM}};
  exe_reg_uops_1_pwflag = _RAND_108[3:0];
  _RAND_109 = {1{`RANDOM}};
  exe_reg_uops_1_pflag_busy = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  exe_reg_uops_1_stale_pflag = _RAND_110[3:0];
  _RAND_111 = {1{`RANDOM}};
  exe_reg_uops_1_op1_sel = _RAND_111[3:0];
  _RAND_112 = {1{`RANDOM}};
  exe_reg_uops_1_op2_sel = _RAND_112[3:0];
  _RAND_113 = {1{`RANDOM}};
  exe_reg_uops_1_split_num = _RAND_113[5:0];
  _RAND_114 = {1{`RANDOM}};
  exe_reg_uops_1_self_index = _RAND_114[5:0];
  _RAND_115 = {1{`RANDOM}};
  exe_reg_uops_1_rob_inst_idx = _RAND_115[5:0];
  _RAND_116 = {1{`RANDOM}};
  exe_reg_uops_1_address_num = _RAND_116[5:0];
  _RAND_117 = {1{`RANDOM}};
  exe_reg_uops_1_uopc = _RAND_117[6:0];
  _RAND_118 = {1{`RANDOM}};
  exe_reg_uops_1_inst = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  exe_reg_uops_1_debug_inst = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  exe_reg_uops_1_is_rvc = _RAND_120[0:0];
  _RAND_121 = {2{`RANDOM}};
  exe_reg_uops_1_debug_pc = _RAND_121[39:0];
  _RAND_122 = {1{`RANDOM}};
  exe_reg_uops_1_iq_type = _RAND_122[2:0];
  _RAND_123 = {1{`RANDOM}};
  exe_reg_uops_1_fu_code = _RAND_123[9:0];
  _RAND_124 = {1{`RANDOM}};
  exe_reg_uops_1_ctrl_br_type = _RAND_124[3:0];
  _RAND_125 = {1{`RANDOM}};
  exe_reg_uops_1_ctrl_op1_sel = _RAND_125[1:0];
  _RAND_126 = {1{`RANDOM}};
  exe_reg_uops_1_ctrl_op2_sel = _RAND_126[2:0];
  _RAND_127 = {1{`RANDOM}};
  exe_reg_uops_1_ctrl_imm_sel = _RAND_127[2:0];
  _RAND_128 = {1{`RANDOM}};
  exe_reg_uops_1_ctrl_op_fcn = _RAND_128[3:0];
  _RAND_129 = {1{`RANDOM}};
  exe_reg_uops_1_ctrl_fcn_dw = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  exe_reg_uops_1_ctrl_csr_cmd = _RAND_130[2:0];
  _RAND_131 = {1{`RANDOM}};
  exe_reg_uops_1_ctrl_is_load = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  exe_reg_uops_1_ctrl_is_sta = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  exe_reg_uops_1_ctrl_is_std = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  exe_reg_uops_1_ctrl_op3_sel = _RAND_134[1:0];
  _RAND_135 = {1{`RANDOM}};
  exe_reg_uops_1_iw_state = _RAND_135[1:0];
  _RAND_136 = {1{`RANDOM}};
  exe_reg_uops_1_iw_p1_poisoned = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  exe_reg_uops_1_iw_p2_poisoned = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  exe_reg_uops_1_is_br = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  exe_reg_uops_1_is_jalr = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  exe_reg_uops_1_is_jal = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  exe_reg_uops_1_is_sfb = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  exe_reg_uops_1_br_mask = _RAND_142[11:0];
  _RAND_143 = {1{`RANDOM}};
  exe_reg_uops_1_br_tag = _RAND_143[3:0];
  _RAND_144 = {1{`RANDOM}};
  exe_reg_uops_1_ftq_idx = _RAND_144[4:0];
  _RAND_145 = {1{`RANDOM}};
  exe_reg_uops_1_edge_inst = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  exe_reg_uops_1_pc_lob = _RAND_146[5:0];
  _RAND_147 = {1{`RANDOM}};
  exe_reg_uops_1_taken = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  exe_reg_uops_1_imm_packed = _RAND_148[19:0];
  _RAND_149 = {1{`RANDOM}};
  exe_reg_uops_1_csr_addr = _RAND_149[11:0];
  _RAND_150 = {1{`RANDOM}};
  exe_reg_uops_1_rob_idx = _RAND_150[5:0];
  _RAND_151 = {1{`RANDOM}};
  exe_reg_uops_1_ldq_idx = _RAND_151[4:0];
  _RAND_152 = {1{`RANDOM}};
  exe_reg_uops_1_stq_idx = _RAND_152[4:0];
  _RAND_153 = {1{`RANDOM}};
  exe_reg_uops_1_rxq_idx = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  exe_reg_uops_1_pdst = _RAND_154[6:0];
  _RAND_155 = {1{`RANDOM}};
  exe_reg_uops_1_prs1 = _RAND_155[6:0];
  _RAND_156 = {1{`RANDOM}};
  exe_reg_uops_1_prs2 = _RAND_156[6:0];
  _RAND_157 = {1{`RANDOM}};
  exe_reg_uops_1_prs3 = _RAND_157[6:0];
  _RAND_158 = {1{`RANDOM}};
  exe_reg_uops_1_ppred = _RAND_158[4:0];
  _RAND_159 = {1{`RANDOM}};
  exe_reg_uops_1_prs1_busy = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  exe_reg_uops_1_prs2_busy = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  exe_reg_uops_1_prs3_busy = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  exe_reg_uops_1_ppred_busy = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  exe_reg_uops_1_stale_pdst = _RAND_163[6:0];
  _RAND_164 = {1{`RANDOM}};
  exe_reg_uops_1_exception = _RAND_164[0:0];
  _RAND_165 = {2{`RANDOM}};
  exe_reg_uops_1_exc_cause = _RAND_165[63:0];
  _RAND_166 = {1{`RANDOM}};
  exe_reg_uops_1_bypassable = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  exe_reg_uops_1_mem_cmd = _RAND_167[4:0];
  _RAND_168 = {1{`RANDOM}};
  exe_reg_uops_1_mem_size = _RAND_168[1:0];
  _RAND_169 = {1{`RANDOM}};
  exe_reg_uops_1_mem_signed = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  exe_reg_uops_1_is_fence = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  exe_reg_uops_1_is_fencei = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  exe_reg_uops_1_is_amo = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  exe_reg_uops_1_uses_ldq = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  exe_reg_uops_1_uses_stq = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  exe_reg_uops_1_is_sys_pc2epc = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  exe_reg_uops_1_is_unique = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  exe_reg_uops_1_flush_on_commit = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  exe_reg_uops_1_ldst_is_rs1 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  exe_reg_uops_1_ldst = _RAND_179[5:0];
  _RAND_180 = {1{`RANDOM}};
  exe_reg_uops_1_lrs1 = _RAND_180[5:0];
  _RAND_181 = {1{`RANDOM}};
  exe_reg_uops_1_lrs2 = _RAND_181[5:0];
  _RAND_182 = {1{`RANDOM}};
  exe_reg_uops_1_lrs3 = _RAND_182[5:0];
  _RAND_183 = {1{`RANDOM}};
  exe_reg_uops_1_ldst_val = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  exe_reg_uops_1_dst_rtype = _RAND_184[1:0];
  _RAND_185 = {1{`RANDOM}};
  exe_reg_uops_1_lrs1_rtype = _RAND_185[1:0];
  _RAND_186 = {1{`RANDOM}};
  exe_reg_uops_1_lrs2_rtype = _RAND_186[1:0];
  _RAND_187 = {1{`RANDOM}};
  exe_reg_uops_1_frs3_en = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  exe_reg_uops_1_fp_val = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  exe_reg_uops_1_fp_single = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  exe_reg_uops_1_xcpt_pf_if = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  exe_reg_uops_1_xcpt_ae_if = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  exe_reg_uops_1_xcpt_ma_if = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  exe_reg_uops_1_bp_debug_if = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  exe_reg_uops_1_bp_xcpt_if = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  exe_reg_uops_1_debug_fsrc = _RAND_195[1:0];
  _RAND_196 = {1{`RANDOM}};
  exe_reg_uops_1_debug_tsrc = _RAND_196[1:0];
  _RAND_197 = {1{`RANDOM}};
  exe_reg_uops_2_switch = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  exe_reg_uops_2_switch_off = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  exe_reg_uops_2_is_unicore = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  exe_reg_uops_2_shift = _RAND_200[2:0];
  _RAND_201 = {1{`RANDOM}};
  exe_reg_uops_2_lrs3_rtype = _RAND_201[1:0];
  _RAND_202 = {1{`RANDOM}};
  exe_reg_uops_2_rflag = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  exe_reg_uops_2_wflag = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  exe_reg_uops_2_prflag = _RAND_204[3:0];
  _RAND_205 = {1{`RANDOM}};
  exe_reg_uops_2_pwflag = _RAND_205[3:0];
  _RAND_206 = {1{`RANDOM}};
  exe_reg_uops_2_pflag_busy = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  exe_reg_uops_2_stale_pflag = _RAND_207[3:0];
  _RAND_208 = {1{`RANDOM}};
  exe_reg_uops_2_op1_sel = _RAND_208[3:0];
  _RAND_209 = {1{`RANDOM}};
  exe_reg_uops_2_op2_sel = _RAND_209[3:0];
  _RAND_210 = {1{`RANDOM}};
  exe_reg_uops_2_split_num = _RAND_210[5:0];
  _RAND_211 = {1{`RANDOM}};
  exe_reg_uops_2_self_index = _RAND_211[5:0];
  _RAND_212 = {1{`RANDOM}};
  exe_reg_uops_2_rob_inst_idx = _RAND_212[5:0];
  _RAND_213 = {1{`RANDOM}};
  exe_reg_uops_2_address_num = _RAND_213[5:0];
  _RAND_214 = {1{`RANDOM}};
  exe_reg_uops_2_uopc = _RAND_214[6:0];
  _RAND_215 = {1{`RANDOM}};
  exe_reg_uops_2_inst = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  exe_reg_uops_2_debug_inst = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  exe_reg_uops_2_is_rvc = _RAND_217[0:0];
  _RAND_218 = {2{`RANDOM}};
  exe_reg_uops_2_debug_pc = _RAND_218[39:0];
  _RAND_219 = {1{`RANDOM}};
  exe_reg_uops_2_iq_type = _RAND_219[2:0];
  _RAND_220 = {1{`RANDOM}};
  exe_reg_uops_2_fu_code = _RAND_220[9:0];
  _RAND_221 = {1{`RANDOM}};
  exe_reg_uops_2_ctrl_br_type = _RAND_221[3:0];
  _RAND_222 = {1{`RANDOM}};
  exe_reg_uops_2_ctrl_op1_sel = _RAND_222[1:0];
  _RAND_223 = {1{`RANDOM}};
  exe_reg_uops_2_ctrl_op2_sel = _RAND_223[2:0];
  _RAND_224 = {1{`RANDOM}};
  exe_reg_uops_2_ctrl_imm_sel = _RAND_224[2:0];
  _RAND_225 = {1{`RANDOM}};
  exe_reg_uops_2_ctrl_op_fcn = _RAND_225[3:0];
  _RAND_226 = {1{`RANDOM}};
  exe_reg_uops_2_ctrl_fcn_dw = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  exe_reg_uops_2_ctrl_csr_cmd = _RAND_227[2:0];
  _RAND_228 = {1{`RANDOM}};
  exe_reg_uops_2_ctrl_is_load = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  exe_reg_uops_2_ctrl_is_sta = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  exe_reg_uops_2_ctrl_is_std = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  exe_reg_uops_2_ctrl_op3_sel = _RAND_231[1:0];
  _RAND_232 = {1{`RANDOM}};
  exe_reg_uops_2_iw_state = _RAND_232[1:0];
  _RAND_233 = {1{`RANDOM}};
  exe_reg_uops_2_iw_p1_poisoned = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  exe_reg_uops_2_iw_p2_poisoned = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  exe_reg_uops_2_is_br = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  exe_reg_uops_2_is_jalr = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  exe_reg_uops_2_is_jal = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  exe_reg_uops_2_is_sfb = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  exe_reg_uops_2_br_mask = _RAND_239[11:0];
  _RAND_240 = {1{`RANDOM}};
  exe_reg_uops_2_br_tag = _RAND_240[3:0];
  _RAND_241 = {1{`RANDOM}};
  exe_reg_uops_2_ftq_idx = _RAND_241[4:0];
  _RAND_242 = {1{`RANDOM}};
  exe_reg_uops_2_edge_inst = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  exe_reg_uops_2_pc_lob = _RAND_243[5:0];
  _RAND_244 = {1{`RANDOM}};
  exe_reg_uops_2_taken = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  exe_reg_uops_2_imm_packed = _RAND_245[19:0];
  _RAND_246 = {1{`RANDOM}};
  exe_reg_uops_2_csr_addr = _RAND_246[11:0];
  _RAND_247 = {1{`RANDOM}};
  exe_reg_uops_2_rob_idx = _RAND_247[5:0];
  _RAND_248 = {1{`RANDOM}};
  exe_reg_uops_2_ldq_idx = _RAND_248[4:0];
  _RAND_249 = {1{`RANDOM}};
  exe_reg_uops_2_stq_idx = _RAND_249[4:0];
  _RAND_250 = {1{`RANDOM}};
  exe_reg_uops_2_rxq_idx = _RAND_250[1:0];
  _RAND_251 = {1{`RANDOM}};
  exe_reg_uops_2_pdst = _RAND_251[6:0];
  _RAND_252 = {1{`RANDOM}};
  exe_reg_uops_2_prs1 = _RAND_252[6:0];
  _RAND_253 = {1{`RANDOM}};
  exe_reg_uops_2_prs2 = _RAND_253[6:0];
  _RAND_254 = {1{`RANDOM}};
  exe_reg_uops_2_prs3 = _RAND_254[6:0];
  _RAND_255 = {1{`RANDOM}};
  exe_reg_uops_2_ppred = _RAND_255[4:0];
  _RAND_256 = {1{`RANDOM}};
  exe_reg_uops_2_prs1_busy = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  exe_reg_uops_2_prs2_busy = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  exe_reg_uops_2_prs3_busy = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  exe_reg_uops_2_ppred_busy = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  exe_reg_uops_2_stale_pdst = _RAND_260[6:0];
  _RAND_261 = {1{`RANDOM}};
  exe_reg_uops_2_exception = _RAND_261[0:0];
  _RAND_262 = {2{`RANDOM}};
  exe_reg_uops_2_exc_cause = _RAND_262[63:0];
  _RAND_263 = {1{`RANDOM}};
  exe_reg_uops_2_bypassable = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  exe_reg_uops_2_mem_cmd = _RAND_264[4:0];
  _RAND_265 = {1{`RANDOM}};
  exe_reg_uops_2_mem_size = _RAND_265[1:0];
  _RAND_266 = {1{`RANDOM}};
  exe_reg_uops_2_mem_signed = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  exe_reg_uops_2_is_fence = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  exe_reg_uops_2_is_fencei = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  exe_reg_uops_2_is_amo = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  exe_reg_uops_2_uses_ldq = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  exe_reg_uops_2_uses_stq = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  exe_reg_uops_2_is_sys_pc2epc = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  exe_reg_uops_2_is_unique = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  exe_reg_uops_2_flush_on_commit = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  exe_reg_uops_2_ldst_is_rs1 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  exe_reg_uops_2_ldst = _RAND_276[5:0];
  _RAND_277 = {1{`RANDOM}};
  exe_reg_uops_2_lrs1 = _RAND_277[5:0];
  _RAND_278 = {1{`RANDOM}};
  exe_reg_uops_2_lrs2 = _RAND_278[5:0];
  _RAND_279 = {1{`RANDOM}};
  exe_reg_uops_2_lrs3 = _RAND_279[5:0];
  _RAND_280 = {1{`RANDOM}};
  exe_reg_uops_2_ldst_val = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  exe_reg_uops_2_dst_rtype = _RAND_281[1:0];
  _RAND_282 = {1{`RANDOM}};
  exe_reg_uops_2_lrs1_rtype = _RAND_282[1:0];
  _RAND_283 = {1{`RANDOM}};
  exe_reg_uops_2_lrs2_rtype = _RAND_283[1:0];
  _RAND_284 = {1{`RANDOM}};
  exe_reg_uops_2_frs3_en = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  exe_reg_uops_2_fp_val = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  exe_reg_uops_2_fp_single = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  exe_reg_uops_2_xcpt_pf_if = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  exe_reg_uops_2_xcpt_ae_if = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  exe_reg_uops_2_xcpt_ma_if = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  exe_reg_uops_2_bp_debug_if = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  exe_reg_uops_2_bp_xcpt_if = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  exe_reg_uops_2_debug_fsrc = _RAND_292[1:0];
  _RAND_293 = {1{`RANDOM}};
  exe_reg_uops_2_debug_tsrc = _RAND_293[1:0];
  _RAND_294 = {2{`RANDOM}};
  exe_reg_rs1_data_0 = _RAND_294[63:0];
  _RAND_295 = {2{`RANDOM}};
  exe_reg_rs1_data_1 = _RAND_295[63:0];
  _RAND_296 = {2{`RANDOM}};
  exe_reg_rs1_data_2 = _RAND_296[63:0];
  _RAND_297 = {2{`RANDOM}};
  exe_reg_rs2_data_0 = _RAND_297[63:0];
  _RAND_298 = {2{`RANDOM}};
  exe_reg_rs2_data_1 = _RAND_298[63:0];
  _RAND_299 = {2{`RANDOM}};
  exe_reg_rs2_data_2 = _RAND_299[63:0];
  _RAND_300 = {2{`RANDOM}};
  exe_reg_rs3_data_0 = _RAND_300[63:0];
  _RAND_301 = {2{`RANDOM}};
  exe_reg_rs3_data_1 = _RAND_301[63:0];
  _RAND_302 = {2{`RANDOM}};
  exe_reg_rs3_data_2 = _RAND_302[63:0];
  _RAND_303 = {1{`RANDOM}};
  exe_reg_flag_data_0 = _RAND_303[3:0];
  _RAND_304 = {1{`RANDOM}};
  exe_reg_flag_data_1 = _RAND_304[3:0];
  _RAND_305 = {1{`RANDOM}};
  exe_reg_flag_data_2 = _RAND_305[3:0];
  _RAND_306 = {1{`RANDOM}};
  REG = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  REG_1_switch = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  REG_1_switch_off = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  REG_1_is_unicore = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  REG_1_shift = _RAND_310[2:0];
  _RAND_311 = {1{`RANDOM}};
  REG_1_lrs3_rtype = _RAND_311[1:0];
  _RAND_312 = {1{`RANDOM}};
  REG_1_rflag = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  REG_1_wflag = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  REG_1_prflag = _RAND_314[3:0];
  _RAND_315 = {1{`RANDOM}};
  REG_1_pwflag = _RAND_315[3:0];
  _RAND_316 = {1{`RANDOM}};
  REG_1_pflag_busy = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  REG_1_stale_pflag = _RAND_317[3:0];
  _RAND_318 = {1{`RANDOM}};
  REG_1_op1_sel = _RAND_318[3:0];
  _RAND_319 = {1{`RANDOM}};
  REG_1_op2_sel = _RAND_319[3:0];
  _RAND_320 = {1{`RANDOM}};
  REG_1_split_num = _RAND_320[5:0];
  _RAND_321 = {1{`RANDOM}};
  REG_1_self_index = _RAND_321[5:0];
  _RAND_322 = {1{`RANDOM}};
  REG_1_rob_inst_idx = _RAND_322[5:0];
  _RAND_323 = {1{`RANDOM}};
  REG_1_address_num = _RAND_323[5:0];
  _RAND_324 = {1{`RANDOM}};
  REG_1_uopc = _RAND_324[6:0];
  _RAND_325 = {1{`RANDOM}};
  REG_1_inst = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  REG_1_debug_inst = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  REG_1_is_rvc = _RAND_327[0:0];
  _RAND_328 = {2{`RANDOM}};
  REG_1_debug_pc = _RAND_328[39:0];
  _RAND_329 = {1{`RANDOM}};
  REG_1_iq_type = _RAND_329[2:0];
  _RAND_330 = {1{`RANDOM}};
  REG_1_fu_code = _RAND_330[9:0];
  _RAND_331 = {1{`RANDOM}};
  REG_1_ctrl_br_type = _RAND_331[3:0];
  _RAND_332 = {1{`RANDOM}};
  REG_1_ctrl_op1_sel = _RAND_332[1:0];
  _RAND_333 = {1{`RANDOM}};
  REG_1_ctrl_op2_sel = _RAND_333[2:0];
  _RAND_334 = {1{`RANDOM}};
  REG_1_ctrl_imm_sel = _RAND_334[2:0];
  _RAND_335 = {1{`RANDOM}};
  REG_1_ctrl_op_fcn = _RAND_335[3:0];
  _RAND_336 = {1{`RANDOM}};
  REG_1_ctrl_fcn_dw = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  REG_1_ctrl_csr_cmd = _RAND_337[2:0];
  _RAND_338 = {1{`RANDOM}};
  REG_1_ctrl_is_load = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  REG_1_ctrl_is_sta = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  REG_1_ctrl_is_std = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  REG_1_ctrl_op3_sel = _RAND_341[1:0];
  _RAND_342 = {1{`RANDOM}};
  REG_1_iw_state = _RAND_342[1:0];
  _RAND_343 = {1{`RANDOM}};
  REG_1_iw_p1_poisoned = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  REG_1_iw_p2_poisoned = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  REG_1_is_br = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  REG_1_is_jalr = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  REG_1_is_jal = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  REG_1_is_sfb = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  REG_1_br_mask = _RAND_349[11:0];
  _RAND_350 = {1{`RANDOM}};
  REG_1_br_tag = _RAND_350[3:0];
  _RAND_351 = {1{`RANDOM}};
  REG_1_ftq_idx = _RAND_351[4:0];
  _RAND_352 = {1{`RANDOM}};
  REG_1_edge_inst = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  REG_1_pc_lob = _RAND_353[5:0];
  _RAND_354 = {1{`RANDOM}};
  REG_1_taken = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  REG_1_imm_packed = _RAND_355[19:0];
  _RAND_356 = {1{`RANDOM}};
  REG_1_csr_addr = _RAND_356[11:0];
  _RAND_357 = {1{`RANDOM}};
  REG_1_rob_idx = _RAND_357[5:0];
  _RAND_358 = {1{`RANDOM}};
  REG_1_ldq_idx = _RAND_358[4:0];
  _RAND_359 = {1{`RANDOM}};
  REG_1_stq_idx = _RAND_359[4:0];
  _RAND_360 = {1{`RANDOM}};
  REG_1_rxq_idx = _RAND_360[1:0];
  _RAND_361 = {1{`RANDOM}};
  REG_1_pdst = _RAND_361[6:0];
  _RAND_362 = {1{`RANDOM}};
  REG_1_prs1 = _RAND_362[6:0];
  _RAND_363 = {1{`RANDOM}};
  REG_1_prs2 = _RAND_363[6:0];
  _RAND_364 = {1{`RANDOM}};
  REG_1_prs3 = _RAND_364[6:0];
  _RAND_365 = {1{`RANDOM}};
  REG_1_ppred = _RAND_365[4:0];
  _RAND_366 = {1{`RANDOM}};
  REG_1_prs1_busy = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  REG_1_prs2_busy = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  REG_1_prs3_busy = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  REG_1_ppred_busy = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  REG_1_stale_pdst = _RAND_370[6:0];
  _RAND_371 = {1{`RANDOM}};
  REG_1_exception = _RAND_371[0:0];
  _RAND_372 = {2{`RANDOM}};
  REG_1_exc_cause = _RAND_372[63:0];
  _RAND_373 = {1{`RANDOM}};
  REG_1_bypassable = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  REG_1_mem_cmd = _RAND_374[4:0];
  _RAND_375 = {1{`RANDOM}};
  REG_1_mem_size = _RAND_375[1:0];
  _RAND_376 = {1{`RANDOM}};
  REG_1_mem_signed = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  REG_1_is_fence = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  REG_1_is_fencei = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  REG_1_is_amo = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  REG_1_uses_ldq = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  REG_1_uses_stq = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  REG_1_is_sys_pc2epc = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  REG_1_is_unique = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  REG_1_flush_on_commit = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  REG_1_ldst_is_rs1 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  REG_1_ldst = _RAND_386[5:0];
  _RAND_387 = {1{`RANDOM}};
  REG_1_lrs1 = _RAND_387[5:0];
  _RAND_388 = {1{`RANDOM}};
  REG_1_lrs2 = _RAND_388[5:0];
  _RAND_389 = {1{`RANDOM}};
  REG_1_lrs3 = _RAND_389[5:0];
  _RAND_390 = {1{`RANDOM}};
  REG_1_ldst_val = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  REG_1_dst_rtype = _RAND_391[1:0];
  _RAND_392 = {1{`RANDOM}};
  REG_1_lrs1_rtype = _RAND_392[1:0];
  _RAND_393 = {1{`RANDOM}};
  REG_1_lrs2_rtype = _RAND_393[1:0];
  _RAND_394 = {1{`RANDOM}};
  REG_1_frs3_en = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  REG_1_fp_val = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  REG_1_fp_single = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  REG_1_xcpt_pf_if = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  REG_1_xcpt_ae_if = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  REG_1_xcpt_ma_if = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  REG_1_bp_debug_if = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  REG_1_bp_xcpt_if = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  REG_1_debug_fsrc = _RAND_402[1:0];
  _RAND_403 = {1{`RANDOM}};
  REG_1_debug_tsrc = _RAND_403[1:0];
  _RAND_404 = {1{`RANDOM}};
  REG_2 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  REG_3_switch = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  REG_3_switch_off = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  REG_3_is_unicore = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  REG_3_shift = _RAND_408[2:0];
  _RAND_409 = {1{`RANDOM}};
  REG_3_lrs3_rtype = _RAND_409[1:0];
  _RAND_410 = {1{`RANDOM}};
  REG_3_rflag = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  REG_3_wflag = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  REG_3_prflag = _RAND_412[3:0];
  _RAND_413 = {1{`RANDOM}};
  REG_3_pwflag = _RAND_413[3:0];
  _RAND_414 = {1{`RANDOM}};
  REG_3_pflag_busy = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  REG_3_stale_pflag = _RAND_415[3:0];
  _RAND_416 = {1{`RANDOM}};
  REG_3_op1_sel = _RAND_416[3:0];
  _RAND_417 = {1{`RANDOM}};
  REG_3_op2_sel = _RAND_417[3:0];
  _RAND_418 = {1{`RANDOM}};
  REG_3_split_num = _RAND_418[5:0];
  _RAND_419 = {1{`RANDOM}};
  REG_3_self_index = _RAND_419[5:0];
  _RAND_420 = {1{`RANDOM}};
  REG_3_rob_inst_idx = _RAND_420[5:0];
  _RAND_421 = {1{`RANDOM}};
  REG_3_address_num = _RAND_421[5:0];
  _RAND_422 = {1{`RANDOM}};
  REG_3_uopc = _RAND_422[6:0];
  _RAND_423 = {1{`RANDOM}};
  REG_3_inst = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  REG_3_debug_inst = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  REG_3_is_rvc = _RAND_425[0:0];
  _RAND_426 = {2{`RANDOM}};
  REG_3_debug_pc = _RAND_426[39:0];
  _RAND_427 = {1{`RANDOM}};
  REG_3_iq_type = _RAND_427[2:0];
  _RAND_428 = {1{`RANDOM}};
  REG_3_fu_code = _RAND_428[9:0];
  _RAND_429 = {1{`RANDOM}};
  REG_3_ctrl_br_type = _RAND_429[3:0];
  _RAND_430 = {1{`RANDOM}};
  REG_3_ctrl_op1_sel = _RAND_430[1:0];
  _RAND_431 = {1{`RANDOM}};
  REG_3_ctrl_op2_sel = _RAND_431[2:0];
  _RAND_432 = {1{`RANDOM}};
  REG_3_ctrl_imm_sel = _RAND_432[2:0];
  _RAND_433 = {1{`RANDOM}};
  REG_3_ctrl_op_fcn = _RAND_433[3:0];
  _RAND_434 = {1{`RANDOM}};
  REG_3_ctrl_fcn_dw = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  REG_3_ctrl_csr_cmd = _RAND_435[2:0];
  _RAND_436 = {1{`RANDOM}};
  REG_3_ctrl_is_load = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  REG_3_ctrl_is_sta = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  REG_3_ctrl_is_std = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  REG_3_ctrl_op3_sel = _RAND_439[1:0];
  _RAND_440 = {1{`RANDOM}};
  REG_3_iw_state = _RAND_440[1:0];
  _RAND_441 = {1{`RANDOM}};
  REG_3_iw_p1_poisoned = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  REG_3_iw_p2_poisoned = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  REG_3_is_br = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  REG_3_is_jalr = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  REG_3_is_jal = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  REG_3_is_sfb = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  REG_3_br_mask = _RAND_447[11:0];
  _RAND_448 = {1{`RANDOM}};
  REG_3_br_tag = _RAND_448[3:0];
  _RAND_449 = {1{`RANDOM}};
  REG_3_ftq_idx = _RAND_449[4:0];
  _RAND_450 = {1{`RANDOM}};
  REG_3_edge_inst = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  REG_3_pc_lob = _RAND_451[5:0];
  _RAND_452 = {1{`RANDOM}};
  REG_3_taken = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  REG_3_imm_packed = _RAND_453[19:0];
  _RAND_454 = {1{`RANDOM}};
  REG_3_csr_addr = _RAND_454[11:0];
  _RAND_455 = {1{`RANDOM}};
  REG_3_rob_idx = _RAND_455[5:0];
  _RAND_456 = {1{`RANDOM}};
  REG_3_ldq_idx = _RAND_456[4:0];
  _RAND_457 = {1{`RANDOM}};
  REG_3_stq_idx = _RAND_457[4:0];
  _RAND_458 = {1{`RANDOM}};
  REG_3_rxq_idx = _RAND_458[1:0];
  _RAND_459 = {1{`RANDOM}};
  REG_3_pdst = _RAND_459[6:0];
  _RAND_460 = {1{`RANDOM}};
  REG_3_prs1 = _RAND_460[6:0];
  _RAND_461 = {1{`RANDOM}};
  REG_3_prs2 = _RAND_461[6:0];
  _RAND_462 = {1{`RANDOM}};
  REG_3_prs3 = _RAND_462[6:0];
  _RAND_463 = {1{`RANDOM}};
  REG_3_ppred = _RAND_463[4:0];
  _RAND_464 = {1{`RANDOM}};
  REG_3_prs1_busy = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  REG_3_prs2_busy = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  REG_3_prs3_busy = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  REG_3_ppred_busy = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  REG_3_stale_pdst = _RAND_468[6:0];
  _RAND_469 = {1{`RANDOM}};
  REG_3_exception = _RAND_469[0:0];
  _RAND_470 = {2{`RANDOM}};
  REG_3_exc_cause = _RAND_470[63:0];
  _RAND_471 = {1{`RANDOM}};
  REG_3_bypassable = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  REG_3_mem_cmd = _RAND_472[4:0];
  _RAND_473 = {1{`RANDOM}};
  REG_3_mem_size = _RAND_473[1:0];
  _RAND_474 = {1{`RANDOM}};
  REG_3_mem_signed = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  REG_3_is_fence = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  REG_3_is_fencei = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  REG_3_is_amo = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  REG_3_uses_ldq = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  REG_3_uses_stq = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  REG_3_is_sys_pc2epc = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  REG_3_is_unique = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  REG_3_flush_on_commit = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  REG_3_ldst_is_rs1 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  REG_3_ldst = _RAND_484[5:0];
  _RAND_485 = {1{`RANDOM}};
  REG_3_lrs1 = _RAND_485[5:0];
  _RAND_486 = {1{`RANDOM}};
  REG_3_lrs2 = _RAND_486[5:0];
  _RAND_487 = {1{`RANDOM}};
  REG_3_lrs3 = _RAND_487[5:0];
  _RAND_488 = {1{`RANDOM}};
  REG_3_ldst_val = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  REG_3_dst_rtype = _RAND_489[1:0];
  _RAND_490 = {1{`RANDOM}};
  REG_3_lrs1_rtype = _RAND_490[1:0];
  _RAND_491 = {1{`RANDOM}};
  REG_3_lrs2_rtype = _RAND_491[1:0];
  _RAND_492 = {1{`RANDOM}};
  REG_3_frs3_en = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  REG_3_fp_val = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  REG_3_fp_single = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  REG_3_xcpt_pf_if = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  REG_3_xcpt_ae_if = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  REG_3_xcpt_ma_if = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  REG_3_bp_debug_if = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  REG_3_bp_xcpt_if = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  REG_3_debug_fsrc = _RAND_500[1:0];
  _RAND_501 = {1{`RANDOM}};
  REG_3_debug_tsrc = _RAND_501[1:0];
  _RAND_502 = {1{`RANDOM}};
  REG_4 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  REG_5_switch = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  REG_5_switch_off = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  REG_5_is_unicore = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  REG_5_shift = _RAND_506[2:0];
  _RAND_507 = {1{`RANDOM}};
  REG_5_lrs3_rtype = _RAND_507[1:0];
  _RAND_508 = {1{`RANDOM}};
  REG_5_rflag = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  REG_5_wflag = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  REG_5_prflag = _RAND_510[3:0];
  _RAND_511 = {1{`RANDOM}};
  REG_5_pwflag = _RAND_511[3:0];
  _RAND_512 = {1{`RANDOM}};
  REG_5_pflag_busy = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  REG_5_stale_pflag = _RAND_513[3:0];
  _RAND_514 = {1{`RANDOM}};
  REG_5_op1_sel = _RAND_514[3:0];
  _RAND_515 = {1{`RANDOM}};
  REG_5_op2_sel = _RAND_515[3:0];
  _RAND_516 = {1{`RANDOM}};
  REG_5_split_num = _RAND_516[5:0];
  _RAND_517 = {1{`RANDOM}};
  REG_5_self_index = _RAND_517[5:0];
  _RAND_518 = {1{`RANDOM}};
  REG_5_rob_inst_idx = _RAND_518[5:0];
  _RAND_519 = {1{`RANDOM}};
  REG_5_address_num = _RAND_519[5:0];
  _RAND_520 = {1{`RANDOM}};
  REG_5_uopc = _RAND_520[6:0];
  _RAND_521 = {1{`RANDOM}};
  REG_5_inst = _RAND_521[31:0];
  _RAND_522 = {1{`RANDOM}};
  REG_5_debug_inst = _RAND_522[31:0];
  _RAND_523 = {1{`RANDOM}};
  REG_5_is_rvc = _RAND_523[0:0];
  _RAND_524 = {2{`RANDOM}};
  REG_5_debug_pc = _RAND_524[39:0];
  _RAND_525 = {1{`RANDOM}};
  REG_5_iq_type = _RAND_525[2:0];
  _RAND_526 = {1{`RANDOM}};
  REG_5_fu_code = _RAND_526[9:0];
  _RAND_527 = {1{`RANDOM}};
  REG_5_ctrl_br_type = _RAND_527[3:0];
  _RAND_528 = {1{`RANDOM}};
  REG_5_ctrl_op1_sel = _RAND_528[1:0];
  _RAND_529 = {1{`RANDOM}};
  REG_5_ctrl_op2_sel = _RAND_529[2:0];
  _RAND_530 = {1{`RANDOM}};
  REG_5_ctrl_imm_sel = _RAND_530[2:0];
  _RAND_531 = {1{`RANDOM}};
  REG_5_ctrl_op_fcn = _RAND_531[3:0];
  _RAND_532 = {1{`RANDOM}};
  REG_5_ctrl_fcn_dw = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  REG_5_ctrl_csr_cmd = _RAND_533[2:0];
  _RAND_534 = {1{`RANDOM}};
  REG_5_ctrl_is_load = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  REG_5_ctrl_is_sta = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  REG_5_ctrl_is_std = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  REG_5_ctrl_op3_sel = _RAND_537[1:0];
  _RAND_538 = {1{`RANDOM}};
  REG_5_iw_state = _RAND_538[1:0];
  _RAND_539 = {1{`RANDOM}};
  REG_5_iw_p1_poisoned = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  REG_5_iw_p2_poisoned = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  REG_5_is_br = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  REG_5_is_jalr = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  REG_5_is_jal = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  REG_5_is_sfb = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  REG_5_br_mask = _RAND_545[11:0];
  _RAND_546 = {1{`RANDOM}};
  REG_5_br_tag = _RAND_546[3:0];
  _RAND_547 = {1{`RANDOM}};
  REG_5_ftq_idx = _RAND_547[4:0];
  _RAND_548 = {1{`RANDOM}};
  REG_5_edge_inst = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  REG_5_pc_lob = _RAND_549[5:0];
  _RAND_550 = {1{`RANDOM}};
  REG_5_taken = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  REG_5_imm_packed = _RAND_551[19:0];
  _RAND_552 = {1{`RANDOM}};
  REG_5_csr_addr = _RAND_552[11:0];
  _RAND_553 = {1{`RANDOM}};
  REG_5_rob_idx = _RAND_553[5:0];
  _RAND_554 = {1{`RANDOM}};
  REG_5_ldq_idx = _RAND_554[4:0];
  _RAND_555 = {1{`RANDOM}};
  REG_5_stq_idx = _RAND_555[4:0];
  _RAND_556 = {1{`RANDOM}};
  REG_5_rxq_idx = _RAND_556[1:0];
  _RAND_557 = {1{`RANDOM}};
  REG_5_pdst = _RAND_557[6:0];
  _RAND_558 = {1{`RANDOM}};
  REG_5_prs1 = _RAND_558[6:0];
  _RAND_559 = {1{`RANDOM}};
  REG_5_prs2 = _RAND_559[6:0];
  _RAND_560 = {1{`RANDOM}};
  REG_5_prs3 = _RAND_560[6:0];
  _RAND_561 = {1{`RANDOM}};
  REG_5_ppred = _RAND_561[4:0];
  _RAND_562 = {1{`RANDOM}};
  REG_5_prs1_busy = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  REG_5_prs2_busy = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  REG_5_prs3_busy = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  REG_5_ppred_busy = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  REG_5_stale_pdst = _RAND_566[6:0];
  _RAND_567 = {1{`RANDOM}};
  REG_5_exception = _RAND_567[0:0];
  _RAND_568 = {2{`RANDOM}};
  REG_5_exc_cause = _RAND_568[63:0];
  _RAND_569 = {1{`RANDOM}};
  REG_5_bypassable = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  REG_5_mem_cmd = _RAND_570[4:0];
  _RAND_571 = {1{`RANDOM}};
  REG_5_mem_size = _RAND_571[1:0];
  _RAND_572 = {1{`RANDOM}};
  REG_5_mem_signed = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  REG_5_is_fence = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  REG_5_is_fencei = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  REG_5_is_amo = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  REG_5_uses_ldq = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  REG_5_uses_stq = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  REG_5_is_sys_pc2epc = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  REG_5_is_unique = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  REG_5_flush_on_commit = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  REG_5_ldst_is_rs1 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  REG_5_ldst = _RAND_582[5:0];
  _RAND_583 = {1{`RANDOM}};
  REG_5_lrs1 = _RAND_583[5:0];
  _RAND_584 = {1{`RANDOM}};
  REG_5_lrs2 = _RAND_584[5:0];
  _RAND_585 = {1{`RANDOM}};
  REG_5_lrs3 = _RAND_585[5:0];
  _RAND_586 = {1{`RANDOM}};
  REG_5_ldst_val = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  REG_5_dst_rtype = _RAND_587[1:0];
  _RAND_588 = {1{`RANDOM}};
  REG_5_lrs1_rtype = _RAND_588[1:0];
  _RAND_589 = {1{`RANDOM}};
  REG_5_lrs2_rtype = _RAND_589[1:0];
  _RAND_590 = {1{`RANDOM}};
  REG_5_frs3_en = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  REG_5_fp_val = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  REG_5_fp_single = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  REG_5_xcpt_pf_if = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  REG_5_xcpt_ae_if = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  REG_5_xcpt_ma_if = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  REG_5_bp_debug_if = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  REG_5_bp_xcpt_if = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  REG_5_debug_fsrc = _RAND_598[1:0];
  _RAND_599 = {1{`RANDOM}};
  REG_5_debug_tsrc = _RAND_599[1:0];
  _RAND_600 = {1{`RANDOM}};
  REG_6 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  REG_7 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  REG_8 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  REG_9 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  REG_10 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  REG_11 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  REG_12 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  REG_13 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  REG_14 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  REG_15 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  REG_16 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  REG_17 = _RAND_611[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
