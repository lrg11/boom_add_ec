module IssueUnitCollapsing(
  input         clock,
  input         reset,
  output        io_dis_uops_0_ready,
  input         io_dis_uops_0_valid,
  input         io_dis_uops_0_bits_switch,
  input         io_dis_uops_0_bits_switch_off,
  input         io_dis_uops_0_bits_is_unicore,
  input  [2:0]  io_dis_uops_0_bits_shift,
  input  [1:0]  io_dis_uops_0_bits_lrs3_rtype,
  input         io_dis_uops_0_bits_rflag,
  input         io_dis_uops_0_bits_wflag,
  input  [3:0]  io_dis_uops_0_bits_prflag,
  input  [3:0]  io_dis_uops_0_bits_pwflag,
  input         io_dis_uops_0_bits_pflag_busy,
  input  [3:0]  io_dis_uops_0_bits_stale_pflag,
  input  [3:0]  io_dis_uops_0_bits_op1_sel,
  input  [3:0]  io_dis_uops_0_bits_op2_sel,
  input  [5:0]  io_dis_uops_0_bits_split_num,
  input  [5:0]  io_dis_uops_0_bits_self_index,
  input  [5:0]  io_dis_uops_0_bits_rob_inst_idx,
  input  [5:0]  io_dis_uops_0_bits_address_num,
  input  [6:0]  io_dis_uops_0_bits_uopc,
  input  [31:0] io_dis_uops_0_bits_inst,
  input  [31:0] io_dis_uops_0_bits_debug_inst,
  input         io_dis_uops_0_bits_is_rvc,
  input  [39:0] io_dis_uops_0_bits_debug_pc,
  input  [2:0]  io_dis_uops_0_bits_iq_type,
  input  [9:0]  io_dis_uops_0_bits_fu_code,
  input  [3:0]  io_dis_uops_0_bits_ctrl_br_type,
  input  [1:0]  io_dis_uops_0_bits_ctrl_op1_sel,
  input  [2:0]  io_dis_uops_0_bits_ctrl_op2_sel,
  input  [2:0]  io_dis_uops_0_bits_ctrl_imm_sel,
  input  [3:0]  io_dis_uops_0_bits_ctrl_op_fcn,
  input         io_dis_uops_0_bits_ctrl_fcn_dw,
  input  [2:0]  io_dis_uops_0_bits_ctrl_csr_cmd,
  input         io_dis_uops_0_bits_ctrl_is_load,
  input         io_dis_uops_0_bits_ctrl_is_sta,
  input         io_dis_uops_0_bits_ctrl_is_std,
  input  [1:0]  io_dis_uops_0_bits_ctrl_op3_sel,
  input  [1:0]  io_dis_uops_0_bits_iw_state,
  input         io_dis_uops_0_bits_iw_p1_poisoned,
  input         io_dis_uops_0_bits_iw_p2_poisoned,
  input         io_dis_uops_0_bits_is_br,
  input         io_dis_uops_0_bits_is_jalr,
  input         io_dis_uops_0_bits_is_jal,
  input         io_dis_uops_0_bits_is_sfb,
  input  [11:0] io_dis_uops_0_bits_br_mask,
  input  [3:0]  io_dis_uops_0_bits_br_tag,
  input  [4:0]  io_dis_uops_0_bits_ftq_idx,
  input         io_dis_uops_0_bits_edge_inst,
  input  [5:0]  io_dis_uops_0_bits_pc_lob,
  input         io_dis_uops_0_bits_taken,
  input  [19:0] io_dis_uops_0_bits_imm_packed,
  input  [11:0] io_dis_uops_0_bits_csr_addr,
  input  [5:0]  io_dis_uops_0_bits_rob_idx,
  input  [4:0]  io_dis_uops_0_bits_ldq_idx,
  input  [4:0]  io_dis_uops_0_bits_stq_idx,
  input  [1:0]  io_dis_uops_0_bits_rxq_idx,
  input  [6:0]  io_dis_uops_0_bits_pdst,
  input  [6:0]  io_dis_uops_0_bits_prs1,
  input  [6:0]  io_dis_uops_0_bits_prs2,
  input  [6:0]  io_dis_uops_0_bits_prs3,
  input  [4:0]  io_dis_uops_0_bits_ppred,
  input         io_dis_uops_0_bits_prs1_busy,
  input         io_dis_uops_0_bits_prs2_busy,
  input         io_dis_uops_0_bits_prs3_busy,
  input         io_dis_uops_0_bits_ppred_busy,
  input  [6:0]  io_dis_uops_0_bits_stale_pdst,
  input         io_dis_uops_0_bits_exception,
  input  [63:0] io_dis_uops_0_bits_exc_cause,
  input         io_dis_uops_0_bits_bypassable,
  input  [4:0]  io_dis_uops_0_bits_mem_cmd,
  input  [1:0]  io_dis_uops_0_bits_mem_size,
  input         io_dis_uops_0_bits_mem_signed,
  input         io_dis_uops_0_bits_is_fence,
  input         io_dis_uops_0_bits_is_fencei,
  input         io_dis_uops_0_bits_is_amo,
  input         io_dis_uops_0_bits_uses_ldq,
  input         io_dis_uops_0_bits_uses_stq,
  input         io_dis_uops_0_bits_is_sys_pc2epc,
  input         io_dis_uops_0_bits_is_unique,
  input         io_dis_uops_0_bits_flush_on_commit,
  input         io_dis_uops_0_bits_ldst_is_rs1,
  input  [5:0]  io_dis_uops_0_bits_ldst,
  input  [5:0]  io_dis_uops_0_bits_lrs1,
  input  [5:0]  io_dis_uops_0_bits_lrs2,
  input  [5:0]  io_dis_uops_0_bits_lrs3,
  input         io_dis_uops_0_bits_ldst_val,
  input  [1:0]  io_dis_uops_0_bits_dst_rtype,
  input  [1:0]  io_dis_uops_0_bits_lrs1_rtype,
  input  [1:0]  io_dis_uops_0_bits_lrs2_rtype,
  input         io_dis_uops_0_bits_frs3_en,
  input         io_dis_uops_0_bits_fp_val,
  input         io_dis_uops_0_bits_fp_single,
  input         io_dis_uops_0_bits_xcpt_pf_if,
  input         io_dis_uops_0_bits_xcpt_ae_if,
  input         io_dis_uops_0_bits_xcpt_ma_if,
  input         io_dis_uops_0_bits_bp_debug_if,
  input         io_dis_uops_0_bits_bp_xcpt_if,
  input  [1:0]  io_dis_uops_0_bits_debug_fsrc,
  input  [1:0]  io_dis_uops_0_bits_debug_tsrc,
  output        io_dis_uops_1_ready,
  input         io_dis_uops_1_valid,
  input         io_dis_uops_1_bits_switch,
  input         io_dis_uops_1_bits_switch_off,
  input         io_dis_uops_1_bits_is_unicore,
  input  [2:0]  io_dis_uops_1_bits_shift,
  input  [1:0]  io_dis_uops_1_bits_lrs3_rtype,
  input         io_dis_uops_1_bits_rflag,
  input         io_dis_uops_1_bits_wflag,
  input  [3:0]  io_dis_uops_1_bits_prflag,
  input  [3:0]  io_dis_uops_1_bits_pwflag,
  input         io_dis_uops_1_bits_pflag_busy,
  input  [3:0]  io_dis_uops_1_bits_stale_pflag,
  input  [3:0]  io_dis_uops_1_bits_op1_sel,
  input  [3:0]  io_dis_uops_1_bits_op2_sel,
  input  [5:0]  io_dis_uops_1_bits_split_num,
  input  [5:0]  io_dis_uops_1_bits_self_index,
  input  [5:0]  io_dis_uops_1_bits_rob_inst_idx,
  input  [5:0]  io_dis_uops_1_bits_address_num,
  input  [6:0]  io_dis_uops_1_bits_uopc,
  input  [31:0] io_dis_uops_1_bits_inst,
  input  [31:0] io_dis_uops_1_bits_debug_inst,
  input         io_dis_uops_1_bits_is_rvc,
  input  [39:0] io_dis_uops_1_bits_debug_pc,
  input  [2:0]  io_dis_uops_1_bits_iq_type,
  input  [9:0]  io_dis_uops_1_bits_fu_code,
  input  [3:0]  io_dis_uops_1_bits_ctrl_br_type,
  input  [1:0]  io_dis_uops_1_bits_ctrl_op1_sel,
  input  [2:0]  io_dis_uops_1_bits_ctrl_op2_sel,
  input  [2:0]  io_dis_uops_1_bits_ctrl_imm_sel,
  input  [3:0]  io_dis_uops_1_bits_ctrl_op_fcn,
  input         io_dis_uops_1_bits_ctrl_fcn_dw,
  input  [2:0]  io_dis_uops_1_bits_ctrl_csr_cmd,
  input         io_dis_uops_1_bits_ctrl_is_load,
  input         io_dis_uops_1_bits_ctrl_is_sta,
  input         io_dis_uops_1_bits_ctrl_is_std,
  input  [1:0]  io_dis_uops_1_bits_ctrl_op3_sel,
  input  [1:0]  io_dis_uops_1_bits_iw_state,
  input         io_dis_uops_1_bits_iw_p1_poisoned,
  input         io_dis_uops_1_bits_iw_p2_poisoned,
  input         io_dis_uops_1_bits_is_br,
  input         io_dis_uops_1_bits_is_jalr,
  input         io_dis_uops_1_bits_is_jal,
  input         io_dis_uops_1_bits_is_sfb,
  input  [11:0] io_dis_uops_1_bits_br_mask,
  input  [3:0]  io_dis_uops_1_bits_br_tag,
  input  [4:0]  io_dis_uops_1_bits_ftq_idx,
  input         io_dis_uops_1_bits_edge_inst,
  input  [5:0]  io_dis_uops_1_bits_pc_lob,
  input         io_dis_uops_1_bits_taken,
  input  [19:0] io_dis_uops_1_bits_imm_packed,
  input  [11:0] io_dis_uops_1_bits_csr_addr,
  input  [5:0]  io_dis_uops_1_bits_rob_idx,
  input  [4:0]  io_dis_uops_1_bits_ldq_idx,
  input  [4:0]  io_dis_uops_1_bits_stq_idx,
  input  [1:0]  io_dis_uops_1_bits_rxq_idx,
  input  [6:0]  io_dis_uops_1_bits_pdst,
  input  [6:0]  io_dis_uops_1_bits_prs1,
  input  [6:0]  io_dis_uops_1_bits_prs2,
  input  [6:0]  io_dis_uops_1_bits_prs3,
  input  [4:0]  io_dis_uops_1_bits_ppred,
  input         io_dis_uops_1_bits_prs1_busy,
  input         io_dis_uops_1_bits_prs2_busy,
  input         io_dis_uops_1_bits_prs3_busy,
  input         io_dis_uops_1_bits_ppred_busy,
  input  [6:0]  io_dis_uops_1_bits_stale_pdst,
  input         io_dis_uops_1_bits_exception,
  input  [63:0] io_dis_uops_1_bits_exc_cause,
  input         io_dis_uops_1_bits_bypassable,
  input  [4:0]  io_dis_uops_1_bits_mem_cmd,
  input  [1:0]  io_dis_uops_1_bits_mem_size,
  input         io_dis_uops_1_bits_mem_signed,
  input         io_dis_uops_1_bits_is_fence,
  input         io_dis_uops_1_bits_is_fencei,
  input         io_dis_uops_1_bits_is_amo,
  input         io_dis_uops_1_bits_uses_ldq,
  input         io_dis_uops_1_bits_uses_stq,
  input         io_dis_uops_1_bits_is_sys_pc2epc,
  input         io_dis_uops_1_bits_is_unique,
  input         io_dis_uops_1_bits_flush_on_commit,
  input         io_dis_uops_1_bits_ldst_is_rs1,
  input  [5:0]  io_dis_uops_1_bits_ldst,
  input  [5:0]  io_dis_uops_1_bits_lrs1,
  input  [5:0]  io_dis_uops_1_bits_lrs2,
  input  [5:0]  io_dis_uops_1_bits_lrs3,
  input         io_dis_uops_1_bits_ldst_val,
  input  [1:0]  io_dis_uops_1_bits_dst_rtype,
  input  [1:0]  io_dis_uops_1_bits_lrs1_rtype,
  input  [1:0]  io_dis_uops_1_bits_lrs2_rtype,
  input         io_dis_uops_1_bits_frs3_en,
  input         io_dis_uops_1_bits_fp_val,
  input         io_dis_uops_1_bits_fp_single,
  input         io_dis_uops_1_bits_xcpt_pf_if,
  input         io_dis_uops_1_bits_xcpt_ae_if,
  input         io_dis_uops_1_bits_xcpt_ma_if,
  input         io_dis_uops_1_bits_bp_debug_if,
  input         io_dis_uops_1_bits_bp_xcpt_if,
  input  [1:0]  io_dis_uops_1_bits_debug_fsrc,
  input  [1:0]  io_dis_uops_1_bits_debug_tsrc,
  output        io_iss_valids_0,
  output        io_iss_uops_0_switch,
  output        io_iss_uops_0_switch_off,
  output        io_iss_uops_0_is_unicore,
  output [2:0]  io_iss_uops_0_shift,
  output [1:0]  io_iss_uops_0_lrs3_rtype,
  output        io_iss_uops_0_rflag,
  output        io_iss_uops_0_wflag,
  output [3:0]  io_iss_uops_0_prflag,
  output [3:0]  io_iss_uops_0_pwflag,
  output        io_iss_uops_0_pflag_busy,
  output [3:0]  io_iss_uops_0_stale_pflag,
  output [3:0]  io_iss_uops_0_op1_sel,
  output [3:0]  io_iss_uops_0_op2_sel,
  output [5:0]  io_iss_uops_0_split_num,
  output [5:0]  io_iss_uops_0_self_index,
  output [5:0]  io_iss_uops_0_rob_inst_idx,
  output [5:0]  io_iss_uops_0_address_num,
  output [6:0]  io_iss_uops_0_uopc,
  output [31:0] io_iss_uops_0_inst,
  output [31:0] io_iss_uops_0_debug_inst,
  output        io_iss_uops_0_is_rvc,
  output [39:0] io_iss_uops_0_debug_pc,
  output [2:0]  io_iss_uops_0_iq_type,
  output [9:0]  io_iss_uops_0_fu_code,
  output [3:0]  io_iss_uops_0_ctrl_br_type,
  output [1:0]  io_iss_uops_0_ctrl_op1_sel,
  output [2:0]  io_iss_uops_0_ctrl_op2_sel,
  output [2:0]  io_iss_uops_0_ctrl_imm_sel,
  output [3:0]  io_iss_uops_0_ctrl_op_fcn,
  output        io_iss_uops_0_ctrl_fcn_dw,
  output [2:0]  io_iss_uops_0_ctrl_csr_cmd,
  output        io_iss_uops_0_ctrl_is_load,
  output        io_iss_uops_0_ctrl_is_sta,
  output        io_iss_uops_0_ctrl_is_std,
  output [1:0]  io_iss_uops_0_ctrl_op3_sel,
  output [1:0]  io_iss_uops_0_iw_state,
  output        io_iss_uops_0_iw_p1_poisoned,
  output        io_iss_uops_0_iw_p2_poisoned,
  output        io_iss_uops_0_is_br,
  output        io_iss_uops_0_is_jalr,
  output        io_iss_uops_0_is_jal,
  output        io_iss_uops_0_is_sfb,
  output [11:0] io_iss_uops_0_br_mask,
  output [3:0]  io_iss_uops_0_br_tag,
  output [4:0]  io_iss_uops_0_ftq_idx,
  output        io_iss_uops_0_edge_inst,
  output [5:0]  io_iss_uops_0_pc_lob,
  output        io_iss_uops_0_taken,
  output [19:0] io_iss_uops_0_imm_packed,
  output [11:0] io_iss_uops_0_csr_addr,
  output [5:0]  io_iss_uops_0_rob_idx,
  output [4:0]  io_iss_uops_0_ldq_idx,
  output [4:0]  io_iss_uops_0_stq_idx,
  output [1:0]  io_iss_uops_0_rxq_idx,
  output [6:0]  io_iss_uops_0_pdst,
  output [6:0]  io_iss_uops_0_prs1,
  output [6:0]  io_iss_uops_0_prs2,
  output [6:0]  io_iss_uops_0_prs3,
  output [4:0]  io_iss_uops_0_ppred,
  output        io_iss_uops_0_prs1_busy,
  output        io_iss_uops_0_prs2_busy,
  output        io_iss_uops_0_prs3_busy,
  output        io_iss_uops_0_ppred_busy,
  output [6:0]  io_iss_uops_0_stale_pdst,
  output        io_iss_uops_0_exception,
  output [63:0] io_iss_uops_0_exc_cause,
  output        io_iss_uops_0_bypassable,
  output [4:0]  io_iss_uops_0_mem_cmd,
  output [1:0]  io_iss_uops_0_mem_size,
  output        io_iss_uops_0_mem_signed,
  output        io_iss_uops_0_is_fence,
  output        io_iss_uops_0_is_fencei,
  output        io_iss_uops_0_is_amo,
  output        io_iss_uops_0_uses_ldq,
  output        io_iss_uops_0_uses_stq,
  output        io_iss_uops_0_is_sys_pc2epc,
  output        io_iss_uops_0_is_unique,
  output        io_iss_uops_0_flush_on_commit,
  output        io_iss_uops_0_ldst_is_rs1,
  output [5:0]  io_iss_uops_0_ldst,
  output [5:0]  io_iss_uops_0_lrs1,
  output [5:0]  io_iss_uops_0_lrs2,
  output [5:0]  io_iss_uops_0_lrs3,
  output        io_iss_uops_0_ldst_val,
  output [1:0]  io_iss_uops_0_dst_rtype,
  output [1:0]  io_iss_uops_0_lrs1_rtype,
  output [1:0]  io_iss_uops_0_lrs2_rtype,
  output        io_iss_uops_0_frs3_en,
  output        io_iss_uops_0_fp_val,
  output        io_iss_uops_0_fp_single,
  output        io_iss_uops_0_xcpt_pf_if,
  output        io_iss_uops_0_xcpt_ae_if,
  output        io_iss_uops_0_xcpt_ma_if,
  output        io_iss_uops_0_bp_debug_if,
  output        io_iss_uops_0_bp_xcpt_if,
  output [1:0]  io_iss_uops_0_debug_fsrc,
  output [1:0]  io_iss_uops_0_debug_tsrc,
  input         io_wakeup_ports_0_valid,
  input  [6:0]  io_wakeup_ports_0_bits_pdst,
  input         io_wakeup_ports_0_bits_poisoned,
  input  [6:0]  io_wakeup_ports_0_bits_pwflag,
  input         io_wakeup_ports_0_bits_flag_valid,
  input         io_wakeup_ports_1_valid,
  input  [6:0]  io_wakeup_ports_1_bits_pdst,
  input         io_wakeup_ports_1_bits_poisoned,
  input  [6:0]  io_wakeup_ports_1_bits_pwflag,
  input         io_wakeup_ports_1_bits_flag_valid,
  input         io_pred_wakeup_port_valid,
  input  [4:0]  io_pred_wakeup_port_bits,
  input         io_spec_ld_wakeup_0_valid,
  input  [6:0]  io_spec_ld_wakeup_0_bits,
  input  [9:0]  io_fu_types_0,
  input  [11:0] io_brupdate_b1_resolve_mask,
  input  [11:0] io_brupdate_b1_mispredict_mask,
  input         io_brupdate_b2_uop_switch,
  input         io_brupdate_b2_uop_switch_off,
  input         io_brupdate_b2_uop_is_unicore,
  input  [2:0]  io_brupdate_b2_uop_shift,
  input  [1:0]  io_brupdate_b2_uop_lrs3_rtype,
  input         io_brupdate_b2_uop_rflag,
  input         io_brupdate_b2_uop_wflag,
  input  [3:0]  io_brupdate_b2_uop_prflag,
  input  [3:0]  io_brupdate_b2_uop_pwflag,
  input         io_brupdate_b2_uop_pflag_busy,
  input  [3:0]  io_brupdate_b2_uop_stale_pflag,
  input  [3:0]  io_brupdate_b2_uop_op1_sel,
  input  [3:0]  io_brupdate_b2_uop_op2_sel,
  input  [5:0]  io_brupdate_b2_uop_split_num,
  input  [5:0]  io_brupdate_b2_uop_self_index,
  input  [5:0]  io_brupdate_b2_uop_rob_inst_idx,
  input  [5:0]  io_brupdate_b2_uop_address_num,
  input  [6:0]  io_brupdate_b2_uop_uopc,
  input  [31:0] io_brupdate_b2_uop_inst,
  input  [31:0] io_brupdate_b2_uop_debug_inst,
  input         io_brupdate_b2_uop_is_rvc,
  input  [39:0] io_brupdate_b2_uop_debug_pc,
  input  [2:0]  io_brupdate_b2_uop_iq_type,
  input  [9:0]  io_brupdate_b2_uop_fu_code,
  input  [3:0]  io_brupdate_b2_uop_ctrl_br_type,
  input  [1:0]  io_brupdate_b2_uop_ctrl_op1_sel,
  input  [2:0]  io_brupdate_b2_uop_ctrl_op2_sel,
  input  [2:0]  io_brupdate_b2_uop_ctrl_imm_sel,
  input  [3:0]  io_brupdate_b2_uop_ctrl_op_fcn,
  input         io_brupdate_b2_uop_ctrl_fcn_dw,
  input  [2:0]  io_brupdate_b2_uop_ctrl_csr_cmd,
  input         io_brupdate_b2_uop_ctrl_is_load,
  input         io_brupdate_b2_uop_ctrl_is_sta,
  input         io_brupdate_b2_uop_ctrl_is_std,
  input  [1:0]  io_brupdate_b2_uop_ctrl_op3_sel,
  input  [1:0]  io_brupdate_b2_uop_iw_state,
  input         io_brupdate_b2_uop_iw_p1_poisoned,
  input         io_brupdate_b2_uop_iw_p2_poisoned,
  input         io_brupdate_b2_uop_is_br,
  input         io_brupdate_b2_uop_is_jalr,
  input         io_brupdate_b2_uop_is_jal,
  input         io_brupdate_b2_uop_is_sfb,
  input  [11:0] io_brupdate_b2_uop_br_mask,
  input  [3:0]  io_brupdate_b2_uop_br_tag,
  input  [4:0]  io_brupdate_b2_uop_ftq_idx,
  input         io_brupdate_b2_uop_edge_inst,
  input  [5:0]  io_brupdate_b2_uop_pc_lob,
  input         io_brupdate_b2_uop_taken,
  input  [19:0] io_brupdate_b2_uop_imm_packed,
  input  [11:0] io_brupdate_b2_uop_csr_addr,
  input  [5:0]  io_brupdate_b2_uop_rob_idx,
  input  [4:0]  io_brupdate_b2_uop_ldq_idx,
  input  [4:0]  io_brupdate_b2_uop_stq_idx,
  input  [1:0]  io_brupdate_b2_uop_rxq_idx,
  input  [6:0]  io_brupdate_b2_uop_pdst,
  input  [6:0]  io_brupdate_b2_uop_prs1,
  input  [6:0]  io_brupdate_b2_uop_prs2,
  input  [6:0]  io_brupdate_b2_uop_prs3,
  input  [4:0]  io_brupdate_b2_uop_ppred,
  input         io_brupdate_b2_uop_prs1_busy,
  input         io_brupdate_b2_uop_prs2_busy,
  input         io_brupdate_b2_uop_prs3_busy,
  input         io_brupdate_b2_uop_ppred_busy,
  input  [6:0]  io_brupdate_b2_uop_stale_pdst,
  input         io_brupdate_b2_uop_exception,
  input  [63:0] io_brupdate_b2_uop_exc_cause,
  input         io_brupdate_b2_uop_bypassable,
  input  [4:0]  io_brupdate_b2_uop_mem_cmd,
  input  [1:0]  io_brupdate_b2_uop_mem_size,
  input         io_brupdate_b2_uop_mem_signed,
  input         io_brupdate_b2_uop_is_fence,
  input         io_brupdate_b2_uop_is_fencei,
  input         io_brupdate_b2_uop_is_amo,
  input         io_brupdate_b2_uop_uses_ldq,
  input         io_brupdate_b2_uop_uses_stq,
  input         io_brupdate_b2_uop_is_sys_pc2epc,
  input         io_brupdate_b2_uop_is_unique,
  input         io_brupdate_b2_uop_flush_on_commit,
  input         io_brupdate_b2_uop_ldst_is_rs1,
  input  [5:0]  io_brupdate_b2_uop_ldst,
  input  [5:0]  io_brupdate_b2_uop_lrs1,
  input  [5:0]  io_brupdate_b2_uop_lrs2,
  input  [5:0]  io_brupdate_b2_uop_lrs3,
  input         io_brupdate_b2_uop_ldst_val,
  input  [1:0]  io_brupdate_b2_uop_dst_rtype,
  input  [1:0]  io_brupdate_b2_uop_lrs1_rtype,
  input  [1:0]  io_brupdate_b2_uop_lrs2_rtype,
  input         io_brupdate_b2_uop_frs3_en,
  input         io_brupdate_b2_uop_fp_val,
  input         io_brupdate_b2_uop_fp_single,
  input         io_brupdate_b2_uop_xcpt_pf_if,
  input         io_brupdate_b2_uop_xcpt_ae_if,
  input         io_brupdate_b2_uop_xcpt_ma_if,
  input         io_brupdate_b2_uop_bp_debug_if,
  input         io_brupdate_b2_uop_bp_xcpt_if,
  input  [1:0]  io_brupdate_b2_uop_debug_fsrc,
  input  [1:0]  io_brupdate_b2_uop_debug_tsrc,
  input         io_brupdate_b2_valid,
  input         io_brupdate_b2_mispredict,
  input         io_brupdate_b2_taken,
  input  [2:0]  io_brupdate_b2_cfi_type,
  input  [1:0]  io_brupdate_b2_pc_sel,
  input  [39:0] io_brupdate_b2_jalr_target,
  input  [31:0] io_brupdate_b2_target_offset,
  input         io_flush_pipeline,
  input         io_ld_miss,
  output        io_event_empty,
  input  [63:0] io_tsc_reg
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  slots_0_clock; // @[issue-unit.scala 157:73]
  wire  slots_0_reset; // @[issue-unit.scala 157:73]
  wire  slots_0_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_0_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_0_io_request; // @[issue-unit.scala 157:73]
  wire  slots_0_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_0_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_0_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_0_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_0_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_0_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_0_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_0_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_0_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_0_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_0_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_0_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_0_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_0_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_0_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_0_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_0_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_0_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_0_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_0_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_0_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_0_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_0_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_0_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_0_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_0_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_0_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_0_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_0_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_0_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_0_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_0_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_0_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_0_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_0_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_0_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_0_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_0_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_0_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_0_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_0_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_0_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_0_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_0_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_0_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_0_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_0_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_0_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_0_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_0_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_0_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_0_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_0_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_0_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_0_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_0_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_0_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_1_clock; // @[issue-unit.scala 157:73]
  wire  slots_1_reset; // @[issue-unit.scala 157:73]
  wire  slots_1_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_1_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_1_io_request; // @[issue-unit.scala 157:73]
  wire  slots_1_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_1_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_1_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_1_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_1_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_1_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_1_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_1_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_1_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_1_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_1_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_1_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_1_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_1_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_1_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_1_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_1_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_1_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_1_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_1_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_1_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_1_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_1_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_1_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_1_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_1_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_1_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_1_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_1_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_1_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_1_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_1_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_1_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_1_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_1_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_1_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_1_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_1_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_1_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_1_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_1_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_1_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_1_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_1_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_1_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_1_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_1_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_1_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_1_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_1_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_1_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_1_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_1_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_1_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_1_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_1_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_1_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_2_clock; // @[issue-unit.scala 157:73]
  wire  slots_2_reset; // @[issue-unit.scala 157:73]
  wire  slots_2_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_2_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_2_io_request; // @[issue-unit.scala 157:73]
  wire  slots_2_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_2_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_2_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_2_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_2_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_2_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_2_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_2_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_2_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_2_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_2_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_2_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_2_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_2_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_2_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_2_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_2_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_2_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_2_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_2_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_2_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_2_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_2_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_2_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_2_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_2_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_2_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_2_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_2_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_2_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_2_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_2_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_2_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_2_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_2_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_2_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_2_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_2_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_2_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_2_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_2_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_2_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_2_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_2_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_2_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_2_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_2_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_2_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_2_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_2_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_2_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_2_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_2_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_2_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_2_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_2_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_2_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_3_clock; // @[issue-unit.scala 157:73]
  wire  slots_3_reset; // @[issue-unit.scala 157:73]
  wire  slots_3_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_3_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_3_io_request; // @[issue-unit.scala 157:73]
  wire  slots_3_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_3_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_3_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_3_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_3_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_3_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_3_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_3_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_3_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_3_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_3_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_3_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_3_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_3_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_3_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_3_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_3_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_3_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_3_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_3_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_3_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_3_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_3_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_3_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_3_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_3_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_3_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_3_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_3_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_3_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_3_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_3_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_3_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_3_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_3_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_3_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_3_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_3_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_3_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_3_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_3_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_3_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_3_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_3_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_3_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_3_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_3_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_3_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_3_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_3_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_3_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_3_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_3_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_3_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_3_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_3_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_3_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_4_clock; // @[issue-unit.scala 157:73]
  wire  slots_4_reset; // @[issue-unit.scala 157:73]
  wire  slots_4_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_4_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_4_io_request; // @[issue-unit.scala 157:73]
  wire  slots_4_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_4_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_4_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_4_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_4_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_4_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_4_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_4_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_4_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_4_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_4_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_4_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_4_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_4_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_4_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_4_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_4_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_4_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_4_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_4_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_4_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_4_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_4_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_4_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_4_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_4_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_4_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_4_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_4_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_4_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_4_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_4_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_4_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_4_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_4_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_4_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_4_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_4_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_4_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_4_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_4_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_4_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_4_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_4_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_4_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_4_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_4_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_4_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_4_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_4_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_4_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_4_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_4_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_4_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_4_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_4_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_4_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_5_clock; // @[issue-unit.scala 157:73]
  wire  slots_5_reset; // @[issue-unit.scala 157:73]
  wire  slots_5_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_5_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_5_io_request; // @[issue-unit.scala 157:73]
  wire  slots_5_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_5_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_5_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_5_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_5_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_5_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_5_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_5_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_5_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_5_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_5_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_5_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_5_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_5_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_5_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_5_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_5_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_5_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_5_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_5_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_5_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_5_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_5_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_5_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_5_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_5_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_5_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_5_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_5_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_5_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_5_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_5_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_5_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_5_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_5_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_5_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_5_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_5_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_5_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_5_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_5_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_5_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_5_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_5_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_5_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_5_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_5_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_5_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_5_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_5_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_5_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_5_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_5_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_5_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_5_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_5_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_5_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_6_clock; // @[issue-unit.scala 157:73]
  wire  slots_6_reset; // @[issue-unit.scala 157:73]
  wire  slots_6_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_6_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_6_io_request; // @[issue-unit.scala 157:73]
  wire  slots_6_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_6_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_6_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_6_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_6_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_6_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_6_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_6_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_6_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_6_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_6_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_6_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_6_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_6_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_6_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_6_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_6_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_6_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_6_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_6_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_6_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_6_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_6_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_6_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_6_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_6_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_6_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_6_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_6_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_6_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_6_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_6_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_6_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_6_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_6_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_6_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_6_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_6_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_6_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_6_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_6_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_6_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_6_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_6_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_6_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_6_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_6_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_6_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_6_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_6_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_6_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_6_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_6_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_6_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_6_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_6_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_6_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_7_clock; // @[issue-unit.scala 157:73]
  wire  slots_7_reset; // @[issue-unit.scala 157:73]
  wire  slots_7_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_7_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_7_io_request; // @[issue-unit.scala 157:73]
  wire  slots_7_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_7_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_7_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_7_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_7_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_7_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_7_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_7_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_7_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_7_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_7_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_7_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_7_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_7_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_7_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_7_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_7_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_7_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_7_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_7_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_7_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_7_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_7_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_7_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_7_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_7_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_7_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_7_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_7_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_7_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_7_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_7_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_7_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_7_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_7_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_7_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_7_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_7_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_7_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_7_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_7_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_7_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_7_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_7_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_7_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_7_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_7_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_7_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_7_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_7_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_7_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_7_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_7_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_7_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_7_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_7_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_7_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_8_clock; // @[issue-unit.scala 157:73]
  wire  slots_8_reset; // @[issue-unit.scala 157:73]
  wire  slots_8_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_8_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_8_io_request; // @[issue-unit.scala 157:73]
  wire  slots_8_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_8_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_8_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_8_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_8_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_8_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_8_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_8_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_8_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_8_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_8_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_8_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_8_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_8_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_8_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_8_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_8_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_8_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_8_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_8_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_8_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_8_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_8_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_8_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_8_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_8_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_8_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_8_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_8_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_8_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_8_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_8_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_8_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_8_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_8_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_8_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_8_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_8_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_8_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_8_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_8_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_8_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_8_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_8_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_8_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_8_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_8_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_8_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_8_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_8_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_8_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_8_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_8_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_8_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_8_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_8_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_8_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_9_clock; // @[issue-unit.scala 157:73]
  wire  slots_9_reset; // @[issue-unit.scala 157:73]
  wire  slots_9_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_9_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_9_io_request; // @[issue-unit.scala 157:73]
  wire  slots_9_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_9_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_9_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_9_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_9_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_9_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_9_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_9_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_9_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_9_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_9_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_9_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_9_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_9_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_9_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_9_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_9_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_9_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_9_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_9_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_9_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_9_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_9_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_9_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_9_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_9_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_9_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_9_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_9_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_9_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_9_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_9_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_9_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_9_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_9_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_9_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_9_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_9_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_9_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_9_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_9_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_9_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_9_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_9_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_9_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_9_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_9_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_9_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_9_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_9_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_9_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_9_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_9_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_9_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_9_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_9_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_9_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_10_clock; // @[issue-unit.scala 157:73]
  wire  slots_10_reset; // @[issue-unit.scala 157:73]
  wire  slots_10_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_10_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_10_io_request; // @[issue-unit.scala 157:73]
  wire  slots_10_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_10_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_10_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_10_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_10_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_10_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_10_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_10_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_10_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_10_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_10_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_10_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_10_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_10_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_10_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_10_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_10_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_10_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_10_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_10_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_10_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_10_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_10_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_10_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_10_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_10_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_10_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_10_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_10_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_10_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_10_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_10_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_10_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_10_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_10_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_10_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_10_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_10_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_10_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_10_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_10_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_10_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_10_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_10_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_10_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_10_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_10_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_10_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_10_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_10_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_10_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_10_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_10_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_10_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_10_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_10_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_10_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_11_clock; // @[issue-unit.scala 157:73]
  wire  slots_11_reset; // @[issue-unit.scala 157:73]
  wire  slots_11_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_11_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_11_io_request; // @[issue-unit.scala 157:73]
  wire  slots_11_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_11_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_11_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_11_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_11_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_11_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_11_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_11_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_11_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_11_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_11_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_11_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_11_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_11_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_11_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_11_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_11_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_11_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_11_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_11_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_11_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_11_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_11_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_11_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_11_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_11_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_11_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_11_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_11_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_11_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_11_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_11_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_11_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_11_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_11_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_11_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_11_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_11_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_11_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_11_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_11_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_11_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_11_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_11_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_11_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_11_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_11_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_11_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_11_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_11_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_11_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_11_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_11_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_11_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_11_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_11_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_11_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_12_clock; // @[issue-unit.scala 157:73]
  wire  slots_12_reset; // @[issue-unit.scala 157:73]
  wire  slots_12_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_12_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_12_io_request; // @[issue-unit.scala 157:73]
  wire  slots_12_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_12_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_12_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_12_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_12_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_12_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_12_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_12_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_12_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_12_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_12_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_12_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_12_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_12_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_12_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_12_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_12_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_12_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_12_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_12_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_12_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_12_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_12_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_12_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_12_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_12_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_12_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_12_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_12_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_12_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_12_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_12_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_12_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_12_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_12_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_12_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_12_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_12_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_12_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_12_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_12_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_12_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_12_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_12_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_12_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_12_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_12_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_12_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_12_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_12_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_12_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_12_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_12_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_12_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_12_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_12_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_12_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_13_clock; // @[issue-unit.scala 157:73]
  wire  slots_13_reset; // @[issue-unit.scala 157:73]
  wire  slots_13_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_13_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_13_io_request; // @[issue-unit.scala 157:73]
  wire  slots_13_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_13_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_13_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_13_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_13_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_13_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_13_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_13_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_13_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_13_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_13_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_13_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_13_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_13_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_13_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_13_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_13_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_13_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_13_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_13_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_13_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_13_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_13_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_13_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_13_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_13_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_13_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_13_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_13_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_13_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_13_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_13_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_13_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_13_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_13_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_13_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_13_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_13_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_13_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_13_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_13_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_13_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_13_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_13_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_13_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_13_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_13_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_13_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_13_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_13_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_13_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_13_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_13_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_13_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_13_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_13_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_13_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_14_clock; // @[issue-unit.scala 157:73]
  wire  slots_14_reset; // @[issue-unit.scala 157:73]
  wire  slots_14_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_14_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_14_io_request; // @[issue-unit.scala 157:73]
  wire  slots_14_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_14_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_14_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_14_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_14_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_14_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_14_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_14_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_14_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_14_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_14_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_14_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_14_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_14_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_14_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_14_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_14_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_14_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_14_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_14_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_14_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_14_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_14_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_14_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_14_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_14_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_14_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_14_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_14_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_14_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_14_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_14_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_14_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_14_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_14_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_14_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_14_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_14_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_14_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_14_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_14_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_14_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_14_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_14_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_14_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_14_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_14_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_14_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_14_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_14_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_14_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_14_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_14_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_14_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_14_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_14_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_14_io_debug_state; // @[issue-unit.scala 157:73]
  wire  slots_15_clock; // @[issue-unit.scala 157:73]
  wire  slots_15_reset; // @[issue-unit.scala 157:73]
  wire  slots_15_io_valid; // @[issue-unit.scala 157:73]
  wire  slots_15_io_will_be_valid; // @[issue-unit.scala 157:73]
  wire  slots_15_io_request; // @[issue-unit.scala 157:73]
  wire  slots_15_io_request_hp; // @[issue-unit.scala 157:73]
  wire  slots_15_io_grant; // @[issue-unit.scala 157:73]
  wire [11:0] slots_15_io_brupdate_b1_resolve_mask; // @[issue-unit.scala 157:73]
  wire [11:0] slots_15_io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_brupdate_b2_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_brupdate_b2_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_brupdate_b2_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_brupdate_b2_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_brupdate_b2_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_brupdate_b2_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_15_io_brupdate_b2_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_15_io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_15_io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_15_io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_15_io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_15_io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_15_io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_brupdate_b2_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_brupdate_b2_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_brupdate_b2_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_brupdate_b2_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_brupdate_b2_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_15_io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_brupdate_b2_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_valid; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_mispredict; // @[issue-unit.scala 157:73]
  wire  slots_15_io_brupdate_b2_taken; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_brupdate_b2_cfi_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_brupdate_b2_pc_sel; // @[issue-unit.scala 157:73]
  wire [39:0] slots_15_io_brupdate_b2_jalr_target; // @[issue-unit.scala 157:73]
  wire [31:0] slots_15_io_brupdate_b2_target_offset; // @[issue-unit.scala 157:73]
  wire  slots_15_io_kill; // @[issue-unit.scala 157:73]
  wire  slots_15_io_clear; // @[issue-unit.scala 157:73]
  wire  slots_15_io_ldspec_miss; // @[issue-unit.scala 157:73]
  wire  slots_15_io_wakeup_ports_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_15_io_wakeup_ports_1_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 157:73]
  wire  slots_15_io_pred_wakeup_port_valid; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_pred_wakeup_port_bits; // @[issue-unit.scala 157:73]
  wire  slots_15_io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_valid; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_switch; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_in_uop_bits_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_rflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_in_uop_bits_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_in_uop_bits_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_in_uop_bits_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_in_uop_bits_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_in_uop_bits_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_in_uop_bits_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_in_uop_bits_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_in_uop_bits_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_in_uop_bits_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_in_uop_bits_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_15_io_in_uop_bits_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_15_io_in_uop_bits_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_15_io_in_uop_bits_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_in_uop_bits_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_15_io_in_uop_bits_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_in_uop_bits_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_in_uop_bits_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_in_uop_bits_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_in_uop_bits_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_in_uop_bits_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_br; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_15_io_in_uop_bits_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_in_uop_bits_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_in_uop_bits_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_in_uop_bits_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_15_io_in_uop_bits_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_15_io_in_uop_bits_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_in_uop_bits_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_in_uop_bits_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_in_uop_bits_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_in_uop_bits_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_in_uop_bits_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_in_uop_bits_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_in_uop_bits_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_in_uop_bits_ppred; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_in_uop_bits_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_15_io_in_uop_bits_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_in_uop_bits_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_in_uop_bits_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_in_uop_bits_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_in_uop_bits_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_in_uop_bits_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_in_uop_bits_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_in_uop_bits_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_out_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_out_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_out_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_out_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_out_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_out_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_out_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_out_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_out_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_out_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_out_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_15_io_out_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_15_io_out_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_15_io_out_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_out_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_15_io_out_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_out_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_15_io_out_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_out_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_out_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_out_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_15_io_out_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_15_io_out_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_out_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_out_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_out_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_out_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_out_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_out_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_out_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_out_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_out_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_15_io_out_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_out_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_out_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_out_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_out_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_out_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_out_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_switch; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_switch_off; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_unicore; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_uop_shift; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_lrs3_rtype; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_rflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_wflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_uop_prflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_uop_pwflag; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_pflag_busy; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_uop_stale_pflag; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_uop_op1_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_uop_op2_sel; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_uop_split_num; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_uop_self_index; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_uop_rob_inst_idx; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_uop_address_num; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_uop_uopc; // @[issue-unit.scala 157:73]
  wire [31:0] slots_15_io_uop_inst; // @[issue-unit.scala 157:73]
  wire [31:0] slots_15_io_uop_debug_inst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_rvc; // @[issue-unit.scala 157:73]
  wire [39:0] slots_15_io_uop_debug_pc; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_uop_iq_type; // @[issue-unit.scala 157:73]
  wire [9:0] slots_15_io_uop_fu_code; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_uop_ctrl_br_type; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_ctrl_op1_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_uop_ctrl_op2_sel; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_uop_ctrl_imm_sel; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_uop_ctrl_op_fcn; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 157:73]
  wire [2:0] slots_15_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_ctrl_is_load; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_ctrl_is_sta; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_ctrl_is_std; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_ctrl_op3_sel; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_iw_state; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_iw_p1_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_iw_p2_poisoned; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_br; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_jalr; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_jal; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_sfb; // @[issue-unit.scala 157:73]
  wire [11:0] slots_15_io_uop_br_mask; // @[issue-unit.scala 157:73]
  wire [3:0] slots_15_io_uop_br_tag; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_uop_ftq_idx; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_edge_inst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_uop_pc_lob; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_taken; // @[issue-unit.scala 157:73]
  wire [19:0] slots_15_io_uop_imm_packed; // @[issue-unit.scala 157:73]
  wire [11:0] slots_15_io_uop_csr_addr; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_uop_rob_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_uop_ldq_idx; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_uop_stq_idx; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_rxq_idx; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_uop_pdst; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_uop_prs1; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_uop_prs2; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_uop_prs3; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_uop_ppred; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_prs1_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_prs2_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_prs3_busy; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_ppred_busy; // @[issue-unit.scala 157:73]
  wire [6:0] slots_15_io_uop_stale_pdst; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_exception; // @[issue-unit.scala 157:73]
  wire [63:0] slots_15_io_uop_exc_cause; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_bypassable; // @[issue-unit.scala 157:73]
  wire [4:0] slots_15_io_uop_mem_cmd; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_mem_size; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_mem_signed; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_fence; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_fencei; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_amo; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_uses_ldq; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_uses_stq; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_sys_pc2epc; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_is_unique; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_flush_on_commit; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_ldst_is_rs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_uop_ldst; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_uop_lrs1; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_uop_lrs2; // @[issue-unit.scala 157:73]
  wire [5:0] slots_15_io_uop_lrs3; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_ldst_val; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_dst_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_lrs1_rtype; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_lrs2_rtype; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_frs3_en; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_fp_val; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_fp_single; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_xcpt_pf_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_xcpt_ae_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_xcpt_ma_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_bp_debug_if; // @[issue-unit.scala 157:73]
  wire  slots_15_io_uop_bp_xcpt_if; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_debug_fsrc; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_uop_debug_tsrc; // @[issue-unit.scala 157:73]
  wire  slots_15_io_debug_p1; // @[issue-unit.scala 157:73]
  wire  slots_15_io_debug_p2; // @[issue-unit.scala 157:73]
  wire  slots_15_io_debug_p3; // @[issue-unit.scala 157:73]
  wire  slots_15_io_debug_ppred; // @[issue-unit.scala 157:73]
  wire [1:0] slots_15_io_debug_state; // @[issue-unit.scala 157:73]
  wire [1:0] uops_16_lrs1_rtype = io_dis_uops_0_bits_uopc == 7'h2 ? 2'h2 : io_dis_uops_0_bits_lrs1_rtype; // @[issue-unit.scala 142:50 issue-unit.scala 143:32 issue-unit.scala 124:17]
  wire  uops_16_prs1_busy = io_dis_uops_0_bits_uopc == 7'h2 ? 1'h0 : io_dis_uops_0_bits_prs1_busy; // @[issue-unit.scala 142:50 issue-unit.scala 144:32 issue-unit.scala 124:17]
  wire [1:0] uops_17_lrs1_rtype = io_dis_uops_1_bits_uopc == 7'h2 ? 2'h2 : io_dis_uops_1_bits_lrs1_rtype; // @[issue-unit.scala 142:50 issue-unit.scala 143:32 issue-unit.scala 124:17]
  wire  uops_17_prs1_busy = io_dis_uops_1_bits_uopc == 7'h2 ? 1'h0 : io_dis_uops_1_bits_prs1_busy; // @[issue-unit.scala 142:50 issue-unit.scala 144:32 issue-unit.scala 124:17]
  wire  issue_slots_0_valid = slots_0_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_valid = slots_1_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_valid = slots_2_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_valid = slots_3_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_valid = slots_4_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_valid = slots_5_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_valid = slots_6_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_valid = slots_7_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_valid = slots_8_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_valid = slots_9_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_valid = slots_10_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_valid = slots_11_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_valid = slots_12_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_valid = slots_13_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_valid = slots_14_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_valid = slots_15_io_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_0_request = slots_0_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_0_uop_fu_code = slots_0_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_332 = issue_slots_0_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_333 = _T_332 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  issue_slots_0_grant = issue_slots_0_request & _T_333; // @[issue-unit-age-ordered.scala 122:40]
  wire  issue_slots_1_request = slots_1_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_1_uop_fu_code = slots_1_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_347 = issue_slots_1_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_348 = _T_347 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_351 = issue_slots_1_request & _T_348; // @[issue-unit-age-ordered.scala 122:40]
  wire  issue_slots_1_grant = issue_slots_1_request & _T_348 & ~issue_slots_0_grant; // @[issue-unit-age-ordered.scala 122:56]
  wire [1:0] _T_57 = issue_slots_0_grant + issue_slots_1_grant; // @[Bitwise.scala 47:55]
  wire  issue_slots_2_request = slots_2_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_2_uop_fu_code = slots_2_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_362 = issue_slots_2_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_363 = _T_362 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_366 = issue_slots_2_request & _T_363; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_357 = _T_351 | issue_slots_0_grant; // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_2_grant = issue_slots_2_request & _T_363 & ~_T_357; // @[issue-unit-age-ordered.scala 122:56]
  wire  issue_slots_3_request = slots_3_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_3_uop_fu_code = slots_3_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_377 = issue_slots_3_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_378 = _T_377 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_381 = issue_slots_3_request & _T_378; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_372 = _T_366 | (_T_351 | issue_slots_0_grant); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_3_grant = issue_slots_3_request & _T_378 & ~_T_372; // @[issue-unit-age-ordered.scala 122:56]
  wire [1:0] _T_59 = issue_slots_2_grant + issue_slots_3_grant; // @[Bitwise.scala 47:55]
  wire [2:0] _T_61 = _T_57 + _T_59; // @[Bitwise.scala 47:55]
  wire  issue_slots_4_request = slots_4_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_4_uop_fu_code = slots_4_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_392 = issue_slots_4_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_393 = _T_392 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_396 = issue_slots_4_request & _T_393; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_387 = _T_381 | (_T_366 | (_T_351 | issue_slots_0_grant)); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_4_grant = issue_slots_4_request & _T_393 & ~_T_387; // @[issue-unit-age-ordered.scala 122:56]
  wire  issue_slots_5_request = slots_5_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_5_uop_fu_code = slots_5_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_407 = issue_slots_5_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_408 = _T_407 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_411 = issue_slots_5_request & _T_408; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_402 = _T_396 | (_T_381 | (_T_366 | (_T_351 | issue_slots_0_grant))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_5_grant = issue_slots_5_request & _T_408 & ~_T_402; // @[issue-unit-age-ordered.scala 122:56]
  wire [1:0] _T_63 = issue_slots_4_grant + issue_slots_5_grant; // @[Bitwise.scala 47:55]
  wire  issue_slots_6_request = slots_6_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_6_uop_fu_code = slots_6_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_422 = issue_slots_6_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_423 = _T_422 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_426 = issue_slots_6_request & _T_423; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_417 = _T_411 | (_T_396 | (_T_381 | (_T_366 | (_T_351 | issue_slots_0_grant)))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_6_grant = issue_slots_6_request & _T_423 & ~_T_417; // @[issue-unit-age-ordered.scala 122:56]
  wire  issue_slots_7_request = slots_7_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_7_uop_fu_code = slots_7_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_437 = issue_slots_7_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_438 = _T_437 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_441 = issue_slots_7_request & _T_438; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_432 = _T_426 | (_T_411 | (_T_396 | (_T_381 | (_T_366 | (_T_351 | issue_slots_0_grant))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_7_grant = issue_slots_7_request & _T_438 & ~_T_432; // @[issue-unit-age-ordered.scala 122:56]
  wire [1:0] _T_65 = issue_slots_6_grant + issue_slots_7_grant; // @[Bitwise.scala 47:55]
  wire [2:0] _T_67 = _T_63 + _T_65; // @[Bitwise.scala 47:55]
  wire [3:0] _T_69 = _T_61 + _T_67; // @[Bitwise.scala 47:55]
  wire  issue_slots_8_request = slots_8_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_8_uop_fu_code = slots_8_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_452 = issue_slots_8_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_453 = _T_452 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_456 = issue_slots_8_request & _T_453; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_447 = _T_441 | (_T_426 | (_T_411 | (_T_396 | (_T_381 | (_T_366 | (_T_351 | issue_slots_0_grant)))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_8_grant = issue_slots_8_request & _T_453 & ~_T_447; // @[issue-unit-age-ordered.scala 122:56]
  wire  issue_slots_9_request = slots_9_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_9_uop_fu_code = slots_9_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_467 = issue_slots_9_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_468 = _T_467 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_471 = issue_slots_9_request & _T_468; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_462 = _T_456 | (_T_441 | (_T_426 | (_T_411 | (_T_396 | (_T_381 | (_T_366 | (_T_351 | issue_slots_0_grant)))))
    )); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_9_grant = issue_slots_9_request & _T_468 & ~_T_462; // @[issue-unit-age-ordered.scala 122:56]
  wire [1:0] _T_71 = issue_slots_8_grant + issue_slots_9_grant; // @[Bitwise.scala 47:55]
  wire  issue_slots_10_request = slots_10_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_10_uop_fu_code = slots_10_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_482 = issue_slots_10_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_483 = _T_482 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_486 = issue_slots_10_request & _T_483; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_477 = _T_471 | (_T_456 | (_T_441 | (_T_426 | (_T_411 | (_T_396 | (_T_381 | (_T_366 | (_T_351 |
    issue_slots_0_grant)))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_10_grant = issue_slots_10_request & _T_483 & ~_T_477; // @[issue-unit-age-ordered.scala 122:56]
  wire  issue_slots_11_request = slots_11_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_11_uop_fu_code = slots_11_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_497 = issue_slots_11_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_498 = _T_497 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_501 = issue_slots_11_request & _T_498; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_492 = _T_486 | (_T_471 | (_T_456 | (_T_441 | (_T_426 | (_T_411 | (_T_396 | (_T_381 | (_T_366 | (_T_351 |
    issue_slots_0_grant))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_11_grant = issue_slots_11_request & _T_498 & ~_T_492; // @[issue-unit-age-ordered.scala 122:56]
  wire [1:0] _T_73 = issue_slots_10_grant + issue_slots_11_grant; // @[Bitwise.scala 47:55]
  wire [2:0] _T_75 = _T_71 + _T_73; // @[Bitwise.scala 47:55]
  wire  issue_slots_12_request = slots_12_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_12_uop_fu_code = slots_12_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_512 = issue_slots_12_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_513 = _T_512 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_516 = issue_slots_12_request & _T_513; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_507 = _T_501 | (_T_486 | (_T_471 | (_T_456 | (_T_441 | (_T_426 | (_T_411 | (_T_396 | (_T_381 | (_T_366 | (
    _T_351 | issue_slots_0_grant)))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_12_grant = issue_slots_12_request & _T_513 & ~_T_507; // @[issue-unit-age-ordered.scala 122:56]
  wire  issue_slots_13_request = slots_13_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_13_uop_fu_code = slots_13_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_527 = issue_slots_13_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_528 = _T_527 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_531 = issue_slots_13_request & _T_528; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_522 = _T_516 | (_T_501 | (_T_486 | (_T_471 | (_T_456 | (_T_441 | (_T_426 | (_T_411 | (_T_396 | (_T_381 | (
    _T_366 | (_T_351 | issue_slots_0_grant))))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_13_grant = issue_slots_13_request & _T_528 & ~_T_522; // @[issue-unit-age-ordered.scala 122:56]
  wire [1:0] _T_77 = issue_slots_12_grant + issue_slots_13_grant; // @[Bitwise.scala 47:55]
  wire  issue_slots_14_request = slots_14_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_14_uop_fu_code = slots_14_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_542 = issue_slots_14_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_543 = _T_542 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_546 = issue_slots_14_request & _T_543; // @[issue-unit-age-ordered.scala 122:40]
  wire  _T_537 = _T_531 | (_T_516 | (_T_501 | (_T_486 | (_T_471 | (_T_456 | (_T_441 | (_T_426 | (_T_411 | (_T_396 | (
    _T_381 | (_T_366 | (_T_351 | issue_slots_0_grant)))))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_14_grant = issue_slots_14_request & _T_543 & ~_T_537; // @[issue-unit-age-ordered.scala 122:56]
  wire  issue_slots_15_request = slots_15_io_request; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_15_uop_fu_code = slots_15_io_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] _T_557 = issue_slots_15_uop_fu_code & io_fu_types_0; // @[issue-unit-age-ordered.scala 120:54]
  wire  _T_558 = _T_557 != 10'h0; // @[issue-unit-age-ordered.scala 120:72]
  wire  _T_552 = _T_546 | (_T_531 | (_T_516 | (_T_501 | (_T_486 | (_T_471 | (_T_456 | (_T_441 | (_T_426 | (_T_411 | (
    _T_396 | (_T_381 | (_T_366 | (_T_351 | issue_slots_0_grant))))))))))))); // @[issue-unit-age-ordered.scala 128:69]
  wire  issue_slots_15_grant = issue_slots_15_request & _T_558 & ~_T_552; // @[issue-unit-age-ordered.scala 122:56]
  wire [1:0] _T_79 = issue_slots_14_grant + issue_slots_15_grant; // @[Bitwise.scala 47:55]
  wire [2:0] _T_81 = _T_77 + _T_79; // @[Bitwise.scala 47:55]
  wire [3:0] _T_83 = _T_75 + _T_81; // @[Bitwise.scala 47:55]
  wire [4:0] _T_85 = _T_69 + _T_83; // @[Bitwise.scala 47:55]
  wire  vacants_0 = ~issue_slots_0_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_1 = ~issue_slots_1_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_2 = ~issue_slots_2_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_3 = ~issue_slots_3_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_4 = ~issue_slots_4_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_5 = ~issue_slots_5_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_6 = ~issue_slots_6_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_7 = ~issue_slots_7_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_8 = ~issue_slots_8_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_9 = ~issue_slots_9_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_10 = ~issue_slots_10_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_11 = ~issue_slots_11_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_12 = ~issue_slots_12_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_13 = ~issue_slots_13_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_14 = ~issue_slots_14_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_15 = ~issue_slots_15_valid; // @[issue-unit-age-ordered.scala 39:38]
  wire  vacants_16 = ~io_dis_uops_0_valid; // @[issue-unit-age-ordered.scala 39:82]
  wire [2:0] _GEN_5 = vacants_0 ? 3'h1 : 3'h0; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_104 = {_GEN_5[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_6 = ~_GEN_5[1] & vacants_1 ? _T_104 : {{1'd0}, _GEN_5[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_7 = _GEN_5[1:0] == 2'h0 & vacants_1 ? 3'h1 : _GEN_6; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_110 = {_GEN_7[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_8 = ~_GEN_7[1] & vacants_2 ? _T_110 : {{1'd0}, _GEN_7[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_9 = _GEN_7[1:0] == 2'h0 & vacants_2 ? 3'h1 : _GEN_8; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_116 = {_GEN_9[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_10 = ~_GEN_9[1] & vacants_3 ? _T_116 : {{1'd0}, _GEN_9[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_11 = _GEN_9[1:0] == 2'h0 & vacants_3 ? 3'h1 : _GEN_10; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_122 = {_GEN_11[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_12 = ~_GEN_11[1] & vacants_4 ? _T_122 : {{1'd0}, _GEN_11[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_13 = _GEN_11[1:0] == 2'h0 & vacants_4 ? 3'h1 : _GEN_12; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_128 = {_GEN_13[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_14 = ~_GEN_13[1] & vacants_5 ? _T_128 : {{1'd0}, _GEN_13[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_15 = _GEN_13[1:0] == 2'h0 & vacants_5 ? 3'h1 : _GEN_14; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_134 = {_GEN_15[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_16 = ~_GEN_15[1] & vacants_6 ? _T_134 : {{1'd0}, _GEN_15[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_17 = _GEN_15[1:0] == 2'h0 & vacants_6 ? 3'h1 : _GEN_16; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_140 = {_GEN_17[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_18 = ~_GEN_17[1] & vacants_7 ? _T_140 : {{1'd0}, _GEN_17[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_19 = _GEN_17[1:0] == 2'h0 & vacants_7 ? 3'h1 : _GEN_18; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_146 = {_GEN_19[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_20 = ~_GEN_19[1] & vacants_8 ? _T_146 : {{1'd0}, _GEN_19[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_21 = _GEN_19[1:0] == 2'h0 & vacants_8 ? 3'h1 : _GEN_20; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_152 = {_GEN_21[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_22 = ~_GEN_21[1] & vacants_9 ? _T_152 : {{1'd0}, _GEN_21[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_23 = _GEN_21[1:0] == 2'h0 & vacants_9 ? 3'h1 : _GEN_22; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_158 = {_GEN_23[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_24 = ~_GEN_23[1] & vacants_10 ? _T_158 : {{1'd0}, _GEN_23[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_25 = _GEN_23[1:0] == 2'h0 & vacants_10 ? 3'h1 : _GEN_24; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_164 = {_GEN_25[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_26 = ~_GEN_25[1] & vacants_11 ? _T_164 : {{1'd0}, _GEN_25[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_27 = _GEN_25[1:0] == 2'h0 & vacants_11 ? 3'h1 : _GEN_26; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_170 = {_GEN_27[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_28 = ~_GEN_27[1] & vacants_12 ? _T_170 : {{1'd0}, _GEN_27[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_29 = _GEN_27[1:0] == 2'h0 & vacants_12 ? 3'h1 : _GEN_28; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_176 = {_GEN_29[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_30 = ~_GEN_29[1] & vacants_13 ? _T_176 : {{1'd0}, _GEN_29[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_31 = _GEN_29[1:0] == 2'h0 & vacants_13 ? 3'h1 : _GEN_30; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_182 = {_GEN_31[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_32 = ~_GEN_31[1] & vacants_14 ? _T_182 : {{1'd0}, _GEN_31[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_33 = _GEN_31[1:0] == 2'h0 & vacants_14 ? 3'h1 : _GEN_32; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_188 = {_GEN_33[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_34 = ~_GEN_33[1] & vacants_15 ? _T_188 : {{1'd0}, _GEN_33[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_35 = _GEN_33[1:0] == 2'h0 & vacants_15 ? 3'h1 : _GEN_34; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire [2:0] _T_194 = {_GEN_35[1:0], 1'h0}; // @[issue-unit-age-ordered.scala 48:26]
  wire [2:0] _GEN_36 = ~_GEN_35[1] & vacants_16 ? _T_194 : {{1'd0}, _GEN_35[1:0]}; // @[issue-unit-age-ordered.scala 47:44 issue-unit-age-ordered.scala 48:13 issue-unit-age-ordered.scala 44:11]
  wire [2:0] _GEN_37 = _GEN_35[1:0] == 2'h0 & vacants_16 ? 3'h1 : _GEN_36; // @[issue-unit-age-ordered.scala 45:37 issue-unit-age-ordered.scala 46:13]
  wire  _T_195 = ~io_dis_uops_0_bits_exception; // @[issue-unit-age-ordered.scala 62:57]
  wire  _T_196 = io_dis_uops_0_valid & _T_195; // @[issue-unit-age-ordered.scala 61:77]
  wire  _T_197 = ~io_dis_uops_0_bits_is_fence; // @[issue-unit-age-ordered.scala 63:57]
  wire  _T_198 = _T_196 & _T_197; // @[issue-unit-age-ordered.scala 62:80]
  wire  _T_199 = ~io_dis_uops_0_bits_is_fencei; // @[issue-unit-age-ordered.scala 64:57]
  wire  will_be_valid_16 = _T_198 & _T_199; // @[issue-unit-age-ordered.scala 63:79]
  wire  _T_200 = ~io_dis_uops_1_bits_exception; // @[issue-unit-age-ordered.scala 62:57]
  wire  _T_201 = io_dis_uops_1_valid & _T_200; // @[issue-unit-age-ordered.scala 61:77]
  wire  _T_202 = ~io_dis_uops_1_bits_is_fence; // @[issue-unit-age-ordered.scala 63:57]
  wire  _T_203 = _T_201 & _T_202; // @[issue-unit-age-ordered.scala 62:80]
  wire  _T_204 = ~io_dis_uops_1_bits_is_fencei; // @[issue-unit-age-ordered.scala 64:57]
  wire  will_be_valid_17 = _T_203 & _T_204; // @[issue-unit-age-ordered.scala 63:79]
  wire  issue_slots_1_will_be_valid = slots_1_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_38 = _GEN_5[1:0] == 2'h1 & issue_slots_1_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire [1:0] issue_slots_1_out_uop_debug_tsrc = slots_1_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_1_out_uop_debug_fsrc = slots_1_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_bp_xcpt_if = slots_1_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_bp_debug_if = slots_1_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_xcpt_ma_if = slots_1_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_xcpt_ae_if = slots_1_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_xcpt_pf_if = slots_1_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_fp_single = slots_1_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_fp_val = slots_1_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_frs3_en = slots_1_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_1_out_uop_lrs2_rtype = slots_1_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_1_out_uop_lrs1_rtype = slots_1_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_1_out_uop_dst_rtype = slots_1_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_ldst_val = slots_1_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_1_out_uop_lrs3 = slots_1_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_1_out_uop_lrs2 = slots_1_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_1_out_uop_lrs1 = slots_1_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_1_out_uop_ldst = slots_1_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_ldst_is_rs1 = slots_1_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_flush_on_commit = slots_1_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_unique = slots_1_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_sys_pc2epc = slots_1_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_uses_stq = slots_1_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_uses_ldq = slots_1_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_amo = slots_1_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_fencei = slots_1_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_fence = slots_1_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_mem_signed = slots_1_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_1_out_uop_mem_size = slots_1_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_1_out_uop_mem_cmd = slots_1_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_bypassable = slots_1_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_1_out_uop_exc_cause = slots_1_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_exception = slots_1_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_1_out_uop_stale_pdst = slots_1_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_ppred_busy = slots_1_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_prs3_busy = slots_1_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_prs2_busy = slots_1_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_prs1_busy = slots_1_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_1_out_uop_ppred = slots_1_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_1_out_uop_prs3 = slots_1_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_1_out_uop_prs2 = slots_1_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_1_out_uop_prs1 = slots_1_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_1_out_uop_pdst = slots_1_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_1_out_uop_rxq_idx = slots_1_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_1_out_uop_stq_idx = slots_1_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_1_out_uop_ldq_idx = slots_1_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_1_out_uop_rob_idx = slots_1_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_1_out_uop_csr_addr = slots_1_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_1_out_uop_imm_packed = slots_1_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_taken = slots_1_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_1_out_uop_pc_lob = slots_1_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_edge_inst = slots_1_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_1_out_uop_ftq_idx = slots_1_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_1_out_uop_br_tag = slots_1_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_1_out_uop_br_mask = slots_1_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_sfb = slots_1_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_jal = slots_1_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_jalr = slots_1_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_br = slots_1_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_iw_p2_poisoned = slots_1_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_iw_p1_poisoned = slots_1_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_1_out_uop_iw_state = slots_1_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_1_out_uop_ctrl_op3_sel = slots_1_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_ctrl_is_std = slots_1_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_ctrl_is_sta = slots_1_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_ctrl_is_load = slots_1_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_1_out_uop_ctrl_csr_cmd = slots_1_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_ctrl_fcn_dw = slots_1_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_1_out_uop_ctrl_op_fcn = slots_1_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_1_out_uop_ctrl_imm_sel = slots_1_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_1_out_uop_ctrl_op2_sel = slots_1_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_1_out_uop_ctrl_op1_sel = slots_1_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_1_out_uop_ctrl_br_type = slots_1_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_1_out_uop_fu_code = slots_1_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_1_out_uop_iq_type = slots_1_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_1_out_uop_debug_pc = slots_1_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_rvc = slots_1_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_1_out_uop_debug_inst = slots_1_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_1_out_uop_inst = slots_1_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_1_out_uop_uopc = slots_1_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_1_out_uop_address_num = slots_1_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_1_out_uop_rob_inst_idx = slots_1_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_1_out_uop_self_index = slots_1_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_1_out_uop_split_num = slots_1_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_1_out_uop_op2_sel = slots_1_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_1_out_uop_op1_sel = slots_1_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_1_out_uop_stale_pflag = slots_1_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_pflag_busy = slots_1_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_1_out_uop_pwflag = slots_1_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_1_out_uop_prflag = slots_1_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_wflag = slots_1_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_rflag = slots_1_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_1_out_uop_lrs3_rtype = slots_1_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_1_out_uop_shift = slots_1_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_is_unicore = slots_1_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_switch_off = slots_1_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_out_uop_switch = slots_1_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_will_be_valid = slots_2_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_0_in_uop_valid = _GEN_7[1:0] == 2'h2 ? issue_slots_2_will_be_valid : _GEN_38; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_2_out_uop_debug_tsrc = slots_2_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_2_out_uop_debug_fsrc = slots_2_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_bp_xcpt_if = slots_2_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_bp_debug_if = slots_2_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_xcpt_ma_if = slots_2_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_xcpt_ae_if = slots_2_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_xcpt_pf_if = slots_2_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_fp_single = slots_2_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_fp_val = slots_2_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_frs3_en = slots_2_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_2_out_uop_lrs2_rtype = slots_2_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_2_out_uop_lrs1_rtype = slots_2_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_2_out_uop_dst_rtype = slots_2_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_ldst_val = slots_2_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_2_out_uop_lrs3 = slots_2_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_2_out_uop_lrs2 = slots_2_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_2_out_uop_lrs1 = slots_2_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_2_out_uop_ldst = slots_2_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_ldst_is_rs1 = slots_2_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_flush_on_commit = slots_2_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_unique = slots_2_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_sys_pc2epc = slots_2_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_uses_stq = slots_2_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_uses_ldq = slots_2_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_amo = slots_2_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_fencei = slots_2_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_fence = slots_2_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_mem_signed = slots_2_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_2_out_uop_mem_size = slots_2_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_2_out_uop_mem_cmd = slots_2_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_bypassable = slots_2_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_2_out_uop_exc_cause = slots_2_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_exception = slots_2_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_2_out_uop_stale_pdst = slots_2_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_ppred_busy = slots_2_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_prs3_busy = slots_2_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_prs2_busy = slots_2_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_prs1_busy = slots_2_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_2_out_uop_ppred = slots_2_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_2_out_uop_prs3 = slots_2_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_2_out_uop_prs2 = slots_2_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_2_out_uop_prs1 = slots_2_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_2_out_uop_pdst = slots_2_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_2_out_uop_rxq_idx = slots_2_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_2_out_uop_stq_idx = slots_2_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_2_out_uop_ldq_idx = slots_2_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_2_out_uop_rob_idx = slots_2_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_2_out_uop_csr_addr = slots_2_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_2_out_uop_imm_packed = slots_2_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_taken = slots_2_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_2_out_uop_pc_lob = slots_2_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_edge_inst = slots_2_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_2_out_uop_ftq_idx = slots_2_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_2_out_uop_br_tag = slots_2_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_2_out_uop_br_mask = slots_2_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_sfb = slots_2_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_jal = slots_2_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_jalr = slots_2_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_br = slots_2_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_iw_p2_poisoned = slots_2_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_iw_p1_poisoned = slots_2_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_2_out_uop_iw_state = slots_2_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_2_out_uop_ctrl_op3_sel = slots_2_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_ctrl_is_std = slots_2_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_ctrl_is_sta = slots_2_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_ctrl_is_load = slots_2_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_2_out_uop_ctrl_csr_cmd = slots_2_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_ctrl_fcn_dw = slots_2_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_2_out_uop_ctrl_op_fcn = slots_2_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_2_out_uop_ctrl_imm_sel = slots_2_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_2_out_uop_ctrl_op2_sel = slots_2_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_2_out_uop_ctrl_op1_sel = slots_2_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_2_out_uop_ctrl_br_type = slots_2_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_2_out_uop_fu_code = slots_2_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_2_out_uop_iq_type = slots_2_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_2_out_uop_debug_pc = slots_2_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_rvc = slots_2_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_2_out_uop_debug_inst = slots_2_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_2_out_uop_inst = slots_2_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_2_out_uop_uopc = slots_2_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_2_out_uop_address_num = slots_2_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_2_out_uop_rob_inst_idx = slots_2_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_2_out_uop_self_index = slots_2_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_2_out_uop_split_num = slots_2_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_2_out_uop_op2_sel = slots_2_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_2_out_uop_op1_sel = slots_2_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_2_out_uop_stale_pflag = slots_2_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_pflag_busy = slots_2_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_2_out_uop_pwflag = slots_2_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_2_out_uop_prflag = slots_2_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_wflag = slots_2_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_rflag = slots_2_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_2_out_uop_lrs3_rtype = slots_2_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_2_out_uop_shift = slots_2_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_is_unicore = slots_2_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_switch_off = slots_2_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_out_uop_switch = slots_2_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_234 = _GEN_7[1:0] == 2'h1 & issue_slots_2_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_3_will_be_valid = slots_3_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_in_uop_valid = _GEN_9[1:0] == 2'h2 ? issue_slots_3_will_be_valid : _GEN_234; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_3_out_uop_debug_tsrc = slots_3_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_3_out_uop_debug_fsrc = slots_3_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_bp_xcpt_if = slots_3_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_bp_debug_if = slots_3_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_xcpt_ma_if = slots_3_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_xcpt_ae_if = slots_3_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_xcpt_pf_if = slots_3_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_fp_single = slots_3_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_fp_val = slots_3_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_frs3_en = slots_3_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_3_out_uop_lrs2_rtype = slots_3_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_3_out_uop_lrs1_rtype = slots_3_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_3_out_uop_dst_rtype = slots_3_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_ldst_val = slots_3_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_3_out_uop_lrs3 = slots_3_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_3_out_uop_lrs2 = slots_3_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_3_out_uop_lrs1 = slots_3_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_3_out_uop_ldst = slots_3_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_ldst_is_rs1 = slots_3_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_flush_on_commit = slots_3_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_unique = slots_3_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_sys_pc2epc = slots_3_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_uses_stq = slots_3_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_uses_ldq = slots_3_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_amo = slots_3_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_fencei = slots_3_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_fence = slots_3_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_mem_signed = slots_3_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_3_out_uop_mem_size = slots_3_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_3_out_uop_mem_cmd = slots_3_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_bypassable = slots_3_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_3_out_uop_exc_cause = slots_3_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_exception = slots_3_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_3_out_uop_stale_pdst = slots_3_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_ppred_busy = slots_3_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_prs3_busy = slots_3_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_prs2_busy = slots_3_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_prs1_busy = slots_3_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_3_out_uop_ppred = slots_3_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_3_out_uop_prs3 = slots_3_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_3_out_uop_prs2 = slots_3_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_3_out_uop_prs1 = slots_3_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_3_out_uop_pdst = slots_3_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_3_out_uop_rxq_idx = slots_3_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_3_out_uop_stq_idx = slots_3_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_3_out_uop_ldq_idx = slots_3_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_3_out_uop_rob_idx = slots_3_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_3_out_uop_csr_addr = slots_3_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_3_out_uop_imm_packed = slots_3_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_taken = slots_3_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_3_out_uop_pc_lob = slots_3_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_edge_inst = slots_3_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_3_out_uop_ftq_idx = slots_3_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_3_out_uop_br_tag = slots_3_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_3_out_uop_br_mask = slots_3_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_sfb = slots_3_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_jal = slots_3_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_jalr = slots_3_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_br = slots_3_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_iw_p2_poisoned = slots_3_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_iw_p1_poisoned = slots_3_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_3_out_uop_iw_state = slots_3_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_3_out_uop_ctrl_op3_sel = slots_3_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_ctrl_is_std = slots_3_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_ctrl_is_sta = slots_3_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_ctrl_is_load = slots_3_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_3_out_uop_ctrl_csr_cmd = slots_3_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_ctrl_fcn_dw = slots_3_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_3_out_uop_ctrl_op_fcn = slots_3_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_3_out_uop_ctrl_imm_sel = slots_3_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_3_out_uop_ctrl_op2_sel = slots_3_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_3_out_uop_ctrl_op1_sel = slots_3_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_3_out_uop_ctrl_br_type = slots_3_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_3_out_uop_fu_code = slots_3_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_3_out_uop_iq_type = slots_3_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_3_out_uop_debug_pc = slots_3_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_rvc = slots_3_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_3_out_uop_debug_inst = slots_3_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_3_out_uop_inst = slots_3_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_3_out_uop_uopc = slots_3_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_3_out_uop_address_num = slots_3_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_3_out_uop_rob_inst_idx = slots_3_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_3_out_uop_self_index = slots_3_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_3_out_uop_split_num = slots_3_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_3_out_uop_op2_sel = slots_3_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_3_out_uop_op1_sel = slots_3_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_3_out_uop_stale_pflag = slots_3_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_pflag_busy = slots_3_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_3_out_uop_pwflag = slots_3_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_3_out_uop_prflag = slots_3_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_wflag = slots_3_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_rflag = slots_3_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_3_out_uop_lrs3_rtype = slots_3_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_3_out_uop_shift = slots_3_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_is_unicore = slots_3_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_switch_off = slots_3_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_out_uop_switch = slots_3_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_1_clear = _GEN_5[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_430 = _GEN_9[1:0] == 2'h1 & issue_slots_3_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_4_will_be_valid = slots_4_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_in_uop_valid = _GEN_11[1:0] == 2'h2 ? issue_slots_4_will_be_valid : _GEN_430; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_4_out_uop_debug_tsrc = slots_4_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_4_out_uop_debug_fsrc = slots_4_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_bp_xcpt_if = slots_4_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_bp_debug_if = slots_4_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_xcpt_ma_if = slots_4_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_xcpt_ae_if = slots_4_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_xcpt_pf_if = slots_4_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_fp_single = slots_4_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_fp_val = slots_4_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_frs3_en = slots_4_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_4_out_uop_lrs2_rtype = slots_4_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_4_out_uop_lrs1_rtype = slots_4_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_4_out_uop_dst_rtype = slots_4_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_ldst_val = slots_4_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_4_out_uop_lrs3 = slots_4_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_4_out_uop_lrs2 = slots_4_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_4_out_uop_lrs1 = slots_4_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_4_out_uop_ldst = slots_4_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_ldst_is_rs1 = slots_4_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_flush_on_commit = slots_4_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_unique = slots_4_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_sys_pc2epc = slots_4_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_uses_stq = slots_4_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_uses_ldq = slots_4_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_amo = slots_4_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_fencei = slots_4_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_fence = slots_4_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_mem_signed = slots_4_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_4_out_uop_mem_size = slots_4_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_4_out_uop_mem_cmd = slots_4_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_bypassable = slots_4_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_4_out_uop_exc_cause = slots_4_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_exception = slots_4_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_4_out_uop_stale_pdst = slots_4_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_ppred_busy = slots_4_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_prs3_busy = slots_4_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_prs2_busy = slots_4_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_prs1_busy = slots_4_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_4_out_uop_ppred = slots_4_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_4_out_uop_prs3 = slots_4_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_4_out_uop_prs2 = slots_4_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_4_out_uop_prs1 = slots_4_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_4_out_uop_pdst = slots_4_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_4_out_uop_rxq_idx = slots_4_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_4_out_uop_stq_idx = slots_4_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_4_out_uop_ldq_idx = slots_4_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_4_out_uop_rob_idx = slots_4_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_4_out_uop_csr_addr = slots_4_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_4_out_uop_imm_packed = slots_4_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_taken = slots_4_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_4_out_uop_pc_lob = slots_4_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_edge_inst = slots_4_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_4_out_uop_ftq_idx = slots_4_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_4_out_uop_br_tag = slots_4_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_4_out_uop_br_mask = slots_4_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_sfb = slots_4_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_jal = slots_4_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_jalr = slots_4_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_br = slots_4_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_iw_p2_poisoned = slots_4_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_iw_p1_poisoned = slots_4_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_4_out_uop_iw_state = slots_4_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_4_out_uop_ctrl_op3_sel = slots_4_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_ctrl_is_std = slots_4_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_ctrl_is_sta = slots_4_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_ctrl_is_load = slots_4_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_4_out_uop_ctrl_csr_cmd = slots_4_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_ctrl_fcn_dw = slots_4_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_4_out_uop_ctrl_op_fcn = slots_4_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_4_out_uop_ctrl_imm_sel = slots_4_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_4_out_uop_ctrl_op2_sel = slots_4_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_4_out_uop_ctrl_op1_sel = slots_4_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_4_out_uop_ctrl_br_type = slots_4_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_4_out_uop_fu_code = slots_4_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_4_out_uop_iq_type = slots_4_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_4_out_uop_debug_pc = slots_4_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_rvc = slots_4_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_4_out_uop_debug_inst = slots_4_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_4_out_uop_inst = slots_4_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_4_out_uop_uopc = slots_4_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_4_out_uop_address_num = slots_4_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_4_out_uop_rob_inst_idx = slots_4_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_4_out_uop_self_index = slots_4_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_4_out_uop_split_num = slots_4_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_4_out_uop_op2_sel = slots_4_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_4_out_uop_op1_sel = slots_4_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_4_out_uop_stale_pflag = slots_4_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_pflag_busy = slots_4_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_4_out_uop_pwflag = slots_4_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_4_out_uop_prflag = slots_4_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_wflag = slots_4_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_rflag = slots_4_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_4_out_uop_lrs3_rtype = slots_4_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_4_out_uop_shift = slots_4_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_is_unicore = slots_4_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_switch_off = slots_4_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_out_uop_switch = slots_4_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_2_clear = _GEN_7[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_626 = _GEN_11[1:0] == 2'h1 & issue_slots_4_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_5_will_be_valid = slots_5_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_in_uop_valid = _GEN_13[1:0] == 2'h2 ? issue_slots_5_will_be_valid : _GEN_626; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_5_out_uop_debug_tsrc = slots_5_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_5_out_uop_debug_fsrc = slots_5_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_bp_xcpt_if = slots_5_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_bp_debug_if = slots_5_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_xcpt_ma_if = slots_5_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_xcpt_ae_if = slots_5_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_xcpt_pf_if = slots_5_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_fp_single = slots_5_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_fp_val = slots_5_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_frs3_en = slots_5_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_5_out_uop_lrs2_rtype = slots_5_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_5_out_uop_lrs1_rtype = slots_5_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_5_out_uop_dst_rtype = slots_5_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_ldst_val = slots_5_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_5_out_uop_lrs3 = slots_5_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_5_out_uop_lrs2 = slots_5_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_5_out_uop_lrs1 = slots_5_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_5_out_uop_ldst = slots_5_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_ldst_is_rs1 = slots_5_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_flush_on_commit = slots_5_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_unique = slots_5_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_sys_pc2epc = slots_5_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_uses_stq = slots_5_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_uses_ldq = slots_5_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_amo = slots_5_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_fencei = slots_5_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_fence = slots_5_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_mem_signed = slots_5_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_5_out_uop_mem_size = slots_5_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_5_out_uop_mem_cmd = slots_5_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_bypassable = slots_5_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_5_out_uop_exc_cause = slots_5_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_exception = slots_5_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_5_out_uop_stale_pdst = slots_5_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_ppred_busy = slots_5_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_prs3_busy = slots_5_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_prs2_busy = slots_5_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_prs1_busy = slots_5_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_5_out_uop_ppred = slots_5_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_5_out_uop_prs3 = slots_5_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_5_out_uop_prs2 = slots_5_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_5_out_uop_prs1 = slots_5_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_5_out_uop_pdst = slots_5_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_5_out_uop_rxq_idx = slots_5_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_5_out_uop_stq_idx = slots_5_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_5_out_uop_ldq_idx = slots_5_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_5_out_uop_rob_idx = slots_5_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_5_out_uop_csr_addr = slots_5_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_5_out_uop_imm_packed = slots_5_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_taken = slots_5_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_5_out_uop_pc_lob = slots_5_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_edge_inst = slots_5_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_5_out_uop_ftq_idx = slots_5_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_5_out_uop_br_tag = slots_5_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_5_out_uop_br_mask = slots_5_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_sfb = slots_5_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_jal = slots_5_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_jalr = slots_5_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_br = slots_5_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_iw_p2_poisoned = slots_5_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_iw_p1_poisoned = slots_5_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_5_out_uop_iw_state = slots_5_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_5_out_uop_ctrl_op3_sel = slots_5_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_ctrl_is_std = slots_5_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_ctrl_is_sta = slots_5_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_ctrl_is_load = slots_5_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_5_out_uop_ctrl_csr_cmd = slots_5_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_ctrl_fcn_dw = slots_5_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_5_out_uop_ctrl_op_fcn = slots_5_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_5_out_uop_ctrl_imm_sel = slots_5_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_5_out_uop_ctrl_op2_sel = slots_5_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_5_out_uop_ctrl_op1_sel = slots_5_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_5_out_uop_ctrl_br_type = slots_5_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_5_out_uop_fu_code = slots_5_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_5_out_uop_iq_type = slots_5_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_5_out_uop_debug_pc = slots_5_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_rvc = slots_5_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_5_out_uop_debug_inst = slots_5_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_5_out_uop_inst = slots_5_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_5_out_uop_uopc = slots_5_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_5_out_uop_address_num = slots_5_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_5_out_uop_rob_inst_idx = slots_5_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_5_out_uop_self_index = slots_5_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_5_out_uop_split_num = slots_5_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_5_out_uop_op2_sel = slots_5_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_5_out_uop_op1_sel = slots_5_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_5_out_uop_stale_pflag = slots_5_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_pflag_busy = slots_5_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_5_out_uop_pwflag = slots_5_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_5_out_uop_prflag = slots_5_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_wflag = slots_5_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_rflag = slots_5_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_5_out_uop_lrs3_rtype = slots_5_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_5_out_uop_shift = slots_5_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_is_unicore = slots_5_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_switch_off = slots_5_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_out_uop_switch = slots_5_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_3_clear = _GEN_9[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_822 = _GEN_13[1:0] == 2'h1 & issue_slots_5_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_6_will_be_valid = slots_6_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_in_uop_valid = _GEN_15[1:0] == 2'h2 ? issue_slots_6_will_be_valid : _GEN_822; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_6_out_uop_debug_tsrc = slots_6_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_6_out_uop_debug_fsrc = slots_6_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_bp_xcpt_if = slots_6_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_bp_debug_if = slots_6_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_xcpt_ma_if = slots_6_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_xcpt_ae_if = slots_6_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_xcpt_pf_if = slots_6_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_fp_single = slots_6_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_fp_val = slots_6_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_frs3_en = slots_6_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_6_out_uop_lrs2_rtype = slots_6_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_6_out_uop_lrs1_rtype = slots_6_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_6_out_uop_dst_rtype = slots_6_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_ldst_val = slots_6_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_6_out_uop_lrs3 = slots_6_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_6_out_uop_lrs2 = slots_6_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_6_out_uop_lrs1 = slots_6_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_6_out_uop_ldst = slots_6_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_ldst_is_rs1 = slots_6_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_flush_on_commit = slots_6_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_unique = slots_6_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_sys_pc2epc = slots_6_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_uses_stq = slots_6_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_uses_ldq = slots_6_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_amo = slots_6_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_fencei = slots_6_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_fence = slots_6_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_mem_signed = slots_6_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_6_out_uop_mem_size = slots_6_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_6_out_uop_mem_cmd = slots_6_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_bypassable = slots_6_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_6_out_uop_exc_cause = slots_6_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_exception = slots_6_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_6_out_uop_stale_pdst = slots_6_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_ppred_busy = slots_6_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_prs3_busy = slots_6_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_prs2_busy = slots_6_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_prs1_busy = slots_6_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_6_out_uop_ppred = slots_6_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_6_out_uop_prs3 = slots_6_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_6_out_uop_prs2 = slots_6_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_6_out_uop_prs1 = slots_6_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_6_out_uop_pdst = slots_6_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_6_out_uop_rxq_idx = slots_6_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_6_out_uop_stq_idx = slots_6_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_6_out_uop_ldq_idx = slots_6_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_6_out_uop_rob_idx = slots_6_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_6_out_uop_csr_addr = slots_6_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_6_out_uop_imm_packed = slots_6_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_taken = slots_6_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_6_out_uop_pc_lob = slots_6_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_edge_inst = slots_6_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_6_out_uop_ftq_idx = slots_6_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_6_out_uop_br_tag = slots_6_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_6_out_uop_br_mask = slots_6_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_sfb = slots_6_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_jal = slots_6_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_jalr = slots_6_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_br = slots_6_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_iw_p2_poisoned = slots_6_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_iw_p1_poisoned = slots_6_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_6_out_uop_iw_state = slots_6_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_6_out_uop_ctrl_op3_sel = slots_6_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_ctrl_is_std = slots_6_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_ctrl_is_sta = slots_6_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_ctrl_is_load = slots_6_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_6_out_uop_ctrl_csr_cmd = slots_6_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_ctrl_fcn_dw = slots_6_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_6_out_uop_ctrl_op_fcn = slots_6_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_6_out_uop_ctrl_imm_sel = slots_6_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_6_out_uop_ctrl_op2_sel = slots_6_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_6_out_uop_ctrl_op1_sel = slots_6_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_6_out_uop_ctrl_br_type = slots_6_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_6_out_uop_fu_code = slots_6_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_6_out_uop_iq_type = slots_6_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_6_out_uop_debug_pc = slots_6_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_rvc = slots_6_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_6_out_uop_debug_inst = slots_6_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_6_out_uop_inst = slots_6_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_6_out_uop_uopc = slots_6_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_6_out_uop_address_num = slots_6_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_6_out_uop_rob_inst_idx = slots_6_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_6_out_uop_self_index = slots_6_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_6_out_uop_split_num = slots_6_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_6_out_uop_op2_sel = slots_6_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_6_out_uop_op1_sel = slots_6_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_6_out_uop_stale_pflag = slots_6_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_pflag_busy = slots_6_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_6_out_uop_pwflag = slots_6_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_6_out_uop_prflag = slots_6_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_wflag = slots_6_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_rflag = slots_6_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_6_out_uop_lrs3_rtype = slots_6_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_6_out_uop_shift = slots_6_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_is_unicore = slots_6_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_switch_off = slots_6_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_out_uop_switch = slots_6_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_4_clear = _GEN_11[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_1018 = _GEN_15[1:0] == 2'h1 & issue_slots_6_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_7_will_be_valid = slots_7_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_in_uop_valid = _GEN_17[1:0] == 2'h2 ? issue_slots_7_will_be_valid : _GEN_1018; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_7_out_uop_debug_tsrc = slots_7_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_7_out_uop_debug_fsrc = slots_7_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_bp_xcpt_if = slots_7_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_bp_debug_if = slots_7_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_xcpt_ma_if = slots_7_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_xcpt_ae_if = slots_7_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_xcpt_pf_if = slots_7_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_fp_single = slots_7_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_fp_val = slots_7_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_frs3_en = slots_7_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_7_out_uop_lrs2_rtype = slots_7_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_7_out_uop_lrs1_rtype = slots_7_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_7_out_uop_dst_rtype = slots_7_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_ldst_val = slots_7_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_7_out_uop_lrs3 = slots_7_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_7_out_uop_lrs2 = slots_7_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_7_out_uop_lrs1 = slots_7_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_7_out_uop_ldst = slots_7_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_ldst_is_rs1 = slots_7_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_flush_on_commit = slots_7_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_unique = slots_7_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_sys_pc2epc = slots_7_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_uses_stq = slots_7_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_uses_ldq = slots_7_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_amo = slots_7_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_fencei = slots_7_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_fence = slots_7_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_mem_signed = slots_7_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_7_out_uop_mem_size = slots_7_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_7_out_uop_mem_cmd = slots_7_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_bypassable = slots_7_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_7_out_uop_exc_cause = slots_7_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_exception = slots_7_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_7_out_uop_stale_pdst = slots_7_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_ppred_busy = slots_7_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_prs3_busy = slots_7_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_prs2_busy = slots_7_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_prs1_busy = slots_7_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_7_out_uop_ppred = slots_7_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_7_out_uop_prs3 = slots_7_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_7_out_uop_prs2 = slots_7_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_7_out_uop_prs1 = slots_7_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_7_out_uop_pdst = slots_7_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_7_out_uop_rxq_idx = slots_7_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_7_out_uop_stq_idx = slots_7_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_7_out_uop_ldq_idx = slots_7_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_7_out_uop_rob_idx = slots_7_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_7_out_uop_csr_addr = slots_7_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_7_out_uop_imm_packed = slots_7_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_taken = slots_7_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_7_out_uop_pc_lob = slots_7_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_edge_inst = slots_7_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_7_out_uop_ftq_idx = slots_7_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_7_out_uop_br_tag = slots_7_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_7_out_uop_br_mask = slots_7_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_sfb = slots_7_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_jal = slots_7_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_jalr = slots_7_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_br = slots_7_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_iw_p2_poisoned = slots_7_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_iw_p1_poisoned = slots_7_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_7_out_uop_iw_state = slots_7_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_7_out_uop_ctrl_op3_sel = slots_7_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_ctrl_is_std = slots_7_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_ctrl_is_sta = slots_7_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_ctrl_is_load = slots_7_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_7_out_uop_ctrl_csr_cmd = slots_7_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_ctrl_fcn_dw = slots_7_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_7_out_uop_ctrl_op_fcn = slots_7_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_7_out_uop_ctrl_imm_sel = slots_7_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_7_out_uop_ctrl_op2_sel = slots_7_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_7_out_uop_ctrl_op1_sel = slots_7_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_7_out_uop_ctrl_br_type = slots_7_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_7_out_uop_fu_code = slots_7_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_7_out_uop_iq_type = slots_7_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_7_out_uop_debug_pc = slots_7_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_rvc = slots_7_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_7_out_uop_debug_inst = slots_7_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_7_out_uop_inst = slots_7_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_7_out_uop_uopc = slots_7_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_7_out_uop_address_num = slots_7_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_7_out_uop_rob_inst_idx = slots_7_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_7_out_uop_self_index = slots_7_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_7_out_uop_split_num = slots_7_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_7_out_uop_op2_sel = slots_7_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_7_out_uop_op1_sel = slots_7_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_7_out_uop_stale_pflag = slots_7_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_pflag_busy = slots_7_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_7_out_uop_pwflag = slots_7_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_7_out_uop_prflag = slots_7_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_wflag = slots_7_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_rflag = slots_7_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_7_out_uop_lrs3_rtype = slots_7_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_7_out_uop_shift = slots_7_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_is_unicore = slots_7_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_switch_off = slots_7_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_out_uop_switch = slots_7_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_5_clear = _GEN_13[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_1214 = _GEN_17[1:0] == 2'h1 & issue_slots_7_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_8_will_be_valid = slots_8_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_in_uop_valid = _GEN_19[1:0] == 2'h2 ? issue_slots_8_will_be_valid : _GEN_1214; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_8_out_uop_debug_tsrc = slots_8_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_8_out_uop_debug_fsrc = slots_8_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_bp_xcpt_if = slots_8_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_bp_debug_if = slots_8_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_xcpt_ma_if = slots_8_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_xcpt_ae_if = slots_8_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_xcpt_pf_if = slots_8_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_fp_single = slots_8_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_fp_val = slots_8_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_frs3_en = slots_8_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_8_out_uop_lrs2_rtype = slots_8_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_8_out_uop_lrs1_rtype = slots_8_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_8_out_uop_dst_rtype = slots_8_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_ldst_val = slots_8_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_8_out_uop_lrs3 = slots_8_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_8_out_uop_lrs2 = slots_8_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_8_out_uop_lrs1 = slots_8_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_8_out_uop_ldst = slots_8_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_ldst_is_rs1 = slots_8_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_flush_on_commit = slots_8_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_unique = slots_8_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_sys_pc2epc = slots_8_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_uses_stq = slots_8_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_uses_ldq = slots_8_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_amo = slots_8_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_fencei = slots_8_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_fence = slots_8_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_mem_signed = slots_8_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_8_out_uop_mem_size = slots_8_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_8_out_uop_mem_cmd = slots_8_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_bypassable = slots_8_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_8_out_uop_exc_cause = slots_8_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_exception = slots_8_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_8_out_uop_stale_pdst = slots_8_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_ppred_busy = slots_8_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_prs3_busy = slots_8_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_prs2_busy = slots_8_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_prs1_busy = slots_8_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_8_out_uop_ppred = slots_8_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_8_out_uop_prs3 = slots_8_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_8_out_uop_prs2 = slots_8_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_8_out_uop_prs1 = slots_8_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_8_out_uop_pdst = slots_8_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_8_out_uop_rxq_idx = slots_8_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_8_out_uop_stq_idx = slots_8_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_8_out_uop_ldq_idx = slots_8_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_8_out_uop_rob_idx = slots_8_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_8_out_uop_csr_addr = slots_8_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_8_out_uop_imm_packed = slots_8_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_taken = slots_8_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_8_out_uop_pc_lob = slots_8_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_edge_inst = slots_8_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_8_out_uop_ftq_idx = slots_8_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_8_out_uop_br_tag = slots_8_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_8_out_uop_br_mask = slots_8_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_sfb = slots_8_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_jal = slots_8_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_jalr = slots_8_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_br = slots_8_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_iw_p2_poisoned = slots_8_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_iw_p1_poisoned = slots_8_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_8_out_uop_iw_state = slots_8_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_8_out_uop_ctrl_op3_sel = slots_8_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_ctrl_is_std = slots_8_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_ctrl_is_sta = slots_8_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_ctrl_is_load = slots_8_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_8_out_uop_ctrl_csr_cmd = slots_8_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_ctrl_fcn_dw = slots_8_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_8_out_uop_ctrl_op_fcn = slots_8_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_8_out_uop_ctrl_imm_sel = slots_8_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_8_out_uop_ctrl_op2_sel = slots_8_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_8_out_uop_ctrl_op1_sel = slots_8_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_8_out_uop_ctrl_br_type = slots_8_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_8_out_uop_fu_code = slots_8_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_8_out_uop_iq_type = slots_8_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_8_out_uop_debug_pc = slots_8_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_rvc = slots_8_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_8_out_uop_debug_inst = slots_8_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_8_out_uop_inst = slots_8_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_8_out_uop_uopc = slots_8_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_8_out_uop_address_num = slots_8_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_8_out_uop_rob_inst_idx = slots_8_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_8_out_uop_self_index = slots_8_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_8_out_uop_split_num = slots_8_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_8_out_uop_op2_sel = slots_8_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_8_out_uop_op1_sel = slots_8_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_8_out_uop_stale_pflag = slots_8_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_pflag_busy = slots_8_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_8_out_uop_pwflag = slots_8_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_8_out_uop_prflag = slots_8_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_wflag = slots_8_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_rflag = slots_8_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_8_out_uop_lrs3_rtype = slots_8_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_8_out_uop_shift = slots_8_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_is_unicore = slots_8_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_switch_off = slots_8_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_out_uop_switch = slots_8_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_6_clear = _GEN_15[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_1410 = _GEN_19[1:0] == 2'h1 & issue_slots_8_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_9_will_be_valid = slots_9_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_in_uop_valid = _GEN_21[1:0] == 2'h2 ? issue_slots_9_will_be_valid : _GEN_1410; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_9_out_uop_debug_tsrc = slots_9_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_9_out_uop_debug_fsrc = slots_9_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_bp_xcpt_if = slots_9_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_bp_debug_if = slots_9_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_xcpt_ma_if = slots_9_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_xcpt_ae_if = slots_9_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_xcpt_pf_if = slots_9_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_fp_single = slots_9_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_fp_val = slots_9_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_frs3_en = slots_9_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_9_out_uop_lrs2_rtype = slots_9_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_9_out_uop_lrs1_rtype = slots_9_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_9_out_uop_dst_rtype = slots_9_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_ldst_val = slots_9_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_9_out_uop_lrs3 = slots_9_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_9_out_uop_lrs2 = slots_9_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_9_out_uop_lrs1 = slots_9_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_9_out_uop_ldst = slots_9_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_ldst_is_rs1 = slots_9_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_flush_on_commit = slots_9_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_unique = slots_9_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_sys_pc2epc = slots_9_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_uses_stq = slots_9_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_uses_ldq = slots_9_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_amo = slots_9_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_fencei = slots_9_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_fence = slots_9_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_mem_signed = slots_9_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_9_out_uop_mem_size = slots_9_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_9_out_uop_mem_cmd = slots_9_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_bypassable = slots_9_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_9_out_uop_exc_cause = slots_9_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_exception = slots_9_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_9_out_uop_stale_pdst = slots_9_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_ppred_busy = slots_9_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_prs3_busy = slots_9_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_prs2_busy = slots_9_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_prs1_busy = slots_9_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_9_out_uop_ppred = slots_9_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_9_out_uop_prs3 = slots_9_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_9_out_uop_prs2 = slots_9_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_9_out_uop_prs1 = slots_9_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_9_out_uop_pdst = slots_9_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_9_out_uop_rxq_idx = slots_9_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_9_out_uop_stq_idx = slots_9_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_9_out_uop_ldq_idx = slots_9_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_9_out_uop_rob_idx = slots_9_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_9_out_uop_csr_addr = slots_9_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_9_out_uop_imm_packed = slots_9_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_taken = slots_9_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_9_out_uop_pc_lob = slots_9_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_edge_inst = slots_9_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_9_out_uop_ftq_idx = slots_9_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_9_out_uop_br_tag = slots_9_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_9_out_uop_br_mask = slots_9_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_sfb = slots_9_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_jal = slots_9_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_jalr = slots_9_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_br = slots_9_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_iw_p2_poisoned = slots_9_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_iw_p1_poisoned = slots_9_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_9_out_uop_iw_state = slots_9_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_9_out_uop_ctrl_op3_sel = slots_9_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_ctrl_is_std = slots_9_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_ctrl_is_sta = slots_9_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_ctrl_is_load = slots_9_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_9_out_uop_ctrl_csr_cmd = slots_9_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_ctrl_fcn_dw = slots_9_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_9_out_uop_ctrl_op_fcn = slots_9_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_9_out_uop_ctrl_imm_sel = slots_9_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_9_out_uop_ctrl_op2_sel = slots_9_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_9_out_uop_ctrl_op1_sel = slots_9_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_9_out_uop_ctrl_br_type = slots_9_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_9_out_uop_fu_code = slots_9_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_9_out_uop_iq_type = slots_9_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_9_out_uop_debug_pc = slots_9_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_rvc = slots_9_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_9_out_uop_debug_inst = slots_9_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_9_out_uop_inst = slots_9_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_9_out_uop_uopc = slots_9_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_9_out_uop_address_num = slots_9_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_9_out_uop_rob_inst_idx = slots_9_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_9_out_uop_self_index = slots_9_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_9_out_uop_split_num = slots_9_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_9_out_uop_op2_sel = slots_9_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_9_out_uop_op1_sel = slots_9_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_9_out_uop_stale_pflag = slots_9_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_pflag_busy = slots_9_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_9_out_uop_pwflag = slots_9_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_9_out_uop_prflag = slots_9_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_wflag = slots_9_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_rflag = slots_9_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_9_out_uop_lrs3_rtype = slots_9_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_9_out_uop_shift = slots_9_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_is_unicore = slots_9_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_switch_off = slots_9_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_out_uop_switch = slots_9_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_7_clear = _GEN_17[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_1606 = _GEN_21[1:0] == 2'h1 & issue_slots_9_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_10_will_be_valid = slots_10_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_in_uop_valid = _GEN_23[1:0] == 2'h2 ? issue_slots_10_will_be_valid : _GEN_1606; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_10_out_uop_debug_tsrc = slots_10_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_10_out_uop_debug_fsrc = slots_10_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_bp_xcpt_if = slots_10_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_bp_debug_if = slots_10_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_xcpt_ma_if = slots_10_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_xcpt_ae_if = slots_10_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_xcpt_pf_if = slots_10_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_fp_single = slots_10_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_fp_val = slots_10_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_frs3_en = slots_10_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_10_out_uop_lrs2_rtype = slots_10_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_10_out_uop_lrs1_rtype = slots_10_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_10_out_uop_dst_rtype = slots_10_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_ldst_val = slots_10_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_10_out_uop_lrs3 = slots_10_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_10_out_uop_lrs2 = slots_10_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_10_out_uop_lrs1 = slots_10_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_10_out_uop_ldst = slots_10_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_ldst_is_rs1 = slots_10_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_flush_on_commit = slots_10_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_unique = slots_10_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_sys_pc2epc = slots_10_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_uses_stq = slots_10_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_uses_ldq = slots_10_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_amo = slots_10_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_fencei = slots_10_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_fence = slots_10_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_mem_signed = slots_10_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_10_out_uop_mem_size = slots_10_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_10_out_uop_mem_cmd = slots_10_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_bypassable = slots_10_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_10_out_uop_exc_cause = slots_10_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_exception = slots_10_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_10_out_uop_stale_pdst = slots_10_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_ppred_busy = slots_10_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_prs3_busy = slots_10_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_prs2_busy = slots_10_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_prs1_busy = slots_10_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_10_out_uop_ppred = slots_10_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_10_out_uop_prs3 = slots_10_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_10_out_uop_prs2 = slots_10_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_10_out_uop_prs1 = slots_10_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_10_out_uop_pdst = slots_10_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_10_out_uop_rxq_idx = slots_10_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_10_out_uop_stq_idx = slots_10_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_10_out_uop_ldq_idx = slots_10_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_10_out_uop_rob_idx = slots_10_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_10_out_uop_csr_addr = slots_10_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_10_out_uop_imm_packed = slots_10_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_taken = slots_10_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_10_out_uop_pc_lob = slots_10_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_edge_inst = slots_10_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_10_out_uop_ftq_idx = slots_10_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_10_out_uop_br_tag = slots_10_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_10_out_uop_br_mask = slots_10_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_sfb = slots_10_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_jal = slots_10_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_jalr = slots_10_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_br = slots_10_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_iw_p2_poisoned = slots_10_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_iw_p1_poisoned = slots_10_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_10_out_uop_iw_state = slots_10_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_10_out_uop_ctrl_op3_sel = slots_10_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_ctrl_is_std = slots_10_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_ctrl_is_sta = slots_10_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_ctrl_is_load = slots_10_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_10_out_uop_ctrl_csr_cmd = slots_10_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_ctrl_fcn_dw = slots_10_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_10_out_uop_ctrl_op_fcn = slots_10_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_10_out_uop_ctrl_imm_sel = slots_10_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_10_out_uop_ctrl_op2_sel = slots_10_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_10_out_uop_ctrl_op1_sel = slots_10_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_10_out_uop_ctrl_br_type = slots_10_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_10_out_uop_fu_code = slots_10_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_10_out_uop_iq_type = slots_10_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_10_out_uop_debug_pc = slots_10_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_rvc = slots_10_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_10_out_uop_debug_inst = slots_10_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_10_out_uop_inst = slots_10_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_10_out_uop_uopc = slots_10_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_10_out_uop_address_num = slots_10_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_10_out_uop_rob_inst_idx = slots_10_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_10_out_uop_self_index = slots_10_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_10_out_uop_split_num = slots_10_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_10_out_uop_op2_sel = slots_10_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_10_out_uop_op1_sel = slots_10_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_10_out_uop_stale_pflag = slots_10_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_pflag_busy = slots_10_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_10_out_uop_pwflag = slots_10_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_10_out_uop_prflag = slots_10_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_wflag = slots_10_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_rflag = slots_10_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_10_out_uop_lrs3_rtype = slots_10_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_10_out_uop_shift = slots_10_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_is_unicore = slots_10_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_switch_off = slots_10_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_out_uop_switch = slots_10_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_8_clear = _GEN_19[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_1802 = _GEN_23[1:0] == 2'h1 & issue_slots_10_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_11_will_be_valid = slots_11_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_in_uop_valid = _GEN_25[1:0] == 2'h2 ? issue_slots_11_will_be_valid : _GEN_1802; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_11_out_uop_debug_tsrc = slots_11_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_11_out_uop_debug_fsrc = slots_11_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_bp_xcpt_if = slots_11_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_bp_debug_if = slots_11_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_xcpt_ma_if = slots_11_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_xcpt_ae_if = slots_11_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_xcpt_pf_if = slots_11_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_fp_single = slots_11_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_fp_val = slots_11_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_frs3_en = slots_11_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_11_out_uop_lrs2_rtype = slots_11_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_11_out_uop_lrs1_rtype = slots_11_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_11_out_uop_dst_rtype = slots_11_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_ldst_val = slots_11_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_11_out_uop_lrs3 = slots_11_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_11_out_uop_lrs2 = slots_11_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_11_out_uop_lrs1 = slots_11_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_11_out_uop_ldst = slots_11_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_ldst_is_rs1 = slots_11_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_flush_on_commit = slots_11_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_unique = slots_11_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_sys_pc2epc = slots_11_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_uses_stq = slots_11_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_uses_ldq = slots_11_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_amo = slots_11_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_fencei = slots_11_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_fence = slots_11_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_mem_signed = slots_11_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_11_out_uop_mem_size = slots_11_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_11_out_uop_mem_cmd = slots_11_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_bypassable = slots_11_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_11_out_uop_exc_cause = slots_11_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_exception = slots_11_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_11_out_uop_stale_pdst = slots_11_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_ppred_busy = slots_11_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_prs3_busy = slots_11_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_prs2_busy = slots_11_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_prs1_busy = slots_11_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_11_out_uop_ppred = slots_11_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_11_out_uop_prs3 = slots_11_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_11_out_uop_prs2 = slots_11_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_11_out_uop_prs1 = slots_11_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_11_out_uop_pdst = slots_11_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_11_out_uop_rxq_idx = slots_11_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_11_out_uop_stq_idx = slots_11_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_11_out_uop_ldq_idx = slots_11_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_11_out_uop_rob_idx = slots_11_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_11_out_uop_csr_addr = slots_11_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_11_out_uop_imm_packed = slots_11_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_taken = slots_11_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_11_out_uop_pc_lob = slots_11_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_edge_inst = slots_11_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_11_out_uop_ftq_idx = slots_11_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_11_out_uop_br_tag = slots_11_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_11_out_uop_br_mask = slots_11_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_sfb = slots_11_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_jal = slots_11_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_jalr = slots_11_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_br = slots_11_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_iw_p2_poisoned = slots_11_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_iw_p1_poisoned = slots_11_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_11_out_uop_iw_state = slots_11_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_11_out_uop_ctrl_op3_sel = slots_11_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_ctrl_is_std = slots_11_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_ctrl_is_sta = slots_11_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_ctrl_is_load = slots_11_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_11_out_uop_ctrl_csr_cmd = slots_11_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_ctrl_fcn_dw = slots_11_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_11_out_uop_ctrl_op_fcn = slots_11_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_11_out_uop_ctrl_imm_sel = slots_11_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_11_out_uop_ctrl_op2_sel = slots_11_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_11_out_uop_ctrl_op1_sel = slots_11_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_11_out_uop_ctrl_br_type = slots_11_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_11_out_uop_fu_code = slots_11_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_11_out_uop_iq_type = slots_11_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_11_out_uop_debug_pc = slots_11_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_rvc = slots_11_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_11_out_uop_debug_inst = slots_11_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_11_out_uop_inst = slots_11_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_11_out_uop_uopc = slots_11_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_11_out_uop_address_num = slots_11_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_11_out_uop_rob_inst_idx = slots_11_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_11_out_uop_self_index = slots_11_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_11_out_uop_split_num = slots_11_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_11_out_uop_op2_sel = slots_11_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_11_out_uop_op1_sel = slots_11_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_11_out_uop_stale_pflag = slots_11_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_pflag_busy = slots_11_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_11_out_uop_pwflag = slots_11_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_11_out_uop_prflag = slots_11_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_wflag = slots_11_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_rflag = slots_11_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_11_out_uop_lrs3_rtype = slots_11_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_11_out_uop_shift = slots_11_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_is_unicore = slots_11_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_switch_off = slots_11_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_out_uop_switch = slots_11_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_9_clear = _GEN_21[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_1998 = _GEN_25[1:0] == 2'h1 & issue_slots_11_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_12_will_be_valid = slots_12_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_in_uop_valid = _GEN_27[1:0] == 2'h2 ? issue_slots_12_will_be_valid : _GEN_1998; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_12_out_uop_debug_tsrc = slots_12_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_12_out_uop_debug_fsrc = slots_12_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_bp_xcpt_if = slots_12_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_bp_debug_if = slots_12_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_xcpt_ma_if = slots_12_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_xcpt_ae_if = slots_12_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_xcpt_pf_if = slots_12_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_fp_single = slots_12_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_fp_val = slots_12_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_frs3_en = slots_12_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_12_out_uop_lrs2_rtype = slots_12_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_12_out_uop_lrs1_rtype = slots_12_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_12_out_uop_dst_rtype = slots_12_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_ldst_val = slots_12_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_12_out_uop_lrs3 = slots_12_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_12_out_uop_lrs2 = slots_12_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_12_out_uop_lrs1 = slots_12_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_12_out_uop_ldst = slots_12_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_ldst_is_rs1 = slots_12_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_flush_on_commit = slots_12_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_unique = slots_12_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_sys_pc2epc = slots_12_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_uses_stq = slots_12_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_uses_ldq = slots_12_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_amo = slots_12_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_fencei = slots_12_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_fence = slots_12_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_mem_signed = slots_12_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_12_out_uop_mem_size = slots_12_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_12_out_uop_mem_cmd = slots_12_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_bypassable = slots_12_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_12_out_uop_exc_cause = slots_12_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_exception = slots_12_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_12_out_uop_stale_pdst = slots_12_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_ppred_busy = slots_12_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_prs3_busy = slots_12_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_prs2_busy = slots_12_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_prs1_busy = slots_12_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_12_out_uop_ppred = slots_12_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_12_out_uop_prs3 = slots_12_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_12_out_uop_prs2 = slots_12_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_12_out_uop_prs1 = slots_12_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_12_out_uop_pdst = slots_12_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_12_out_uop_rxq_idx = slots_12_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_12_out_uop_stq_idx = slots_12_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_12_out_uop_ldq_idx = slots_12_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_12_out_uop_rob_idx = slots_12_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_12_out_uop_csr_addr = slots_12_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_12_out_uop_imm_packed = slots_12_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_taken = slots_12_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_12_out_uop_pc_lob = slots_12_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_edge_inst = slots_12_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_12_out_uop_ftq_idx = slots_12_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_12_out_uop_br_tag = slots_12_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_12_out_uop_br_mask = slots_12_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_sfb = slots_12_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_jal = slots_12_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_jalr = slots_12_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_br = slots_12_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_iw_p2_poisoned = slots_12_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_iw_p1_poisoned = slots_12_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_12_out_uop_iw_state = slots_12_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_12_out_uop_ctrl_op3_sel = slots_12_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_ctrl_is_std = slots_12_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_ctrl_is_sta = slots_12_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_ctrl_is_load = slots_12_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_12_out_uop_ctrl_csr_cmd = slots_12_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_ctrl_fcn_dw = slots_12_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_12_out_uop_ctrl_op_fcn = slots_12_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_12_out_uop_ctrl_imm_sel = slots_12_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_12_out_uop_ctrl_op2_sel = slots_12_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_12_out_uop_ctrl_op1_sel = slots_12_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_12_out_uop_ctrl_br_type = slots_12_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_12_out_uop_fu_code = slots_12_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_12_out_uop_iq_type = slots_12_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_12_out_uop_debug_pc = slots_12_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_rvc = slots_12_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_12_out_uop_debug_inst = slots_12_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_12_out_uop_inst = slots_12_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_12_out_uop_uopc = slots_12_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_12_out_uop_address_num = slots_12_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_12_out_uop_rob_inst_idx = slots_12_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_12_out_uop_self_index = slots_12_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_12_out_uop_split_num = slots_12_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_12_out_uop_op2_sel = slots_12_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_12_out_uop_op1_sel = slots_12_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_12_out_uop_stale_pflag = slots_12_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_pflag_busy = slots_12_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_12_out_uop_pwflag = slots_12_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_12_out_uop_prflag = slots_12_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_wflag = slots_12_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_rflag = slots_12_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_12_out_uop_lrs3_rtype = slots_12_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_12_out_uop_shift = slots_12_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_is_unicore = slots_12_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_switch_off = slots_12_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_out_uop_switch = slots_12_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_10_clear = _GEN_23[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_2194 = _GEN_27[1:0] == 2'h1 & issue_slots_12_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_13_will_be_valid = slots_13_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_in_uop_valid = _GEN_29[1:0] == 2'h2 ? issue_slots_13_will_be_valid : _GEN_2194; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_13_out_uop_debug_tsrc = slots_13_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_13_out_uop_debug_fsrc = slots_13_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_bp_xcpt_if = slots_13_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_bp_debug_if = slots_13_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_xcpt_ma_if = slots_13_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_xcpt_ae_if = slots_13_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_xcpt_pf_if = slots_13_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_fp_single = slots_13_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_fp_val = slots_13_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_frs3_en = slots_13_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_13_out_uop_lrs2_rtype = slots_13_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_13_out_uop_lrs1_rtype = slots_13_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_13_out_uop_dst_rtype = slots_13_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_ldst_val = slots_13_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_13_out_uop_lrs3 = slots_13_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_13_out_uop_lrs2 = slots_13_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_13_out_uop_lrs1 = slots_13_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_13_out_uop_ldst = slots_13_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_ldst_is_rs1 = slots_13_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_flush_on_commit = slots_13_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_unique = slots_13_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_sys_pc2epc = slots_13_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_uses_stq = slots_13_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_uses_ldq = slots_13_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_amo = slots_13_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_fencei = slots_13_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_fence = slots_13_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_mem_signed = slots_13_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_13_out_uop_mem_size = slots_13_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_13_out_uop_mem_cmd = slots_13_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_bypassable = slots_13_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_13_out_uop_exc_cause = slots_13_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_exception = slots_13_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_13_out_uop_stale_pdst = slots_13_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_ppred_busy = slots_13_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_prs3_busy = slots_13_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_prs2_busy = slots_13_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_prs1_busy = slots_13_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_13_out_uop_ppred = slots_13_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_13_out_uop_prs3 = slots_13_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_13_out_uop_prs2 = slots_13_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_13_out_uop_prs1 = slots_13_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_13_out_uop_pdst = slots_13_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_13_out_uop_rxq_idx = slots_13_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_13_out_uop_stq_idx = slots_13_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_13_out_uop_ldq_idx = slots_13_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_13_out_uop_rob_idx = slots_13_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_13_out_uop_csr_addr = slots_13_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_13_out_uop_imm_packed = slots_13_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_taken = slots_13_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_13_out_uop_pc_lob = slots_13_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_edge_inst = slots_13_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_13_out_uop_ftq_idx = slots_13_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_13_out_uop_br_tag = slots_13_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_13_out_uop_br_mask = slots_13_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_sfb = slots_13_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_jal = slots_13_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_jalr = slots_13_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_br = slots_13_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_iw_p2_poisoned = slots_13_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_iw_p1_poisoned = slots_13_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_13_out_uop_iw_state = slots_13_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_13_out_uop_ctrl_op3_sel = slots_13_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_ctrl_is_std = slots_13_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_ctrl_is_sta = slots_13_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_ctrl_is_load = slots_13_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_13_out_uop_ctrl_csr_cmd = slots_13_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_ctrl_fcn_dw = slots_13_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_13_out_uop_ctrl_op_fcn = slots_13_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_13_out_uop_ctrl_imm_sel = slots_13_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_13_out_uop_ctrl_op2_sel = slots_13_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_13_out_uop_ctrl_op1_sel = slots_13_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_13_out_uop_ctrl_br_type = slots_13_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_13_out_uop_fu_code = slots_13_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_13_out_uop_iq_type = slots_13_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_13_out_uop_debug_pc = slots_13_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_rvc = slots_13_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_13_out_uop_debug_inst = slots_13_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_13_out_uop_inst = slots_13_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_13_out_uop_uopc = slots_13_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_13_out_uop_address_num = slots_13_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_13_out_uop_rob_inst_idx = slots_13_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_13_out_uop_self_index = slots_13_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_13_out_uop_split_num = slots_13_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_13_out_uop_op2_sel = slots_13_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_13_out_uop_op1_sel = slots_13_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_13_out_uop_stale_pflag = slots_13_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_pflag_busy = slots_13_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_13_out_uop_pwflag = slots_13_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_13_out_uop_prflag = slots_13_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_wflag = slots_13_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_rflag = slots_13_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_13_out_uop_lrs3_rtype = slots_13_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_13_out_uop_shift = slots_13_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_is_unicore = slots_13_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_switch_off = slots_13_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_out_uop_switch = slots_13_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_11_clear = _GEN_25[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_2390 = _GEN_29[1:0] == 2'h1 & issue_slots_13_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_14_will_be_valid = slots_14_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_in_uop_valid = _GEN_31[1:0] == 2'h2 ? issue_slots_14_will_be_valid : _GEN_2390; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_14_out_uop_debug_tsrc = slots_14_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_14_out_uop_debug_fsrc = slots_14_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_bp_xcpt_if = slots_14_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_bp_debug_if = slots_14_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_xcpt_ma_if = slots_14_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_xcpt_ae_if = slots_14_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_xcpt_pf_if = slots_14_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_fp_single = slots_14_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_fp_val = slots_14_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_frs3_en = slots_14_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_14_out_uop_lrs2_rtype = slots_14_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_14_out_uop_lrs1_rtype = slots_14_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_14_out_uop_dst_rtype = slots_14_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_ldst_val = slots_14_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_14_out_uop_lrs3 = slots_14_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_14_out_uop_lrs2 = slots_14_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_14_out_uop_lrs1 = slots_14_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_14_out_uop_ldst = slots_14_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_ldst_is_rs1 = slots_14_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_flush_on_commit = slots_14_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_unique = slots_14_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_sys_pc2epc = slots_14_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_uses_stq = slots_14_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_uses_ldq = slots_14_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_amo = slots_14_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_fencei = slots_14_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_fence = slots_14_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_mem_signed = slots_14_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_14_out_uop_mem_size = slots_14_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_14_out_uop_mem_cmd = slots_14_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_bypassable = slots_14_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_14_out_uop_exc_cause = slots_14_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_exception = slots_14_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_14_out_uop_stale_pdst = slots_14_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_ppred_busy = slots_14_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_prs3_busy = slots_14_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_prs2_busy = slots_14_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_prs1_busy = slots_14_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_14_out_uop_ppred = slots_14_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_14_out_uop_prs3 = slots_14_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_14_out_uop_prs2 = slots_14_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_14_out_uop_prs1 = slots_14_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_14_out_uop_pdst = slots_14_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_14_out_uop_rxq_idx = slots_14_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_14_out_uop_stq_idx = slots_14_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_14_out_uop_ldq_idx = slots_14_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_14_out_uop_rob_idx = slots_14_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_14_out_uop_csr_addr = slots_14_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_14_out_uop_imm_packed = slots_14_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_taken = slots_14_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_14_out_uop_pc_lob = slots_14_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_edge_inst = slots_14_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_14_out_uop_ftq_idx = slots_14_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_14_out_uop_br_tag = slots_14_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_14_out_uop_br_mask = slots_14_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_sfb = slots_14_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_jal = slots_14_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_jalr = slots_14_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_br = slots_14_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_iw_p2_poisoned = slots_14_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_iw_p1_poisoned = slots_14_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_14_out_uop_iw_state = slots_14_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_14_out_uop_ctrl_op3_sel = slots_14_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_ctrl_is_std = slots_14_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_ctrl_is_sta = slots_14_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_ctrl_is_load = slots_14_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_14_out_uop_ctrl_csr_cmd = slots_14_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_ctrl_fcn_dw = slots_14_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_14_out_uop_ctrl_op_fcn = slots_14_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_14_out_uop_ctrl_imm_sel = slots_14_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_14_out_uop_ctrl_op2_sel = slots_14_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_14_out_uop_ctrl_op1_sel = slots_14_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_14_out_uop_ctrl_br_type = slots_14_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_14_out_uop_fu_code = slots_14_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_14_out_uop_iq_type = slots_14_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_14_out_uop_debug_pc = slots_14_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_rvc = slots_14_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_14_out_uop_debug_inst = slots_14_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_14_out_uop_inst = slots_14_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_14_out_uop_uopc = slots_14_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_14_out_uop_address_num = slots_14_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_14_out_uop_rob_inst_idx = slots_14_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_14_out_uop_self_index = slots_14_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_14_out_uop_split_num = slots_14_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_14_out_uop_op2_sel = slots_14_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_14_out_uop_op1_sel = slots_14_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_14_out_uop_stale_pflag = slots_14_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_pflag_busy = slots_14_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_14_out_uop_pwflag = slots_14_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_14_out_uop_prflag = slots_14_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_wflag = slots_14_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_rflag = slots_14_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_14_out_uop_lrs3_rtype = slots_14_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_14_out_uop_shift = slots_14_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_is_unicore = slots_14_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_switch_off = slots_14_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_14_out_uop_switch = slots_14_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_12_clear = _GEN_27[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_2586 = _GEN_31[1:0] == 2'h1 & issue_slots_14_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_15_will_be_valid = slots_15_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_in_uop_valid = _GEN_33[1:0] == 2'h2 ? issue_slots_15_will_be_valid : _GEN_2586; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire [1:0] issue_slots_15_out_uop_debug_tsrc = slots_15_io_out_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_out_uop_debug_fsrc = slots_15_io_out_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_bp_xcpt_if = slots_15_io_out_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_bp_debug_if = slots_15_io_out_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_xcpt_ma_if = slots_15_io_out_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_xcpt_ae_if = slots_15_io_out_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_xcpt_pf_if = slots_15_io_out_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_fp_single = slots_15_io_out_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_fp_val = slots_15_io_out_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_frs3_en = slots_15_io_out_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_out_uop_lrs2_rtype = slots_15_io_out_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_out_uop_lrs1_rtype = slots_15_io_out_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_out_uop_dst_rtype = slots_15_io_out_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_ldst_val = slots_15_io_out_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_out_uop_lrs3 = slots_15_io_out_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_out_uop_lrs2 = slots_15_io_out_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_out_uop_lrs1 = slots_15_io_out_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_out_uop_ldst = slots_15_io_out_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_ldst_is_rs1 = slots_15_io_out_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_flush_on_commit = slots_15_io_out_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_unique = slots_15_io_out_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_sys_pc2epc = slots_15_io_out_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_uses_stq = slots_15_io_out_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_uses_ldq = slots_15_io_out_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_amo = slots_15_io_out_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_fencei = slots_15_io_out_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_fence = slots_15_io_out_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_mem_signed = slots_15_io_out_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_out_uop_mem_size = slots_15_io_out_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_15_out_uop_mem_cmd = slots_15_io_out_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_bypassable = slots_15_io_out_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_15_out_uop_exc_cause = slots_15_io_out_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_exception = slots_15_io_out_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_15_out_uop_stale_pdst = slots_15_io_out_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_ppred_busy = slots_15_io_out_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_prs3_busy = slots_15_io_out_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_prs2_busy = slots_15_io_out_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_prs1_busy = slots_15_io_out_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_15_out_uop_ppred = slots_15_io_out_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_15_out_uop_prs3 = slots_15_io_out_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_15_out_uop_prs2 = slots_15_io_out_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_15_out_uop_prs1 = slots_15_io_out_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_15_out_uop_pdst = slots_15_io_out_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_out_uop_rxq_idx = slots_15_io_out_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_15_out_uop_stq_idx = slots_15_io_out_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_15_out_uop_ldq_idx = slots_15_io_out_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_out_uop_rob_idx = slots_15_io_out_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_15_out_uop_csr_addr = slots_15_io_out_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_15_out_uop_imm_packed = slots_15_io_out_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_taken = slots_15_io_out_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_out_uop_pc_lob = slots_15_io_out_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_edge_inst = slots_15_io_out_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_15_out_uop_ftq_idx = slots_15_io_out_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_out_uop_br_tag = slots_15_io_out_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_15_out_uop_br_mask = slots_15_io_out_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_sfb = slots_15_io_out_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_jal = slots_15_io_out_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_jalr = slots_15_io_out_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_br = slots_15_io_out_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_iw_p2_poisoned = slots_15_io_out_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_iw_p1_poisoned = slots_15_io_out_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_out_uop_iw_state = slots_15_io_out_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_out_uop_ctrl_op3_sel = slots_15_io_out_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_ctrl_is_std = slots_15_io_out_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_ctrl_is_sta = slots_15_io_out_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_ctrl_is_load = slots_15_io_out_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_15_out_uop_ctrl_csr_cmd = slots_15_io_out_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_ctrl_fcn_dw = slots_15_io_out_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_out_uop_ctrl_op_fcn = slots_15_io_out_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_15_out_uop_ctrl_imm_sel = slots_15_io_out_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_15_out_uop_ctrl_op2_sel = slots_15_io_out_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_out_uop_ctrl_op1_sel = slots_15_io_out_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_out_uop_ctrl_br_type = slots_15_io_out_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [9:0] issue_slots_15_out_uop_fu_code = slots_15_io_out_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_15_out_uop_iq_type = slots_15_io_out_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_15_out_uop_debug_pc = slots_15_io_out_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_rvc = slots_15_io_out_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_15_out_uop_debug_inst = slots_15_io_out_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_15_out_uop_inst = slots_15_io_out_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_15_out_uop_uopc = slots_15_io_out_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_out_uop_address_num = slots_15_io_out_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_out_uop_rob_inst_idx = slots_15_io_out_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_out_uop_self_index = slots_15_io_out_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_out_uop_split_num = slots_15_io_out_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_out_uop_op2_sel = slots_15_io_out_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_out_uop_op1_sel = slots_15_io_out_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_out_uop_stale_pflag = slots_15_io_out_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_pflag_busy = slots_15_io_out_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_out_uop_pwflag = slots_15_io_out_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_out_uop_prflag = slots_15_io_out_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_wflag = slots_15_io_out_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_rflag = slots_15_io_out_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_out_uop_lrs3_rtype = slots_15_io_out_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_15_out_uop_shift = slots_15_io_out_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_is_unicore = slots_15_io_out_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_switch_off = slots_15_io_out_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_out_uop_switch = slots_15_io_out_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_13_clear = _GEN_29[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_2782 = _GEN_33[1:0] == 2'h1 & issue_slots_15_will_be_valid; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_14_in_uop_valid = _GEN_35[1:0] == 2'h2 ? will_be_valid_16 : _GEN_2782; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire  issue_slots_14_clear = _GEN_31[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  _GEN_2978 = _GEN_35[1:0] == 2'h1 & will_be_valid_16; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37 issue-unit-age-ordered.scala 68:33]
  wire  issue_slots_15_in_uop_valid = _GEN_37[1:0] == 2'h2 ? will_be_valid_17 : _GEN_2978; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  wire  issue_slots_15_clear = _GEN_33[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  wire  issue_slots_0_will_be_valid = slots_0_io_will_be_valid; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  will_be_available_0 = ~issue_slots_0_will_be_valid & ~issue_slots_0_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_1 = (~issue_slots_1_will_be_valid | issue_slots_1_clear) & ~issue_slots_1_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_2 = (~issue_slots_2_will_be_valid | issue_slots_2_clear) & ~issue_slots_2_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_3 = (~issue_slots_3_will_be_valid | issue_slots_3_clear) & ~issue_slots_3_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_4 = (~issue_slots_4_will_be_valid | issue_slots_4_clear) & ~issue_slots_4_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_5 = (~issue_slots_5_will_be_valid | issue_slots_5_clear) & ~issue_slots_5_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_6 = (~issue_slots_6_will_be_valid | issue_slots_6_clear) & ~issue_slots_6_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_7 = (~issue_slots_7_will_be_valid | issue_slots_7_clear) & ~issue_slots_7_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_8 = (~issue_slots_8_will_be_valid | issue_slots_8_clear) & ~issue_slots_8_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_9 = (~issue_slots_9_will_be_valid | issue_slots_9_clear) & ~issue_slots_9_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_10 = (~issue_slots_10_will_be_valid | issue_slots_10_clear) & ~issue_slots_10_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_11 = (~issue_slots_11_will_be_valid | issue_slots_11_clear) & ~issue_slots_11_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_12 = (~issue_slots_12_will_be_valid | issue_slots_12_clear) & ~issue_slots_12_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_13 = (~issue_slots_13_will_be_valid | issue_slots_13_clear) & ~issue_slots_13_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_14 = (~issue_slots_14_will_be_valid | issue_slots_14_clear) & ~issue_slots_14_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire  will_be_available_15 = (~issue_slots_15_will_be_valid | issue_slots_15_clear) & ~issue_slots_15_in_uop_valid; // @[issue-unit-age-ordered.scala 84:85]
  wire [1:0] _T_301 = will_be_available_0 + will_be_available_1; // @[Bitwise.scala 47:55]
  wire [1:0] _T_303 = will_be_available_2 + will_be_available_3; // @[Bitwise.scala 47:55]
  wire [2:0] _T_305 = _T_301 + _T_303; // @[Bitwise.scala 47:55]
  wire [1:0] _T_307 = will_be_available_4 + will_be_available_5; // @[Bitwise.scala 47:55]
  wire [1:0] _T_309 = will_be_available_6 + will_be_available_7; // @[Bitwise.scala 47:55]
  wire [2:0] _T_311 = _T_307 + _T_309; // @[Bitwise.scala 47:55]
  wire [3:0] _T_313 = _T_305 + _T_311; // @[Bitwise.scala 47:55]
  wire [1:0] _T_315 = will_be_available_8 + will_be_available_9; // @[Bitwise.scala 47:55]
  wire [1:0] _T_317 = will_be_available_10 + will_be_available_11; // @[Bitwise.scala 47:55]
  wire [2:0] _T_319 = _T_315 + _T_317; // @[Bitwise.scala 47:55]
  wire [1:0] _T_321 = will_be_available_12 + will_be_available_13; // @[Bitwise.scala 47:55]
  wire [1:0] _T_323 = will_be_available_14 + will_be_available_15; // @[Bitwise.scala 47:55]
  wire [2:0] _T_325 = _T_321 + _T_323; // @[Bitwise.scala 47:55]
  wire [3:0] _T_327 = _T_319 + _T_325; // @[Bitwise.scala 47:55]
  wire [4:0] num_available = _T_313 + _T_327; // @[Bitwise.scala 47:55]
  reg  REG; // @[issue-unit-age-ordered.scala 87:36]
  reg  REG_1; // @[issue-unit-age-ordered.scala 87:36]
  wire [1:0] issue_slots_0_uop_debug_tsrc = slots_0_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3175 = issue_slots_0_grant ? issue_slots_0_uop_debug_tsrc : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_0_uop_debug_fsrc = slots_0_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3176 = issue_slots_0_grant ? issue_slots_0_uop_debug_fsrc : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_bp_xcpt_if = slots_0_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3177 = issue_slots_0_grant & issue_slots_0_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_bp_debug_if = slots_0_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3178 = issue_slots_0_grant & issue_slots_0_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_xcpt_ma_if = slots_0_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3179 = issue_slots_0_grant & issue_slots_0_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_xcpt_ae_if = slots_0_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3180 = issue_slots_0_grant & issue_slots_0_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_xcpt_pf_if = slots_0_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3181 = issue_slots_0_grant & issue_slots_0_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_fp_single = slots_0_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3182 = issue_slots_0_grant & issue_slots_0_uop_fp_single; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_fp_val = slots_0_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3183 = issue_slots_0_grant & issue_slots_0_uop_fp_val; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_frs3_en = slots_0_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3184 = issue_slots_0_grant & issue_slots_0_uop_frs3_en; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_0_uop_lrs2_rtype = slots_0_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3185 = issue_slots_0_grant ? issue_slots_0_uop_lrs2_rtype : 2'h2; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 102:31]
  wire [1:0] issue_slots_0_uop_lrs1_rtype = slots_0_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3186 = issue_slots_0_grant ? issue_slots_0_uop_lrs1_rtype : 2'h2; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 101:31]
  wire [1:0] issue_slots_0_uop_dst_rtype = slots_0_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3187 = issue_slots_0_grant ? issue_slots_0_uop_dst_rtype : 2'h2; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_ldst_val = slots_0_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3188 = issue_slots_0_grant & issue_slots_0_uop_ldst_val; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_lrs3 = slots_0_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3189 = issue_slots_0_grant ? issue_slots_0_uop_lrs3 : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_lrs2 = slots_0_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3190 = issue_slots_0_grant ? issue_slots_0_uop_lrs2 : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_lrs1 = slots_0_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3191 = issue_slots_0_grant ? issue_slots_0_uop_lrs1 : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_ldst = slots_0_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3192 = issue_slots_0_grant ? issue_slots_0_uop_ldst : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_ldst_is_rs1 = slots_0_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3193 = issue_slots_0_grant & issue_slots_0_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_flush_on_commit = slots_0_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3194 = issue_slots_0_grant & issue_slots_0_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_unique = slots_0_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3195 = issue_slots_0_grant & issue_slots_0_uop_is_unique; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_sys_pc2epc = slots_0_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3196 = issue_slots_0_grant & issue_slots_0_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_uses_stq = slots_0_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3197 = issue_slots_0_grant & issue_slots_0_uop_uses_stq; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_uses_ldq = slots_0_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3198 = issue_slots_0_grant & issue_slots_0_uop_uses_ldq; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_amo = slots_0_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3199 = issue_slots_0_grant & issue_slots_0_uop_is_amo; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_fencei = slots_0_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3200 = issue_slots_0_grant & issue_slots_0_uop_is_fencei; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_fence = slots_0_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3201 = issue_slots_0_grant & issue_slots_0_uop_is_fence; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_mem_signed = slots_0_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3202 = issue_slots_0_grant & issue_slots_0_uop_mem_signed; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_0_uop_mem_size = slots_0_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3203 = issue_slots_0_grant ? issue_slots_0_uop_mem_size : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [4:0] issue_slots_0_uop_mem_cmd = slots_0_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3204 = issue_slots_0_grant ? issue_slots_0_uop_mem_cmd : 5'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_bypassable = slots_0_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3205 = issue_slots_0_grant & issue_slots_0_uop_bypassable; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [63:0] issue_slots_0_uop_exc_cause = slots_0_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_3206 = issue_slots_0_grant ? issue_slots_0_uop_exc_cause : 64'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_exception = slots_0_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3207 = issue_slots_0_grant & issue_slots_0_uop_exception; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [6:0] issue_slots_0_uop_stale_pdst = slots_0_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3208 = issue_slots_0_grant ? issue_slots_0_uop_stale_pdst : 7'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_ppred_busy = slots_0_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3209 = issue_slots_0_grant & issue_slots_0_uop_ppred_busy; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_prs3_busy = slots_0_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3210 = issue_slots_0_grant & issue_slots_0_uop_prs3_busy; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_prs2_busy = slots_0_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3211 = issue_slots_0_grant & issue_slots_0_uop_prs2_busy; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_prs1_busy = slots_0_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3212 = issue_slots_0_grant & issue_slots_0_uop_prs1_busy; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [4:0] issue_slots_0_uop_ppred = slots_0_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3213 = issue_slots_0_grant ? issue_slots_0_uop_ppred : 5'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [6:0] issue_slots_0_uop_prs3 = slots_0_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3214 = issue_slots_0_grant ? issue_slots_0_uop_prs3 : 7'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 100:25]
  wire [6:0] issue_slots_0_uop_prs2 = slots_0_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3215 = issue_slots_0_grant ? issue_slots_0_uop_prs2 : 7'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 99:25]
  wire [6:0] issue_slots_0_uop_prs1 = slots_0_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3216 = issue_slots_0_grant ? issue_slots_0_uop_prs1 : 7'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 98:25]
  wire [6:0] issue_slots_0_uop_pdst = slots_0_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3217 = issue_slots_0_grant ? issue_slots_0_uop_pdst : 7'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_0_uop_rxq_idx = slots_0_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3218 = issue_slots_0_grant ? issue_slots_0_uop_rxq_idx : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [4:0] issue_slots_0_uop_stq_idx = slots_0_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3219 = issue_slots_0_grant ? issue_slots_0_uop_stq_idx : 5'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [4:0] issue_slots_0_uop_ldq_idx = slots_0_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3220 = issue_slots_0_grant ? issue_slots_0_uop_ldq_idx : 5'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_rob_idx = slots_0_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3221 = issue_slots_0_grant ? issue_slots_0_uop_rob_idx : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [11:0] issue_slots_0_uop_csr_addr = slots_0_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_3222 = issue_slots_0_grant ? issue_slots_0_uop_csr_addr : 12'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [19:0] issue_slots_0_uop_imm_packed = slots_0_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_3223 = issue_slots_0_grant ? issue_slots_0_uop_imm_packed : 20'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_taken = slots_0_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3224 = issue_slots_0_grant & issue_slots_0_uop_taken; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_pc_lob = slots_0_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3225 = issue_slots_0_grant ? issue_slots_0_uop_pc_lob : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_edge_inst = slots_0_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3226 = issue_slots_0_grant & issue_slots_0_uop_edge_inst; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [4:0] issue_slots_0_uop_ftq_idx = slots_0_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3227 = issue_slots_0_grant ? issue_slots_0_uop_ftq_idx : 5'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] issue_slots_0_uop_br_tag = slots_0_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3228 = issue_slots_0_grant ? issue_slots_0_uop_br_tag : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [11:0] issue_slots_0_uop_br_mask = slots_0_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_3229 = issue_slots_0_grant ? issue_slots_0_uop_br_mask : 12'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_sfb = slots_0_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3230 = issue_slots_0_grant & issue_slots_0_uop_is_sfb; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_jal = slots_0_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3231 = issue_slots_0_grant & issue_slots_0_uop_is_jal; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_jalr = slots_0_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3232 = issue_slots_0_grant & issue_slots_0_uop_is_jalr; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_br = slots_0_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3233 = issue_slots_0_grant & issue_slots_0_uop_is_br; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_iw_p2_poisoned = slots_0_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3234 = issue_slots_0_grant & issue_slots_0_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_iw_p1_poisoned = slots_0_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3235 = issue_slots_0_grant & issue_slots_0_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_0_uop_iw_state = slots_0_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3236 = issue_slots_0_grant ? issue_slots_0_uop_iw_state : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_0_uop_ctrl_op3_sel = slots_0_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3237 = issue_slots_0_grant ? issue_slots_0_uop_ctrl_op3_sel : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_ctrl_is_std = slots_0_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3238 = issue_slots_0_grant & issue_slots_0_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_ctrl_is_sta = slots_0_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3239 = issue_slots_0_grant & issue_slots_0_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_ctrl_is_load = slots_0_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3240 = issue_slots_0_grant & issue_slots_0_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [2:0] issue_slots_0_uop_ctrl_csr_cmd = slots_0_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3241 = issue_slots_0_grant ? issue_slots_0_uop_ctrl_csr_cmd : 3'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_ctrl_fcn_dw = slots_0_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3242 = issue_slots_0_grant & issue_slots_0_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] issue_slots_0_uop_ctrl_op_fcn = slots_0_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3243 = issue_slots_0_grant ? issue_slots_0_uop_ctrl_op_fcn : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [2:0] issue_slots_0_uop_ctrl_imm_sel = slots_0_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3244 = issue_slots_0_grant ? issue_slots_0_uop_ctrl_imm_sel : 3'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [2:0] issue_slots_0_uop_ctrl_op2_sel = slots_0_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3245 = issue_slots_0_grant ? issue_slots_0_uop_ctrl_op2_sel : 3'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_0_uop_ctrl_op1_sel = slots_0_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3246 = issue_slots_0_grant ? issue_slots_0_uop_ctrl_op1_sel : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] issue_slots_0_uop_ctrl_br_type = slots_0_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3247 = issue_slots_0_grant ? issue_slots_0_uop_ctrl_br_type : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [9:0] _GEN_3248 = issue_slots_0_grant ? issue_slots_0_uop_fu_code : 10'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [2:0] issue_slots_0_uop_iq_type = slots_0_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3249 = issue_slots_0_grant ? issue_slots_0_uop_iq_type : 3'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [39:0] issue_slots_0_uop_debug_pc = slots_0_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_3250 = issue_slots_0_grant ? issue_slots_0_uop_debug_pc : 40'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_rvc = slots_0_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3251 = issue_slots_0_grant & issue_slots_0_uop_is_rvc; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [31:0] issue_slots_0_uop_debug_inst = slots_0_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_3252 = issue_slots_0_grant ? issue_slots_0_uop_debug_inst : 32'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [31:0] issue_slots_0_uop_inst = slots_0_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_3253 = issue_slots_0_grant ? issue_slots_0_uop_inst : 32'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [6:0] issue_slots_0_uop_uopc = slots_0_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3254 = issue_slots_0_grant ? issue_slots_0_uop_uopc : 7'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_address_num = slots_0_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3255 = issue_slots_0_grant ? issue_slots_0_uop_address_num : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_rob_inst_idx = slots_0_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3256 = issue_slots_0_grant ? issue_slots_0_uop_rob_inst_idx : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_self_index = slots_0_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3257 = issue_slots_0_grant ? issue_slots_0_uop_self_index : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [5:0] issue_slots_0_uop_split_num = slots_0_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3258 = issue_slots_0_grant ? issue_slots_0_uop_split_num : 6'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] issue_slots_0_uop_op2_sel = slots_0_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3259 = issue_slots_0_grant ? issue_slots_0_uop_op2_sel : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] issue_slots_0_uop_op1_sel = slots_0_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3260 = issue_slots_0_grant ? issue_slots_0_uop_op1_sel : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] issue_slots_0_uop_stale_pflag = slots_0_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3261 = issue_slots_0_grant ? issue_slots_0_uop_stale_pflag : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_pflag_busy = slots_0_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3262 = issue_slots_0_grant & issue_slots_0_uop_pflag_busy; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] issue_slots_0_uop_pwflag = slots_0_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3263 = issue_slots_0_grant ? issue_slots_0_uop_pwflag : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [3:0] issue_slots_0_uop_prflag = slots_0_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3264 = issue_slots_0_grant ? issue_slots_0_uop_prflag : 4'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 105:27]
  wire  issue_slots_0_uop_wflag = slots_0_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3265 = issue_slots_0_grant & issue_slots_0_uop_wflag; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_rflag = slots_0_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3266 = issue_slots_0_grant & issue_slots_0_uop_rflag; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 106:26]
  wire [1:0] issue_slots_0_uop_lrs3_rtype = slots_0_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3267 = issue_slots_0_grant ? issue_slots_0_uop_lrs3_rtype : 2'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [2:0] issue_slots_0_uop_shift = slots_0_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3268 = issue_slots_0_grant ? issue_slots_0_uop_shift : 3'h0; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_is_unicore = slots_0_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3269 = issue_slots_0_grant & issue_slots_0_uop_is_unicore; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_switch_off = slots_0_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3270 = issue_slots_0_grant & issue_slots_0_uop_switch_off; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire  issue_slots_0_uop_switch = slots_0_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3271 = issue_slots_0_grant & issue_slots_0_uop_switch; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24 issue-unit-age-ordered.scala 96:22]
  wire [1:0] issue_slots_1_uop_debug_tsrc = slots_1_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3274 = issue_slots_1_grant ? issue_slots_1_uop_debug_tsrc : _GEN_3175; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_1_uop_debug_fsrc = slots_1_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3275 = issue_slots_1_grant ? issue_slots_1_uop_debug_fsrc : _GEN_3176; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_bp_xcpt_if = slots_1_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3276 = issue_slots_1_grant ? issue_slots_1_uop_bp_xcpt_if : _GEN_3177; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_bp_debug_if = slots_1_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3277 = issue_slots_1_grant ? issue_slots_1_uop_bp_debug_if : _GEN_3178; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_xcpt_ma_if = slots_1_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3278 = issue_slots_1_grant ? issue_slots_1_uop_xcpt_ma_if : _GEN_3179; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_xcpt_ae_if = slots_1_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3279 = issue_slots_1_grant ? issue_slots_1_uop_xcpt_ae_if : _GEN_3180; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_xcpt_pf_if = slots_1_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3280 = issue_slots_1_grant ? issue_slots_1_uop_xcpt_pf_if : _GEN_3181; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_fp_single = slots_1_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3281 = issue_slots_1_grant ? issue_slots_1_uop_fp_single : _GEN_3182; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_fp_val = slots_1_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3282 = issue_slots_1_grant ? issue_slots_1_uop_fp_val : _GEN_3183; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_frs3_en = slots_1_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3283 = issue_slots_1_grant ? issue_slots_1_uop_frs3_en : _GEN_3184; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_1_uop_lrs2_rtype = slots_1_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3284 = issue_slots_1_grant ? issue_slots_1_uop_lrs2_rtype : _GEN_3185; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_1_uop_lrs1_rtype = slots_1_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3285 = issue_slots_1_grant ? issue_slots_1_uop_lrs1_rtype : _GEN_3186; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_1_uop_dst_rtype = slots_1_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3286 = issue_slots_1_grant ? issue_slots_1_uop_dst_rtype : _GEN_3187; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_ldst_val = slots_1_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3287 = issue_slots_1_grant ? issue_slots_1_uop_ldst_val : _GEN_3188; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_1_uop_lrs3 = slots_1_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3288 = issue_slots_1_grant ? issue_slots_1_uop_lrs3 : _GEN_3189; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_1_uop_lrs2 = slots_1_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3289 = issue_slots_1_grant ? issue_slots_1_uop_lrs2 : _GEN_3190; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_1_uop_lrs1 = slots_1_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3290 = issue_slots_1_grant ? issue_slots_1_uop_lrs1 : _GEN_3191; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_1_uop_ldst = slots_1_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3291 = issue_slots_1_grant ? issue_slots_1_uop_ldst : _GEN_3192; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_ldst_is_rs1 = slots_1_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3292 = issue_slots_1_grant ? issue_slots_1_uop_ldst_is_rs1 : _GEN_3193; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_flush_on_commit = slots_1_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3293 = issue_slots_1_grant ? issue_slots_1_uop_flush_on_commit : _GEN_3194; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_unique = slots_1_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3294 = issue_slots_1_grant ? issue_slots_1_uop_is_unique : _GEN_3195; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_sys_pc2epc = slots_1_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3295 = issue_slots_1_grant ? issue_slots_1_uop_is_sys_pc2epc : _GEN_3196; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_uses_stq = slots_1_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3296 = issue_slots_1_grant ? issue_slots_1_uop_uses_stq : _GEN_3197; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_uses_ldq = slots_1_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3297 = issue_slots_1_grant ? issue_slots_1_uop_uses_ldq : _GEN_3198; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_amo = slots_1_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3298 = issue_slots_1_grant ? issue_slots_1_uop_is_amo : _GEN_3199; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_fencei = slots_1_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3299 = issue_slots_1_grant ? issue_slots_1_uop_is_fencei : _GEN_3200; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_fence = slots_1_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3300 = issue_slots_1_grant ? issue_slots_1_uop_is_fence : _GEN_3201; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_mem_signed = slots_1_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3301 = issue_slots_1_grant ? issue_slots_1_uop_mem_signed : _GEN_3202; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_1_uop_mem_size = slots_1_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3302 = issue_slots_1_grant ? issue_slots_1_uop_mem_size : _GEN_3203; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_1_uop_mem_cmd = slots_1_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3303 = issue_slots_1_grant ? issue_slots_1_uop_mem_cmd : _GEN_3204; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_bypassable = slots_1_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3304 = issue_slots_1_grant ? issue_slots_1_uop_bypassable : _GEN_3205; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_1_uop_exc_cause = slots_1_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_3305 = issue_slots_1_grant ? issue_slots_1_uop_exc_cause : _GEN_3206; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_exception = slots_1_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3306 = issue_slots_1_grant ? issue_slots_1_uop_exception : _GEN_3207; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_1_uop_stale_pdst = slots_1_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3307 = issue_slots_1_grant ? issue_slots_1_uop_stale_pdst : _GEN_3208; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_ppred_busy = slots_1_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3308 = issue_slots_1_grant ? issue_slots_1_uop_ppred_busy : _GEN_3209; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_prs3_busy = slots_1_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3309 = issue_slots_1_grant ? issue_slots_1_uop_prs3_busy : _GEN_3210; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_prs2_busy = slots_1_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3310 = issue_slots_1_grant ? issue_slots_1_uop_prs2_busy : _GEN_3211; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_prs1_busy = slots_1_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3311 = issue_slots_1_grant ? issue_slots_1_uop_prs1_busy : _GEN_3212; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_1_uop_ppred = slots_1_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3312 = issue_slots_1_grant ? issue_slots_1_uop_ppred : _GEN_3213; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_1_uop_prs3 = slots_1_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3313 = issue_slots_1_grant ? issue_slots_1_uop_prs3 : _GEN_3214; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_1_uop_prs2 = slots_1_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3314 = issue_slots_1_grant ? issue_slots_1_uop_prs2 : _GEN_3215; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_1_uop_prs1 = slots_1_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3315 = issue_slots_1_grant ? issue_slots_1_uop_prs1 : _GEN_3216; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_1_uop_pdst = slots_1_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3316 = issue_slots_1_grant ? issue_slots_1_uop_pdst : _GEN_3217; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_1_uop_rxq_idx = slots_1_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3317 = issue_slots_1_grant ? issue_slots_1_uop_rxq_idx : _GEN_3218; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_1_uop_stq_idx = slots_1_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3318 = issue_slots_1_grant ? issue_slots_1_uop_stq_idx : _GEN_3219; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_1_uop_ldq_idx = slots_1_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3319 = issue_slots_1_grant ? issue_slots_1_uop_ldq_idx : _GEN_3220; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_1_uop_rob_idx = slots_1_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3320 = issue_slots_1_grant ? issue_slots_1_uop_rob_idx : _GEN_3221; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_1_uop_csr_addr = slots_1_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_3321 = issue_slots_1_grant ? issue_slots_1_uop_csr_addr : _GEN_3222; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_1_uop_imm_packed = slots_1_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_3322 = issue_slots_1_grant ? issue_slots_1_uop_imm_packed : _GEN_3223; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_taken = slots_1_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3323 = issue_slots_1_grant ? issue_slots_1_uop_taken : _GEN_3224; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_1_uop_pc_lob = slots_1_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3324 = issue_slots_1_grant ? issue_slots_1_uop_pc_lob : _GEN_3225; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_edge_inst = slots_1_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3325 = issue_slots_1_grant ? issue_slots_1_uop_edge_inst : _GEN_3226; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_1_uop_ftq_idx = slots_1_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3326 = issue_slots_1_grant ? issue_slots_1_uop_ftq_idx : _GEN_3227; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_1_uop_br_tag = slots_1_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3327 = issue_slots_1_grant ? issue_slots_1_uop_br_tag : _GEN_3228; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_1_uop_br_mask = slots_1_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_3328 = issue_slots_1_grant ? issue_slots_1_uop_br_mask : _GEN_3229; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_sfb = slots_1_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3329 = issue_slots_1_grant ? issue_slots_1_uop_is_sfb : _GEN_3230; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_jal = slots_1_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3330 = issue_slots_1_grant ? issue_slots_1_uop_is_jal : _GEN_3231; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_jalr = slots_1_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3331 = issue_slots_1_grant ? issue_slots_1_uop_is_jalr : _GEN_3232; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_br = slots_1_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3332 = issue_slots_1_grant ? issue_slots_1_uop_is_br : _GEN_3233; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_iw_p2_poisoned = slots_1_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3333 = issue_slots_1_grant ? issue_slots_1_uop_iw_p2_poisoned : _GEN_3234; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_iw_p1_poisoned = slots_1_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3334 = issue_slots_1_grant ? issue_slots_1_uop_iw_p1_poisoned : _GEN_3235; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_1_uop_iw_state = slots_1_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3335 = issue_slots_1_grant ? issue_slots_1_uop_iw_state : _GEN_3236; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_1_uop_ctrl_op3_sel = slots_1_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3336 = issue_slots_1_grant ? issue_slots_1_uop_ctrl_op3_sel : _GEN_3237; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_ctrl_is_std = slots_1_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3337 = issue_slots_1_grant ? issue_slots_1_uop_ctrl_is_std : _GEN_3238; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_ctrl_is_sta = slots_1_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3338 = issue_slots_1_grant ? issue_slots_1_uop_ctrl_is_sta : _GEN_3239; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_ctrl_is_load = slots_1_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3339 = issue_slots_1_grant ? issue_slots_1_uop_ctrl_is_load : _GEN_3240; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_1_uop_ctrl_csr_cmd = slots_1_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3340 = issue_slots_1_grant ? issue_slots_1_uop_ctrl_csr_cmd : _GEN_3241; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_ctrl_fcn_dw = slots_1_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3341 = issue_slots_1_grant ? issue_slots_1_uop_ctrl_fcn_dw : _GEN_3242; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_1_uop_ctrl_op_fcn = slots_1_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3342 = issue_slots_1_grant ? issue_slots_1_uop_ctrl_op_fcn : _GEN_3243; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_1_uop_ctrl_imm_sel = slots_1_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3343 = issue_slots_1_grant ? issue_slots_1_uop_ctrl_imm_sel : _GEN_3244; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_1_uop_ctrl_op2_sel = slots_1_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3344 = issue_slots_1_grant ? issue_slots_1_uop_ctrl_op2_sel : _GEN_3245; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_1_uop_ctrl_op1_sel = slots_1_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3345 = issue_slots_1_grant ? issue_slots_1_uop_ctrl_op1_sel : _GEN_3246; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_1_uop_ctrl_br_type = slots_1_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3346 = issue_slots_1_grant ? issue_slots_1_uop_ctrl_br_type : _GEN_3247; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_3347 = issue_slots_1_grant ? issue_slots_1_uop_fu_code : _GEN_3248; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_1_uop_iq_type = slots_1_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3348 = issue_slots_1_grant ? issue_slots_1_uop_iq_type : _GEN_3249; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_1_uop_debug_pc = slots_1_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_3349 = issue_slots_1_grant ? issue_slots_1_uop_debug_pc : _GEN_3250; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_rvc = slots_1_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3350 = issue_slots_1_grant ? issue_slots_1_uop_is_rvc : _GEN_3251; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_1_uop_debug_inst = slots_1_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_3351 = issue_slots_1_grant ? issue_slots_1_uop_debug_inst : _GEN_3252; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_1_uop_inst = slots_1_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_3352 = issue_slots_1_grant ? issue_slots_1_uop_inst : _GEN_3253; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_1_uop_uopc = slots_1_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3353 = issue_slots_1_grant ? issue_slots_1_uop_uopc : _GEN_3254; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_1_uop_address_num = slots_1_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3354 = issue_slots_1_grant ? issue_slots_1_uop_address_num : _GEN_3255; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_1_uop_rob_inst_idx = slots_1_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3355 = issue_slots_1_grant ? issue_slots_1_uop_rob_inst_idx : _GEN_3256; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_1_uop_self_index = slots_1_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3356 = issue_slots_1_grant ? issue_slots_1_uop_self_index : _GEN_3257; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_1_uop_split_num = slots_1_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3357 = issue_slots_1_grant ? issue_slots_1_uop_split_num : _GEN_3258; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_1_uop_op2_sel = slots_1_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3358 = issue_slots_1_grant ? issue_slots_1_uop_op2_sel : _GEN_3259; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_1_uop_op1_sel = slots_1_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3359 = issue_slots_1_grant ? issue_slots_1_uop_op1_sel : _GEN_3260; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_1_uop_stale_pflag = slots_1_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3360 = issue_slots_1_grant ? issue_slots_1_uop_stale_pflag : _GEN_3261; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_pflag_busy = slots_1_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3361 = issue_slots_1_grant ? issue_slots_1_uop_pflag_busy : _GEN_3262; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_1_uop_pwflag = slots_1_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3362 = issue_slots_1_grant ? issue_slots_1_uop_pwflag : _GEN_3263; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_1_uop_prflag = slots_1_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3363 = issue_slots_1_grant ? issue_slots_1_uop_prflag : _GEN_3264; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_wflag = slots_1_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3364 = issue_slots_1_grant ? issue_slots_1_uop_wflag : _GEN_3265; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_rflag = slots_1_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3365 = issue_slots_1_grant ? issue_slots_1_uop_rflag : _GEN_3266; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_1_uop_lrs3_rtype = slots_1_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3366 = issue_slots_1_grant ? issue_slots_1_uop_lrs3_rtype : _GEN_3267; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_1_uop_shift = slots_1_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3367 = issue_slots_1_grant ? issue_slots_1_uop_shift : _GEN_3268; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_is_unicore = slots_1_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3368 = issue_slots_1_grant ? issue_slots_1_uop_is_unicore : _GEN_3269; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_switch_off = slots_1_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3369 = issue_slots_1_grant ? issue_slots_1_uop_switch_off : _GEN_3270; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_1_uop_switch = slots_1_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3370 = issue_slots_1_grant ? issue_slots_1_uop_switch : _GEN_3271; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_debug_tsrc = slots_2_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3373 = issue_slots_2_grant ? issue_slots_2_uop_debug_tsrc : _GEN_3274; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_debug_fsrc = slots_2_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3374 = issue_slots_2_grant ? issue_slots_2_uop_debug_fsrc : _GEN_3275; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_bp_xcpt_if = slots_2_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3375 = issue_slots_2_grant ? issue_slots_2_uop_bp_xcpt_if : _GEN_3276; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_bp_debug_if = slots_2_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3376 = issue_slots_2_grant ? issue_slots_2_uop_bp_debug_if : _GEN_3277; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_xcpt_ma_if = slots_2_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3377 = issue_slots_2_grant ? issue_slots_2_uop_xcpt_ma_if : _GEN_3278; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_xcpt_ae_if = slots_2_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3378 = issue_slots_2_grant ? issue_slots_2_uop_xcpt_ae_if : _GEN_3279; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_xcpt_pf_if = slots_2_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3379 = issue_slots_2_grant ? issue_slots_2_uop_xcpt_pf_if : _GEN_3280; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_fp_single = slots_2_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3380 = issue_slots_2_grant ? issue_slots_2_uop_fp_single : _GEN_3281; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_fp_val = slots_2_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3381 = issue_slots_2_grant ? issue_slots_2_uop_fp_val : _GEN_3282; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_frs3_en = slots_2_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3382 = issue_slots_2_grant ? issue_slots_2_uop_frs3_en : _GEN_3283; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_lrs2_rtype = slots_2_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3383 = issue_slots_2_grant ? issue_slots_2_uop_lrs2_rtype : _GEN_3284; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_lrs1_rtype = slots_2_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3384 = issue_slots_2_grant ? issue_slots_2_uop_lrs1_rtype : _GEN_3285; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_dst_rtype = slots_2_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3385 = issue_slots_2_grant ? issue_slots_2_uop_dst_rtype : _GEN_3286; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_ldst_val = slots_2_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3386 = issue_slots_2_grant ? issue_slots_2_uop_ldst_val : _GEN_3287; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_2_uop_lrs3 = slots_2_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3387 = issue_slots_2_grant ? issue_slots_2_uop_lrs3 : _GEN_3288; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_2_uop_lrs2 = slots_2_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3388 = issue_slots_2_grant ? issue_slots_2_uop_lrs2 : _GEN_3289; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_2_uop_lrs1 = slots_2_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3389 = issue_slots_2_grant ? issue_slots_2_uop_lrs1 : _GEN_3290; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_2_uop_ldst = slots_2_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3390 = issue_slots_2_grant ? issue_slots_2_uop_ldst : _GEN_3291; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_ldst_is_rs1 = slots_2_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3391 = issue_slots_2_grant ? issue_slots_2_uop_ldst_is_rs1 : _GEN_3292; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_flush_on_commit = slots_2_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3392 = issue_slots_2_grant ? issue_slots_2_uop_flush_on_commit : _GEN_3293; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_unique = slots_2_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3393 = issue_slots_2_grant ? issue_slots_2_uop_is_unique : _GEN_3294; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_sys_pc2epc = slots_2_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3394 = issue_slots_2_grant ? issue_slots_2_uop_is_sys_pc2epc : _GEN_3295; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_uses_stq = slots_2_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3395 = issue_slots_2_grant ? issue_slots_2_uop_uses_stq : _GEN_3296; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_uses_ldq = slots_2_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3396 = issue_slots_2_grant ? issue_slots_2_uop_uses_ldq : _GEN_3297; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_amo = slots_2_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3397 = issue_slots_2_grant ? issue_slots_2_uop_is_amo : _GEN_3298; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_fencei = slots_2_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3398 = issue_slots_2_grant ? issue_slots_2_uop_is_fencei : _GEN_3299; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_fence = slots_2_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3399 = issue_slots_2_grant ? issue_slots_2_uop_is_fence : _GEN_3300; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_mem_signed = slots_2_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3400 = issue_slots_2_grant ? issue_slots_2_uop_mem_signed : _GEN_3301; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_mem_size = slots_2_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3401 = issue_slots_2_grant ? issue_slots_2_uop_mem_size : _GEN_3302; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_2_uop_mem_cmd = slots_2_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3402 = issue_slots_2_grant ? issue_slots_2_uop_mem_cmd : _GEN_3303; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_bypassable = slots_2_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3403 = issue_slots_2_grant ? issue_slots_2_uop_bypassable : _GEN_3304; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_2_uop_exc_cause = slots_2_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_3404 = issue_slots_2_grant ? issue_slots_2_uop_exc_cause : _GEN_3305; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_exception = slots_2_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3405 = issue_slots_2_grant ? issue_slots_2_uop_exception : _GEN_3306; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_2_uop_stale_pdst = slots_2_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3406 = issue_slots_2_grant ? issue_slots_2_uop_stale_pdst : _GEN_3307; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_ppred_busy = slots_2_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3407 = issue_slots_2_grant ? issue_slots_2_uop_ppred_busy : _GEN_3308; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_prs3_busy = slots_2_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3408 = issue_slots_2_grant ? issue_slots_2_uop_prs3_busy : _GEN_3309; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_prs2_busy = slots_2_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3409 = issue_slots_2_grant ? issue_slots_2_uop_prs2_busy : _GEN_3310; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_prs1_busy = slots_2_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3410 = issue_slots_2_grant ? issue_slots_2_uop_prs1_busy : _GEN_3311; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_2_uop_ppred = slots_2_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3411 = issue_slots_2_grant ? issue_slots_2_uop_ppred : _GEN_3312; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_2_uop_prs3 = slots_2_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3412 = issue_slots_2_grant ? issue_slots_2_uop_prs3 : _GEN_3313; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_2_uop_prs2 = slots_2_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3413 = issue_slots_2_grant ? issue_slots_2_uop_prs2 : _GEN_3314; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_2_uop_prs1 = slots_2_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3414 = issue_slots_2_grant ? issue_slots_2_uop_prs1 : _GEN_3315; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_2_uop_pdst = slots_2_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3415 = issue_slots_2_grant ? issue_slots_2_uop_pdst : _GEN_3316; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_rxq_idx = slots_2_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3416 = issue_slots_2_grant ? issue_slots_2_uop_rxq_idx : _GEN_3317; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_2_uop_stq_idx = slots_2_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3417 = issue_slots_2_grant ? issue_slots_2_uop_stq_idx : _GEN_3318; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_2_uop_ldq_idx = slots_2_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3418 = issue_slots_2_grant ? issue_slots_2_uop_ldq_idx : _GEN_3319; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_2_uop_rob_idx = slots_2_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3419 = issue_slots_2_grant ? issue_slots_2_uop_rob_idx : _GEN_3320; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_2_uop_csr_addr = slots_2_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_3420 = issue_slots_2_grant ? issue_slots_2_uop_csr_addr : _GEN_3321; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_2_uop_imm_packed = slots_2_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_3421 = issue_slots_2_grant ? issue_slots_2_uop_imm_packed : _GEN_3322; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_taken = slots_2_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3422 = issue_slots_2_grant ? issue_slots_2_uop_taken : _GEN_3323; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_2_uop_pc_lob = slots_2_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3423 = issue_slots_2_grant ? issue_slots_2_uop_pc_lob : _GEN_3324; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_edge_inst = slots_2_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3424 = issue_slots_2_grant ? issue_slots_2_uop_edge_inst : _GEN_3325; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_2_uop_ftq_idx = slots_2_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3425 = issue_slots_2_grant ? issue_slots_2_uop_ftq_idx : _GEN_3326; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_2_uop_br_tag = slots_2_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3426 = issue_slots_2_grant ? issue_slots_2_uop_br_tag : _GEN_3327; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_2_uop_br_mask = slots_2_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_3427 = issue_slots_2_grant ? issue_slots_2_uop_br_mask : _GEN_3328; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_sfb = slots_2_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3428 = issue_slots_2_grant ? issue_slots_2_uop_is_sfb : _GEN_3329; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_jal = slots_2_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3429 = issue_slots_2_grant ? issue_slots_2_uop_is_jal : _GEN_3330; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_jalr = slots_2_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3430 = issue_slots_2_grant ? issue_slots_2_uop_is_jalr : _GEN_3331; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_br = slots_2_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3431 = issue_slots_2_grant ? issue_slots_2_uop_is_br : _GEN_3332; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_iw_p2_poisoned = slots_2_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3432 = issue_slots_2_grant ? issue_slots_2_uop_iw_p2_poisoned : _GEN_3333; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_iw_p1_poisoned = slots_2_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3433 = issue_slots_2_grant ? issue_slots_2_uop_iw_p1_poisoned : _GEN_3334; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_iw_state = slots_2_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3434 = issue_slots_2_grant ? issue_slots_2_uop_iw_state : _GEN_3335; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_ctrl_op3_sel = slots_2_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3435 = issue_slots_2_grant ? issue_slots_2_uop_ctrl_op3_sel : _GEN_3336; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_ctrl_is_std = slots_2_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3436 = issue_slots_2_grant ? issue_slots_2_uop_ctrl_is_std : _GEN_3337; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_ctrl_is_sta = slots_2_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3437 = issue_slots_2_grant ? issue_slots_2_uop_ctrl_is_sta : _GEN_3338; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_ctrl_is_load = slots_2_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3438 = issue_slots_2_grant ? issue_slots_2_uop_ctrl_is_load : _GEN_3339; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_2_uop_ctrl_csr_cmd = slots_2_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3439 = issue_slots_2_grant ? issue_slots_2_uop_ctrl_csr_cmd : _GEN_3340; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_ctrl_fcn_dw = slots_2_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3440 = issue_slots_2_grant ? issue_slots_2_uop_ctrl_fcn_dw : _GEN_3341; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_2_uop_ctrl_op_fcn = slots_2_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3441 = issue_slots_2_grant ? issue_slots_2_uop_ctrl_op_fcn : _GEN_3342; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_2_uop_ctrl_imm_sel = slots_2_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3442 = issue_slots_2_grant ? issue_slots_2_uop_ctrl_imm_sel : _GEN_3343; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_2_uop_ctrl_op2_sel = slots_2_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3443 = issue_slots_2_grant ? issue_slots_2_uop_ctrl_op2_sel : _GEN_3344; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_ctrl_op1_sel = slots_2_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3444 = issue_slots_2_grant ? issue_slots_2_uop_ctrl_op1_sel : _GEN_3345; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_2_uop_ctrl_br_type = slots_2_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3445 = issue_slots_2_grant ? issue_slots_2_uop_ctrl_br_type : _GEN_3346; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_3446 = issue_slots_2_grant ? issue_slots_2_uop_fu_code : _GEN_3347; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_2_uop_iq_type = slots_2_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3447 = issue_slots_2_grant ? issue_slots_2_uop_iq_type : _GEN_3348; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_2_uop_debug_pc = slots_2_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_3448 = issue_slots_2_grant ? issue_slots_2_uop_debug_pc : _GEN_3349; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_rvc = slots_2_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3449 = issue_slots_2_grant ? issue_slots_2_uop_is_rvc : _GEN_3350; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_2_uop_debug_inst = slots_2_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_3450 = issue_slots_2_grant ? issue_slots_2_uop_debug_inst : _GEN_3351; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_2_uop_inst = slots_2_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_3451 = issue_slots_2_grant ? issue_slots_2_uop_inst : _GEN_3352; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_2_uop_uopc = slots_2_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3452 = issue_slots_2_grant ? issue_slots_2_uop_uopc : _GEN_3353; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_2_uop_address_num = slots_2_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3453 = issue_slots_2_grant ? issue_slots_2_uop_address_num : _GEN_3354; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_2_uop_rob_inst_idx = slots_2_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3454 = issue_slots_2_grant ? issue_slots_2_uop_rob_inst_idx : _GEN_3355; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_2_uop_self_index = slots_2_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3455 = issue_slots_2_grant ? issue_slots_2_uop_self_index : _GEN_3356; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_2_uop_split_num = slots_2_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3456 = issue_slots_2_grant ? issue_slots_2_uop_split_num : _GEN_3357; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_2_uop_op2_sel = slots_2_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3457 = issue_slots_2_grant ? issue_slots_2_uop_op2_sel : _GEN_3358; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_2_uop_op1_sel = slots_2_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3458 = issue_slots_2_grant ? issue_slots_2_uop_op1_sel : _GEN_3359; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_2_uop_stale_pflag = slots_2_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3459 = issue_slots_2_grant ? issue_slots_2_uop_stale_pflag : _GEN_3360; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_pflag_busy = slots_2_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3460 = issue_slots_2_grant ? issue_slots_2_uop_pflag_busy : _GEN_3361; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_2_uop_pwflag = slots_2_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3461 = issue_slots_2_grant ? issue_slots_2_uop_pwflag : _GEN_3362; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_2_uop_prflag = slots_2_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3462 = issue_slots_2_grant ? issue_slots_2_uop_prflag : _GEN_3363; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_wflag = slots_2_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3463 = issue_slots_2_grant ? issue_slots_2_uop_wflag : _GEN_3364; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_rflag = slots_2_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3464 = issue_slots_2_grant ? issue_slots_2_uop_rflag : _GEN_3365; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_2_uop_lrs3_rtype = slots_2_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3465 = issue_slots_2_grant ? issue_slots_2_uop_lrs3_rtype : _GEN_3366; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_2_uop_shift = slots_2_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3466 = issue_slots_2_grant ? issue_slots_2_uop_shift : _GEN_3367; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_is_unicore = slots_2_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3467 = issue_slots_2_grant ? issue_slots_2_uop_is_unicore : _GEN_3368; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_switch_off = slots_2_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3468 = issue_slots_2_grant ? issue_slots_2_uop_switch_off : _GEN_3369; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_2_uop_switch = slots_2_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3469 = issue_slots_2_grant ? issue_slots_2_uop_switch : _GEN_3370; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_debug_tsrc = slots_3_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3472 = issue_slots_3_grant ? issue_slots_3_uop_debug_tsrc : _GEN_3373; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_debug_fsrc = slots_3_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3473 = issue_slots_3_grant ? issue_slots_3_uop_debug_fsrc : _GEN_3374; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_bp_xcpt_if = slots_3_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3474 = issue_slots_3_grant ? issue_slots_3_uop_bp_xcpt_if : _GEN_3375; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_bp_debug_if = slots_3_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3475 = issue_slots_3_grant ? issue_slots_3_uop_bp_debug_if : _GEN_3376; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_xcpt_ma_if = slots_3_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3476 = issue_slots_3_grant ? issue_slots_3_uop_xcpt_ma_if : _GEN_3377; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_xcpt_ae_if = slots_3_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3477 = issue_slots_3_grant ? issue_slots_3_uop_xcpt_ae_if : _GEN_3378; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_xcpt_pf_if = slots_3_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3478 = issue_slots_3_grant ? issue_slots_3_uop_xcpt_pf_if : _GEN_3379; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_fp_single = slots_3_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3479 = issue_slots_3_grant ? issue_slots_3_uop_fp_single : _GEN_3380; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_fp_val = slots_3_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3480 = issue_slots_3_grant ? issue_slots_3_uop_fp_val : _GEN_3381; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_frs3_en = slots_3_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3481 = issue_slots_3_grant ? issue_slots_3_uop_frs3_en : _GEN_3382; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_lrs2_rtype = slots_3_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3482 = issue_slots_3_grant ? issue_slots_3_uop_lrs2_rtype : _GEN_3383; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_lrs1_rtype = slots_3_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3483 = issue_slots_3_grant ? issue_slots_3_uop_lrs1_rtype : _GEN_3384; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_dst_rtype = slots_3_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3484 = issue_slots_3_grant ? issue_slots_3_uop_dst_rtype : _GEN_3385; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_ldst_val = slots_3_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3485 = issue_slots_3_grant ? issue_slots_3_uop_ldst_val : _GEN_3386; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_3_uop_lrs3 = slots_3_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3486 = issue_slots_3_grant ? issue_slots_3_uop_lrs3 : _GEN_3387; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_3_uop_lrs2 = slots_3_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3487 = issue_slots_3_grant ? issue_slots_3_uop_lrs2 : _GEN_3388; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_3_uop_lrs1 = slots_3_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3488 = issue_slots_3_grant ? issue_slots_3_uop_lrs1 : _GEN_3389; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_3_uop_ldst = slots_3_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3489 = issue_slots_3_grant ? issue_slots_3_uop_ldst : _GEN_3390; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_ldst_is_rs1 = slots_3_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3490 = issue_slots_3_grant ? issue_slots_3_uop_ldst_is_rs1 : _GEN_3391; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_flush_on_commit = slots_3_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3491 = issue_slots_3_grant ? issue_slots_3_uop_flush_on_commit : _GEN_3392; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_unique = slots_3_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3492 = issue_slots_3_grant ? issue_slots_3_uop_is_unique : _GEN_3393; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_sys_pc2epc = slots_3_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3493 = issue_slots_3_grant ? issue_slots_3_uop_is_sys_pc2epc : _GEN_3394; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_uses_stq = slots_3_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3494 = issue_slots_3_grant ? issue_slots_3_uop_uses_stq : _GEN_3395; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_uses_ldq = slots_3_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3495 = issue_slots_3_grant ? issue_slots_3_uop_uses_ldq : _GEN_3396; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_amo = slots_3_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3496 = issue_slots_3_grant ? issue_slots_3_uop_is_amo : _GEN_3397; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_fencei = slots_3_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3497 = issue_slots_3_grant ? issue_slots_3_uop_is_fencei : _GEN_3398; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_fence = slots_3_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3498 = issue_slots_3_grant ? issue_slots_3_uop_is_fence : _GEN_3399; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_mem_signed = slots_3_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3499 = issue_slots_3_grant ? issue_slots_3_uop_mem_signed : _GEN_3400; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_mem_size = slots_3_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3500 = issue_slots_3_grant ? issue_slots_3_uop_mem_size : _GEN_3401; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_3_uop_mem_cmd = slots_3_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3501 = issue_slots_3_grant ? issue_slots_3_uop_mem_cmd : _GEN_3402; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_bypassable = slots_3_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3502 = issue_slots_3_grant ? issue_slots_3_uop_bypassable : _GEN_3403; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_3_uop_exc_cause = slots_3_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_3503 = issue_slots_3_grant ? issue_slots_3_uop_exc_cause : _GEN_3404; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_exception = slots_3_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3504 = issue_slots_3_grant ? issue_slots_3_uop_exception : _GEN_3405; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_3_uop_stale_pdst = slots_3_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3505 = issue_slots_3_grant ? issue_slots_3_uop_stale_pdst : _GEN_3406; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_ppred_busy = slots_3_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3506 = issue_slots_3_grant ? issue_slots_3_uop_ppred_busy : _GEN_3407; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_prs3_busy = slots_3_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3507 = issue_slots_3_grant ? issue_slots_3_uop_prs3_busy : _GEN_3408; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_prs2_busy = slots_3_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3508 = issue_slots_3_grant ? issue_slots_3_uop_prs2_busy : _GEN_3409; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_prs1_busy = slots_3_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3509 = issue_slots_3_grant ? issue_slots_3_uop_prs1_busy : _GEN_3410; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_3_uop_ppred = slots_3_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3510 = issue_slots_3_grant ? issue_slots_3_uop_ppred : _GEN_3411; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_3_uop_prs3 = slots_3_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3511 = issue_slots_3_grant ? issue_slots_3_uop_prs3 : _GEN_3412; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_3_uop_prs2 = slots_3_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3512 = issue_slots_3_grant ? issue_slots_3_uop_prs2 : _GEN_3413; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_3_uop_prs1 = slots_3_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3513 = issue_slots_3_grant ? issue_slots_3_uop_prs1 : _GEN_3414; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_3_uop_pdst = slots_3_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3514 = issue_slots_3_grant ? issue_slots_3_uop_pdst : _GEN_3415; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_rxq_idx = slots_3_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3515 = issue_slots_3_grant ? issue_slots_3_uop_rxq_idx : _GEN_3416; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_3_uop_stq_idx = slots_3_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3516 = issue_slots_3_grant ? issue_slots_3_uop_stq_idx : _GEN_3417; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_3_uop_ldq_idx = slots_3_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3517 = issue_slots_3_grant ? issue_slots_3_uop_ldq_idx : _GEN_3418; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_3_uop_rob_idx = slots_3_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3518 = issue_slots_3_grant ? issue_slots_3_uop_rob_idx : _GEN_3419; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_3_uop_csr_addr = slots_3_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_3519 = issue_slots_3_grant ? issue_slots_3_uop_csr_addr : _GEN_3420; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_3_uop_imm_packed = slots_3_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_3520 = issue_slots_3_grant ? issue_slots_3_uop_imm_packed : _GEN_3421; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_taken = slots_3_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3521 = issue_slots_3_grant ? issue_slots_3_uop_taken : _GEN_3422; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_3_uop_pc_lob = slots_3_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3522 = issue_slots_3_grant ? issue_slots_3_uop_pc_lob : _GEN_3423; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_edge_inst = slots_3_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3523 = issue_slots_3_grant ? issue_slots_3_uop_edge_inst : _GEN_3424; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_3_uop_ftq_idx = slots_3_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3524 = issue_slots_3_grant ? issue_slots_3_uop_ftq_idx : _GEN_3425; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_3_uop_br_tag = slots_3_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3525 = issue_slots_3_grant ? issue_slots_3_uop_br_tag : _GEN_3426; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_3_uop_br_mask = slots_3_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_3526 = issue_slots_3_grant ? issue_slots_3_uop_br_mask : _GEN_3427; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_sfb = slots_3_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3527 = issue_slots_3_grant ? issue_slots_3_uop_is_sfb : _GEN_3428; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_jal = slots_3_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3528 = issue_slots_3_grant ? issue_slots_3_uop_is_jal : _GEN_3429; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_jalr = slots_3_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3529 = issue_slots_3_grant ? issue_slots_3_uop_is_jalr : _GEN_3430; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_br = slots_3_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3530 = issue_slots_3_grant ? issue_slots_3_uop_is_br : _GEN_3431; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_iw_p2_poisoned = slots_3_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3531 = issue_slots_3_grant ? issue_slots_3_uop_iw_p2_poisoned : _GEN_3432; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_iw_p1_poisoned = slots_3_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3532 = issue_slots_3_grant ? issue_slots_3_uop_iw_p1_poisoned : _GEN_3433; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_iw_state = slots_3_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3533 = issue_slots_3_grant ? issue_slots_3_uop_iw_state : _GEN_3434; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_ctrl_op3_sel = slots_3_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3534 = issue_slots_3_grant ? issue_slots_3_uop_ctrl_op3_sel : _GEN_3435; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_ctrl_is_std = slots_3_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3535 = issue_slots_3_grant ? issue_slots_3_uop_ctrl_is_std : _GEN_3436; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_ctrl_is_sta = slots_3_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3536 = issue_slots_3_grant ? issue_slots_3_uop_ctrl_is_sta : _GEN_3437; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_ctrl_is_load = slots_3_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3537 = issue_slots_3_grant ? issue_slots_3_uop_ctrl_is_load : _GEN_3438; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_3_uop_ctrl_csr_cmd = slots_3_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3538 = issue_slots_3_grant ? issue_slots_3_uop_ctrl_csr_cmd : _GEN_3439; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_ctrl_fcn_dw = slots_3_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3539 = issue_slots_3_grant ? issue_slots_3_uop_ctrl_fcn_dw : _GEN_3440; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_3_uop_ctrl_op_fcn = slots_3_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3540 = issue_slots_3_grant ? issue_slots_3_uop_ctrl_op_fcn : _GEN_3441; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_3_uop_ctrl_imm_sel = slots_3_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3541 = issue_slots_3_grant ? issue_slots_3_uop_ctrl_imm_sel : _GEN_3442; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_3_uop_ctrl_op2_sel = slots_3_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3542 = issue_slots_3_grant ? issue_slots_3_uop_ctrl_op2_sel : _GEN_3443; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_ctrl_op1_sel = slots_3_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3543 = issue_slots_3_grant ? issue_slots_3_uop_ctrl_op1_sel : _GEN_3444; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_3_uop_ctrl_br_type = slots_3_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3544 = issue_slots_3_grant ? issue_slots_3_uop_ctrl_br_type : _GEN_3445; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_3545 = issue_slots_3_grant ? issue_slots_3_uop_fu_code : _GEN_3446; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_3_uop_iq_type = slots_3_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3546 = issue_slots_3_grant ? issue_slots_3_uop_iq_type : _GEN_3447; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_3_uop_debug_pc = slots_3_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_3547 = issue_slots_3_grant ? issue_slots_3_uop_debug_pc : _GEN_3448; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_rvc = slots_3_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3548 = issue_slots_3_grant ? issue_slots_3_uop_is_rvc : _GEN_3449; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_3_uop_debug_inst = slots_3_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_3549 = issue_slots_3_grant ? issue_slots_3_uop_debug_inst : _GEN_3450; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_3_uop_inst = slots_3_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_3550 = issue_slots_3_grant ? issue_slots_3_uop_inst : _GEN_3451; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_3_uop_uopc = slots_3_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3551 = issue_slots_3_grant ? issue_slots_3_uop_uopc : _GEN_3452; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_3_uop_address_num = slots_3_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3552 = issue_slots_3_grant ? issue_slots_3_uop_address_num : _GEN_3453; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_3_uop_rob_inst_idx = slots_3_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3553 = issue_slots_3_grant ? issue_slots_3_uop_rob_inst_idx : _GEN_3454; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_3_uop_self_index = slots_3_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3554 = issue_slots_3_grant ? issue_slots_3_uop_self_index : _GEN_3455; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_3_uop_split_num = slots_3_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3555 = issue_slots_3_grant ? issue_slots_3_uop_split_num : _GEN_3456; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_3_uop_op2_sel = slots_3_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3556 = issue_slots_3_grant ? issue_slots_3_uop_op2_sel : _GEN_3457; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_3_uop_op1_sel = slots_3_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3557 = issue_slots_3_grant ? issue_slots_3_uop_op1_sel : _GEN_3458; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_3_uop_stale_pflag = slots_3_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3558 = issue_slots_3_grant ? issue_slots_3_uop_stale_pflag : _GEN_3459; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_pflag_busy = slots_3_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3559 = issue_slots_3_grant ? issue_slots_3_uop_pflag_busy : _GEN_3460; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_3_uop_pwflag = slots_3_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3560 = issue_slots_3_grant ? issue_slots_3_uop_pwflag : _GEN_3461; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_3_uop_prflag = slots_3_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3561 = issue_slots_3_grant ? issue_slots_3_uop_prflag : _GEN_3462; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_wflag = slots_3_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3562 = issue_slots_3_grant ? issue_slots_3_uop_wflag : _GEN_3463; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_rflag = slots_3_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3563 = issue_slots_3_grant ? issue_slots_3_uop_rflag : _GEN_3464; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_3_uop_lrs3_rtype = slots_3_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3564 = issue_slots_3_grant ? issue_slots_3_uop_lrs3_rtype : _GEN_3465; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_3_uop_shift = slots_3_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3565 = issue_slots_3_grant ? issue_slots_3_uop_shift : _GEN_3466; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_is_unicore = slots_3_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3566 = issue_slots_3_grant ? issue_slots_3_uop_is_unicore : _GEN_3467; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_switch_off = slots_3_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3567 = issue_slots_3_grant ? issue_slots_3_uop_switch_off : _GEN_3468; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_3_uop_switch = slots_3_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3568 = issue_slots_3_grant ? issue_slots_3_uop_switch : _GEN_3469; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_debug_tsrc = slots_4_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3571 = issue_slots_4_grant ? issue_slots_4_uop_debug_tsrc : _GEN_3472; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_debug_fsrc = slots_4_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3572 = issue_slots_4_grant ? issue_slots_4_uop_debug_fsrc : _GEN_3473; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_bp_xcpt_if = slots_4_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3573 = issue_slots_4_grant ? issue_slots_4_uop_bp_xcpt_if : _GEN_3474; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_bp_debug_if = slots_4_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3574 = issue_slots_4_grant ? issue_slots_4_uop_bp_debug_if : _GEN_3475; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_xcpt_ma_if = slots_4_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3575 = issue_slots_4_grant ? issue_slots_4_uop_xcpt_ma_if : _GEN_3476; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_xcpt_ae_if = slots_4_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3576 = issue_slots_4_grant ? issue_slots_4_uop_xcpt_ae_if : _GEN_3477; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_xcpt_pf_if = slots_4_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3577 = issue_slots_4_grant ? issue_slots_4_uop_xcpt_pf_if : _GEN_3478; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_fp_single = slots_4_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3578 = issue_slots_4_grant ? issue_slots_4_uop_fp_single : _GEN_3479; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_fp_val = slots_4_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3579 = issue_slots_4_grant ? issue_slots_4_uop_fp_val : _GEN_3480; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_frs3_en = slots_4_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3580 = issue_slots_4_grant ? issue_slots_4_uop_frs3_en : _GEN_3481; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_lrs2_rtype = slots_4_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3581 = issue_slots_4_grant ? issue_slots_4_uop_lrs2_rtype : _GEN_3482; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_lrs1_rtype = slots_4_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3582 = issue_slots_4_grant ? issue_slots_4_uop_lrs1_rtype : _GEN_3483; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_dst_rtype = slots_4_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3583 = issue_slots_4_grant ? issue_slots_4_uop_dst_rtype : _GEN_3484; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_ldst_val = slots_4_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3584 = issue_slots_4_grant ? issue_slots_4_uop_ldst_val : _GEN_3485; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_4_uop_lrs3 = slots_4_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3585 = issue_slots_4_grant ? issue_slots_4_uop_lrs3 : _GEN_3486; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_4_uop_lrs2 = slots_4_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3586 = issue_slots_4_grant ? issue_slots_4_uop_lrs2 : _GEN_3487; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_4_uop_lrs1 = slots_4_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3587 = issue_slots_4_grant ? issue_slots_4_uop_lrs1 : _GEN_3488; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_4_uop_ldst = slots_4_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3588 = issue_slots_4_grant ? issue_slots_4_uop_ldst : _GEN_3489; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_ldst_is_rs1 = slots_4_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3589 = issue_slots_4_grant ? issue_slots_4_uop_ldst_is_rs1 : _GEN_3490; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_flush_on_commit = slots_4_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3590 = issue_slots_4_grant ? issue_slots_4_uop_flush_on_commit : _GEN_3491; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_unique = slots_4_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3591 = issue_slots_4_grant ? issue_slots_4_uop_is_unique : _GEN_3492; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_sys_pc2epc = slots_4_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3592 = issue_slots_4_grant ? issue_slots_4_uop_is_sys_pc2epc : _GEN_3493; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_uses_stq = slots_4_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3593 = issue_slots_4_grant ? issue_slots_4_uop_uses_stq : _GEN_3494; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_uses_ldq = slots_4_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3594 = issue_slots_4_grant ? issue_slots_4_uop_uses_ldq : _GEN_3495; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_amo = slots_4_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3595 = issue_slots_4_grant ? issue_slots_4_uop_is_amo : _GEN_3496; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_fencei = slots_4_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3596 = issue_slots_4_grant ? issue_slots_4_uop_is_fencei : _GEN_3497; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_fence = slots_4_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3597 = issue_slots_4_grant ? issue_slots_4_uop_is_fence : _GEN_3498; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_mem_signed = slots_4_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3598 = issue_slots_4_grant ? issue_slots_4_uop_mem_signed : _GEN_3499; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_mem_size = slots_4_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3599 = issue_slots_4_grant ? issue_slots_4_uop_mem_size : _GEN_3500; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_4_uop_mem_cmd = slots_4_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3600 = issue_slots_4_grant ? issue_slots_4_uop_mem_cmd : _GEN_3501; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_bypassable = slots_4_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3601 = issue_slots_4_grant ? issue_slots_4_uop_bypassable : _GEN_3502; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_4_uop_exc_cause = slots_4_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_3602 = issue_slots_4_grant ? issue_slots_4_uop_exc_cause : _GEN_3503; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_exception = slots_4_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3603 = issue_slots_4_grant ? issue_slots_4_uop_exception : _GEN_3504; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_4_uop_stale_pdst = slots_4_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3604 = issue_slots_4_grant ? issue_slots_4_uop_stale_pdst : _GEN_3505; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_ppred_busy = slots_4_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3605 = issue_slots_4_grant ? issue_slots_4_uop_ppred_busy : _GEN_3506; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_prs3_busy = slots_4_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3606 = issue_slots_4_grant ? issue_slots_4_uop_prs3_busy : _GEN_3507; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_prs2_busy = slots_4_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3607 = issue_slots_4_grant ? issue_slots_4_uop_prs2_busy : _GEN_3508; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_prs1_busy = slots_4_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3608 = issue_slots_4_grant ? issue_slots_4_uop_prs1_busy : _GEN_3509; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_4_uop_ppred = slots_4_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3609 = issue_slots_4_grant ? issue_slots_4_uop_ppred : _GEN_3510; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_4_uop_prs3 = slots_4_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3610 = issue_slots_4_grant ? issue_slots_4_uop_prs3 : _GEN_3511; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_4_uop_prs2 = slots_4_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3611 = issue_slots_4_grant ? issue_slots_4_uop_prs2 : _GEN_3512; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_4_uop_prs1 = slots_4_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3612 = issue_slots_4_grant ? issue_slots_4_uop_prs1 : _GEN_3513; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_4_uop_pdst = slots_4_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3613 = issue_slots_4_grant ? issue_slots_4_uop_pdst : _GEN_3514; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_rxq_idx = slots_4_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3614 = issue_slots_4_grant ? issue_slots_4_uop_rxq_idx : _GEN_3515; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_4_uop_stq_idx = slots_4_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3615 = issue_slots_4_grant ? issue_slots_4_uop_stq_idx : _GEN_3516; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_4_uop_ldq_idx = slots_4_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3616 = issue_slots_4_grant ? issue_slots_4_uop_ldq_idx : _GEN_3517; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_4_uop_rob_idx = slots_4_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3617 = issue_slots_4_grant ? issue_slots_4_uop_rob_idx : _GEN_3518; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_4_uop_csr_addr = slots_4_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_3618 = issue_slots_4_grant ? issue_slots_4_uop_csr_addr : _GEN_3519; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_4_uop_imm_packed = slots_4_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_3619 = issue_slots_4_grant ? issue_slots_4_uop_imm_packed : _GEN_3520; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_taken = slots_4_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3620 = issue_slots_4_grant ? issue_slots_4_uop_taken : _GEN_3521; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_4_uop_pc_lob = slots_4_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3621 = issue_slots_4_grant ? issue_slots_4_uop_pc_lob : _GEN_3522; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_edge_inst = slots_4_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3622 = issue_slots_4_grant ? issue_slots_4_uop_edge_inst : _GEN_3523; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_4_uop_ftq_idx = slots_4_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3623 = issue_slots_4_grant ? issue_slots_4_uop_ftq_idx : _GEN_3524; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_4_uop_br_tag = slots_4_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3624 = issue_slots_4_grant ? issue_slots_4_uop_br_tag : _GEN_3525; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_4_uop_br_mask = slots_4_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_3625 = issue_slots_4_grant ? issue_slots_4_uop_br_mask : _GEN_3526; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_sfb = slots_4_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3626 = issue_slots_4_grant ? issue_slots_4_uop_is_sfb : _GEN_3527; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_jal = slots_4_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3627 = issue_slots_4_grant ? issue_slots_4_uop_is_jal : _GEN_3528; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_jalr = slots_4_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3628 = issue_slots_4_grant ? issue_slots_4_uop_is_jalr : _GEN_3529; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_br = slots_4_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3629 = issue_slots_4_grant ? issue_slots_4_uop_is_br : _GEN_3530; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_iw_p2_poisoned = slots_4_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3630 = issue_slots_4_grant ? issue_slots_4_uop_iw_p2_poisoned : _GEN_3531; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_iw_p1_poisoned = slots_4_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3631 = issue_slots_4_grant ? issue_slots_4_uop_iw_p1_poisoned : _GEN_3532; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_iw_state = slots_4_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3632 = issue_slots_4_grant ? issue_slots_4_uop_iw_state : _GEN_3533; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_ctrl_op3_sel = slots_4_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3633 = issue_slots_4_grant ? issue_slots_4_uop_ctrl_op3_sel : _GEN_3534; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_ctrl_is_std = slots_4_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3634 = issue_slots_4_grant ? issue_slots_4_uop_ctrl_is_std : _GEN_3535; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_ctrl_is_sta = slots_4_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3635 = issue_slots_4_grant ? issue_slots_4_uop_ctrl_is_sta : _GEN_3536; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_ctrl_is_load = slots_4_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3636 = issue_slots_4_grant ? issue_slots_4_uop_ctrl_is_load : _GEN_3537; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_4_uop_ctrl_csr_cmd = slots_4_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3637 = issue_slots_4_grant ? issue_slots_4_uop_ctrl_csr_cmd : _GEN_3538; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_ctrl_fcn_dw = slots_4_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3638 = issue_slots_4_grant ? issue_slots_4_uop_ctrl_fcn_dw : _GEN_3539; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_4_uop_ctrl_op_fcn = slots_4_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3639 = issue_slots_4_grant ? issue_slots_4_uop_ctrl_op_fcn : _GEN_3540; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_4_uop_ctrl_imm_sel = slots_4_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3640 = issue_slots_4_grant ? issue_slots_4_uop_ctrl_imm_sel : _GEN_3541; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_4_uop_ctrl_op2_sel = slots_4_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3641 = issue_slots_4_grant ? issue_slots_4_uop_ctrl_op2_sel : _GEN_3542; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_ctrl_op1_sel = slots_4_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3642 = issue_slots_4_grant ? issue_slots_4_uop_ctrl_op1_sel : _GEN_3543; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_4_uop_ctrl_br_type = slots_4_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3643 = issue_slots_4_grant ? issue_slots_4_uop_ctrl_br_type : _GEN_3544; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_3644 = issue_slots_4_grant ? issue_slots_4_uop_fu_code : _GEN_3545; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_4_uop_iq_type = slots_4_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3645 = issue_slots_4_grant ? issue_slots_4_uop_iq_type : _GEN_3546; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_4_uop_debug_pc = slots_4_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_3646 = issue_slots_4_grant ? issue_slots_4_uop_debug_pc : _GEN_3547; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_rvc = slots_4_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3647 = issue_slots_4_grant ? issue_slots_4_uop_is_rvc : _GEN_3548; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_4_uop_debug_inst = slots_4_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_3648 = issue_slots_4_grant ? issue_slots_4_uop_debug_inst : _GEN_3549; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_4_uop_inst = slots_4_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_3649 = issue_slots_4_grant ? issue_slots_4_uop_inst : _GEN_3550; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_4_uop_uopc = slots_4_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3650 = issue_slots_4_grant ? issue_slots_4_uop_uopc : _GEN_3551; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_4_uop_address_num = slots_4_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3651 = issue_slots_4_grant ? issue_slots_4_uop_address_num : _GEN_3552; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_4_uop_rob_inst_idx = slots_4_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3652 = issue_slots_4_grant ? issue_slots_4_uop_rob_inst_idx : _GEN_3553; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_4_uop_self_index = slots_4_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3653 = issue_slots_4_grant ? issue_slots_4_uop_self_index : _GEN_3554; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_4_uop_split_num = slots_4_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3654 = issue_slots_4_grant ? issue_slots_4_uop_split_num : _GEN_3555; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_4_uop_op2_sel = slots_4_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3655 = issue_slots_4_grant ? issue_slots_4_uop_op2_sel : _GEN_3556; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_4_uop_op1_sel = slots_4_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3656 = issue_slots_4_grant ? issue_slots_4_uop_op1_sel : _GEN_3557; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_4_uop_stale_pflag = slots_4_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3657 = issue_slots_4_grant ? issue_slots_4_uop_stale_pflag : _GEN_3558; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_pflag_busy = slots_4_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3658 = issue_slots_4_grant ? issue_slots_4_uop_pflag_busy : _GEN_3559; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_4_uop_pwflag = slots_4_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3659 = issue_slots_4_grant ? issue_slots_4_uop_pwflag : _GEN_3560; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_4_uop_prflag = slots_4_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3660 = issue_slots_4_grant ? issue_slots_4_uop_prflag : _GEN_3561; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_wflag = slots_4_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3661 = issue_slots_4_grant ? issue_slots_4_uop_wflag : _GEN_3562; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_rflag = slots_4_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3662 = issue_slots_4_grant ? issue_slots_4_uop_rflag : _GEN_3563; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_4_uop_lrs3_rtype = slots_4_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3663 = issue_slots_4_grant ? issue_slots_4_uop_lrs3_rtype : _GEN_3564; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_4_uop_shift = slots_4_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3664 = issue_slots_4_grant ? issue_slots_4_uop_shift : _GEN_3565; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_is_unicore = slots_4_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3665 = issue_slots_4_grant ? issue_slots_4_uop_is_unicore : _GEN_3566; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_switch_off = slots_4_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3666 = issue_slots_4_grant ? issue_slots_4_uop_switch_off : _GEN_3567; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_4_uop_switch = slots_4_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3667 = issue_slots_4_grant ? issue_slots_4_uop_switch : _GEN_3568; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_debug_tsrc = slots_5_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3670 = issue_slots_5_grant ? issue_slots_5_uop_debug_tsrc : _GEN_3571; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_debug_fsrc = slots_5_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3671 = issue_slots_5_grant ? issue_slots_5_uop_debug_fsrc : _GEN_3572; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_bp_xcpt_if = slots_5_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3672 = issue_slots_5_grant ? issue_slots_5_uop_bp_xcpt_if : _GEN_3573; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_bp_debug_if = slots_5_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3673 = issue_slots_5_grant ? issue_slots_5_uop_bp_debug_if : _GEN_3574; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_xcpt_ma_if = slots_5_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3674 = issue_slots_5_grant ? issue_slots_5_uop_xcpt_ma_if : _GEN_3575; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_xcpt_ae_if = slots_5_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3675 = issue_slots_5_grant ? issue_slots_5_uop_xcpt_ae_if : _GEN_3576; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_xcpt_pf_if = slots_5_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3676 = issue_slots_5_grant ? issue_slots_5_uop_xcpt_pf_if : _GEN_3577; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_fp_single = slots_5_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3677 = issue_slots_5_grant ? issue_slots_5_uop_fp_single : _GEN_3578; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_fp_val = slots_5_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3678 = issue_slots_5_grant ? issue_slots_5_uop_fp_val : _GEN_3579; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_frs3_en = slots_5_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3679 = issue_slots_5_grant ? issue_slots_5_uop_frs3_en : _GEN_3580; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_lrs2_rtype = slots_5_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3680 = issue_slots_5_grant ? issue_slots_5_uop_lrs2_rtype : _GEN_3581; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_lrs1_rtype = slots_5_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3681 = issue_slots_5_grant ? issue_slots_5_uop_lrs1_rtype : _GEN_3582; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_dst_rtype = slots_5_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3682 = issue_slots_5_grant ? issue_slots_5_uop_dst_rtype : _GEN_3583; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_ldst_val = slots_5_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3683 = issue_slots_5_grant ? issue_slots_5_uop_ldst_val : _GEN_3584; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_5_uop_lrs3 = slots_5_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3684 = issue_slots_5_grant ? issue_slots_5_uop_lrs3 : _GEN_3585; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_5_uop_lrs2 = slots_5_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3685 = issue_slots_5_grant ? issue_slots_5_uop_lrs2 : _GEN_3586; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_5_uop_lrs1 = slots_5_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3686 = issue_slots_5_grant ? issue_slots_5_uop_lrs1 : _GEN_3587; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_5_uop_ldst = slots_5_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3687 = issue_slots_5_grant ? issue_slots_5_uop_ldst : _GEN_3588; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_ldst_is_rs1 = slots_5_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3688 = issue_slots_5_grant ? issue_slots_5_uop_ldst_is_rs1 : _GEN_3589; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_flush_on_commit = slots_5_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3689 = issue_slots_5_grant ? issue_slots_5_uop_flush_on_commit : _GEN_3590; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_unique = slots_5_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3690 = issue_slots_5_grant ? issue_slots_5_uop_is_unique : _GEN_3591; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_sys_pc2epc = slots_5_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3691 = issue_slots_5_grant ? issue_slots_5_uop_is_sys_pc2epc : _GEN_3592; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_uses_stq = slots_5_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3692 = issue_slots_5_grant ? issue_slots_5_uop_uses_stq : _GEN_3593; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_uses_ldq = slots_5_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3693 = issue_slots_5_grant ? issue_slots_5_uop_uses_ldq : _GEN_3594; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_amo = slots_5_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3694 = issue_slots_5_grant ? issue_slots_5_uop_is_amo : _GEN_3595; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_fencei = slots_5_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3695 = issue_slots_5_grant ? issue_slots_5_uop_is_fencei : _GEN_3596; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_fence = slots_5_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3696 = issue_slots_5_grant ? issue_slots_5_uop_is_fence : _GEN_3597; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_mem_signed = slots_5_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3697 = issue_slots_5_grant ? issue_slots_5_uop_mem_signed : _GEN_3598; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_mem_size = slots_5_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3698 = issue_slots_5_grant ? issue_slots_5_uop_mem_size : _GEN_3599; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_5_uop_mem_cmd = slots_5_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3699 = issue_slots_5_grant ? issue_slots_5_uop_mem_cmd : _GEN_3600; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_bypassable = slots_5_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3700 = issue_slots_5_grant ? issue_slots_5_uop_bypassable : _GEN_3601; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_5_uop_exc_cause = slots_5_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_3701 = issue_slots_5_grant ? issue_slots_5_uop_exc_cause : _GEN_3602; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_exception = slots_5_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3702 = issue_slots_5_grant ? issue_slots_5_uop_exception : _GEN_3603; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_5_uop_stale_pdst = slots_5_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3703 = issue_slots_5_grant ? issue_slots_5_uop_stale_pdst : _GEN_3604; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_ppred_busy = slots_5_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3704 = issue_slots_5_grant ? issue_slots_5_uop_ppred_busy : _GEN_3605; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_prs3_busy = slots_5_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3705 = issue_slots_5_grant ? issue_slots_5_uop_prs3_busy : _GEN_3606; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_prs2_busy = slots_5_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3706 = issue_slots_5_grant ? issue_slots_5_uop_prs2_busy : _GEN_3607; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_prs1_busy = slots_5_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3707 = issue_slots_5_grant ? issue_slots_5_uop_prs1_busy : _GEN_3608; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_5_uop_ppred = slots_5_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3708 = issue_slots_5_grant ? issue_slots_5_uop_ppred : _GEN_3609; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_5_uop_prs3 = slots_5_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3709 = issue_slots_5_grant ? issue_slots_5_uop_prs3 : _GEN_3610; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_5_uop_prs2 = slots_5_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3710 = issue_slots_5_grant ? issue_slots_5_uop_prs2 : _GEN_3611; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_5_uop_prs1 = slots_5_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3711 = issue_slots_5_grant ? issue_slots_5_uop_prs1 : _GEN_3612; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_5_uop_pdst = slots_5_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3712 = issue_slots_5_grant ? issue_slots_5_uop_pdst : _GEN_3613; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_rxq_idx = slots_5_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3713 = issue_slots_5_grant ? issue_slots_5_uop_rxq_idx : _GEN_3614; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_5_uop_stq_idx = slots_5_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3714 = issue_slots_5_grant ? issue_slots_5_uop_stq_idx : _GEN_3615; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_5_uop_ldq_idx = slots_5_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3715 = issue_slots_5_grant ? issue_slots_5_uop_ldq_idx : _GEN_3616; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_5_uop_rob_idx = slots_5_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3716 = issue_slots_5_grant ? issue_slots_5_uop_rob_idx : _GEN_3617; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_5_uop_csr_addr = slots_5_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_3717 = issue_slots_5_grant ? issue_slots_5_uop_csr_addr : _GEN_3618; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_5_uop_imm_packed = slots_5_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_3718 = issue_slots_5_grant ? issue_slots_5_uop_imm_packed : _GEN_3619; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_taken = slots_5_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3719 = issue_slots_5_grant ? issue_slots_5_uop_taken : _GEN_3620; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_5_uop_pc_lob = slots_5_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3720 = issue_slots_5_grant ? issue_slots_5_uop_pc_lob : _GEN_3621; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_edge_inst = slots_5_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3721 = issue_slots_5_grant ? issue_slots_5_uop_edge_inst : _GEN_3622; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_5_uop_ftq_idx = slots_5_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3722 = issue_slots_5_grant ? issue_slots_5_uop_ftq_idx : _GEN_3623; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_5_uop_br_tag = slots_5_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3723 = issue_slots_5_grant ? issue_slots_5_uop_br_tag : _GEN_3624; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_5_uop_br_mask = slots_5_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_3724 = issue_slots_5_grant ? issue_slots_5_uop_br_mask : _GEN_3625; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_sfb = slots_5_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3725 = issue_slots_5_grant ? issue_slots_5_uop_is_sfb : _GEN_3626; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_jal = slots_5_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3726 = issue_slots_5_grant ? issue_slots_5_uop_is_jal : _GEN_3627; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_jalr = slots_5_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3727 = issue_slots_5_grant ? issue_slots_5_uop_is_jalr : _GEN_3628; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_br = slots_5_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3728 = issue_slots_5_grant ? issue_slots_5_uop_is_br : _GEN_3629; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_iw_p2_poisoned = slots_5_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3729 = issue_slots_5_grant ? issue_slots_5_uop_iw_p2_poisoned : _GEN_3630; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_iw_p1_poisoned = slots_5_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3730 = issue_slots_5_grant ? issue_slots_5_uop_iw_p1_poisoned : _GEN_3631; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_iw_state = slots_5_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3731 = issue_slots_5_grant ? issue_slots_5_uop_iw_state : _GEN_3632; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_ctrl_op3_sel = slots_5_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3732 = issue_slots_5_grant ? issue_slots_5_uop_ctrl_op3_sel : _GEN_3633; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_ctrl_is_std = slots_5_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3733 = issue_slots_5_grant ? issue_slots_5_uop_ctrl_is_std : _GEN_3634; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_ctrl_is_sta = slots_5_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3734 = issue_slots_5_grant ? issue_slots_5_uop_ctrl_is_sta : _GEN_3635; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_ctrl_is_load = slots_5_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3735 = issue_slots_5_grant ? issue_slots_5_uop_ctrl_is_load : _GEN_3636; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_5_uop_ctrl_csr_cmd = slots_5_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3736 = issue_slots_5_grant ? issue_slots_5_uop_ctrl_csr_cmd : _GEN_3637; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_ctrl_fcn_dw = slots_5_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3737 = issue_slots_5_grant ? issue_slots_5_uop_ctrl_fcn_dw : _GEN_3638; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_5_uop_ctrl_op_fcn = slots_5_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3738 = issue_slots_5_grant ? issue_slots_5_uop_ctrl_op_fcn : _GEN_3639; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_5_uop_ctrl_imm_sel = slots_5_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3739 = issue_slots_5_grant ? issue_slots_5_uop_ctrl_imm_sel : _GEN_3640; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_5_uop_ctrl_op2_sel = slots_5_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3740 = issue_slots_5_grant ? issue_slots_5_uop_ctrl_op2_sel : _GEN_3641; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_ctrl_op1_sel = slots_5_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3741 = issue_slots_5_grant ? issue_slots_5_uop_ctrl_op1_sel : _GEN_3642; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_5_uop_ctrl_br_type = slots_5_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3742 = issue_slots_5_grant ? issue_slots_5_uop_ctrl_br_type : _GEN_3643; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_3743 = issue_slots_5_grant ? issue_slots_5_uop_fu_code : _GEN_3644; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_5_uop_iq_type = slots_5_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3744 = issue_slots_5_grant ? issue_slots_5_uop_iq_type : _GEN_3645; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_5_uop_debug_pc = slots_5_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_3745 = issue_slots_5_grant ? issue_slots_5_uop_debug_pc : _GEN_3646; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_rvc = slots_5_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3746 = issue_slots_5_grant ? issue_slots_5_uop_is_rvc : _GEN_3647; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_5_uop_debug_inst = slots_5_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_3747 = issue_slots_5_grant ? issue_slots_5_uop_debug_inst : _GEN_3648; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_5_uop_inst = slots_5_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_3748 = issue_slots_5_grant ? issue_slots_5_uop_inst : _GEN_3649; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_5_uop_uopc = slots_5_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3749 = issue_slots_5_grant ? issue_slots_5_uop_uopc : _GEN_3650; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_5_uop_address_num = slots_5_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3750 = issue_slots_5_grant ? issue_slots_5_uop_address_num : _GEN_3651; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_5_uop_rob_inst_idx = slots_5_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3751 = issue_slots_5_grant ? issue_slots_5_uop_rob_inst_idx : _GEN_3652; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_5_uop_self_index = slots_5_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3752 = issue_slots_5_grant ? issue_slots_5_uop_self_index : _GEN_3653; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_5_uop_split_num = slots_5_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3753 = issue_slots_5_grant ? issue_slots_5_uop_split_num : _GEN_3654; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_5_uop_op2_sel = slots_5_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3754 = issue_slots_5_grant ? issue_slots_5_uop_op2_sel : _GEN_3655; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_5_uop_op1_sel = slots_5_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3755 = issue_slots_5_grant ? issue_slots_5_uop_op1_sel : _GEN_3656; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_5_uop_stale_pflag = slots_5_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3756 = issue_slots_5_grant ? issue_slots_5_uop_stale_pflag : _GEN_3657; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_pflag_busy = slots_5_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3757 = issue_slots_5_grant ? issue_slots_5_uop_pflag_busy : _GEN_3658; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_5_uop_pwflag = slots_5_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3758 = issue_slots_5_grant ? issue_slots_5_uop_pwflag : _GEN_3659; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_5_uop_prflag = slots_5_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3759 = issue_slots_5_grant ? issue_slots_5_uop_prflag : _GEN_3660; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_wflag = slots_5_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3760 = issue_slots_5_grant ? issue_slots_5_uop_wflag : _GEN_3661; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_rflag = slots_5_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3761 = issue_slots_5_grant ? issue_slots_5_uop_rflag : _GEN_3662; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_5_uop_lrs3_rtype = slots_5_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3762 = issue_slots_5_grant ? issue_slots_5_uop_lrs3_rtype : _GEN_3663; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_5_uop_shift = slots_5_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3763 = issue_slots_5_grant ? issue_slots_5_uop_shift : _GEN_3664; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_is_unicore = slots_5_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3764 = issue_slots_5_grant ? issue_slots_5_uop_is_unicore : _GEN_3665; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_switch_off = slots_5_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3765 = issue_slots_5_grant ? issue_slots_5_uop_switch_off : _GEN_3666; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_5_uop_switch = slots_5_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3766 = issue_slots_5_grant ? issue_slots_5_uop_switch : _GEN_3667; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_debug_tsrc = slots_6_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3769 = issue_slots_6_grant ? issue_slots_6_uop_debug_tsrc : _GEN_3670; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_debug_fsrc = slots_6_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3770 = issue_slots_6_grant ? issue_slots_6_uop_debug_fsrc : _GEN_3671; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_bp_xcpt_if = slots_6_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3771 = issue_slots_6_grant ? issue_slots_6_uop_bp_xcpt_if : _GEN_3672; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_bp_debug_if = slots_6_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3772 = issue_slots_6_grant ? issue_slots_6_uop_bp_debug_if : _GEN_3673; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_xcpt_ma_if = slots_6_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3773 = issue_slots_6_grant ? issue_slots_6_uop_xcpt_ma_if : _GEN_3674; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_xcpt_ae_if = slots_6_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3774 = issue_slots_6_grant ? issue_slots_6_uop_xcpt_ae_if : _GEN_3675; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_xcpt_pf_if = slots_6_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3775 = issue_slots_6_grant ? issue_slots_6_uop_xcpt_pf_if : _GEN_3676; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_fp_single = slots_6_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3776 = issue_slots_6_grant ? issue_slots_6_uop_fp_single : _GEN_3677; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_fp_val = slots_6_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3777 = issue_slots_6_grant ? issue_slots_6_uop_fp_val : _GEN_3678; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_frs3_en = slots_6_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3778 = issue_slots_6_grant ? issue_slots_6_uop_frs3_en : _GEN_3679; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_lrs2_rtype = slots_6_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3779 = issue_slots_6_grant ? issue_slots_6_uop_lrs2_rtype : _GEN_3680; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_lrs1_rtype = slots_6_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3780 = issue_slots_6_grant ? issue_slots_6_uop_lrs1_rtype : _GEN_3681; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_dst_rtype = slots_6_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3781 = issue_slots_6_grant ? issue_slots_6_uop_dst_rtype : _GEN_3682; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_ldst_val = slots_6_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3782 = issue_slots_6_grant ? issue_slots_6_uop_ldst_val : _GEN_3683; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_6_uop_lrs3 = slots_6_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3783 = issue_slots_6_grant ? issue_slots_6_uop_lrs3 : _GEN_3684; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_6_uop_lrs2 = slots_6_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3784 = issue_slots_6_grant ? issue_slots_6_uop_lrs2 : _GEN_3685; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_6_uop_lrs1 = slots_6_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3785 = issue_slots_6_grant ? issue_slots_6_uop_lrs1 : _GEN_3686; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_6_uop_ldst = slots_6_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3786 = issue_slots_6_grant ? issue_slots_6_uop_ldst : _GEN_3687; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_ldst_is_rs1 = slots_6_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3787 = issue_slots_6_grant ? issue_slots_6_uop_ldst_is_rs1 : _GEN_3688; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_flush_on_commit = slots_6_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3788 = issue_slots_6_grant ? issue_slots_6_uop_flush_on_commit : _GEN_3689; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_unique = slots_6_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3789 = issue_slots_6_grant ? issue_slots_6_uop_is_unique : _GEN_3690; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_sys_pc2epc = slots_6_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3790 = issue_slots_6_grant ? issue_slots_6_uop_is_sys_pc2epc : _GEN_3691; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_uses_stq = slots_6_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3791 = issue_slots_6_grant ? issue_slots_6_uop_uses_stq : _GEN_3692; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_uses_ldq = slots_6_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3792 = issue_slots_6_grant ? issue_slots_6_uop_uses_ldq : _GEN_3693; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_amo = slots_6_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3793 = issue_slots_6_grant ? issue_slots_6_uop_is_amo : _GEN_3694; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_fencei = slots_6_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3794 = issue_slots_6_grant ? issue_slots_6_uop_is_fencei : _GEN_3695; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_fence = slots_6_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3795 = issue_slots_6_grant ? issue_slots_6_uop_is_fence : _GEN_3696; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_mem_signed = slots_6_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3796 = issue_slots_6_grant ? issue_slots_6_uop_mem_signed : _GEN_3697; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_mem_size = slots_6_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3797 = issue_slots_6_grant ? issue_slots_6_uop_mem_size : _GEN_3698; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_6_uop_mem_cmd = slots_6_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3798 = issue_slots_6_grant ? issue_slots_6_uop_mem_cmd : _GEN_3699; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_bypassable = slots_6_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3799 = issue_slots_6_grant ? issue_slots_6_uop_bypassable : _GEN_3700; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_6_uop_exc_cause = slots_6_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_3800 = issue_slots_6_grant ? issue_slots_6_uop_exc_cause : _GEN_3701; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_exception = slots_6_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3801 = issue_slots_6_grant ? issue_slots_6_uop_exception : _GEN_3702; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_6_uop_stale_pdst = slots_6_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3802 = issue_slots_6_grant ? issue_slots_6_uop_stale_pdst : _GEN_3703; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_ppred_busy = slots_6_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3803 = issue_slots_6_grant ? issue_slots_6_uop_ppred_busy : _GEN_3704; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_prs3_busy = slots_6_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3804 = issue_slots_6_grant ? issue_slots_6_uop_prs3_busy : _GEN_3705; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_prs2_busy = slots_6_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3805 = issue_slots_6_grant ? issue_slots_6_uop_prs2_busy : _GEN_3706; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_prs1_busy = slots_6_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3806 = issue_slots_6_grant ? issue_slots_6_uop_prs1_busy : _GEN_3707; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_6_uop_ppred = slots_6_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3807 = issue_slots_6_grant ? issue_slots_6_uop_ppred : _GEN_3708; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_6_uop_prs3 = slots_6_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3808 = issue_slots_6_grant ? issue_slots_6_uop_prs3 : _GEN_3709; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_6_uop_prs2 = slots_6_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3809 = issue_slots_6_grant ? issue_slots_6_uop_prs2 : _GEN_3710; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_6_uop_prs1 = slots_6_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3810 = issue_slots_6_grant ? issue_slots_6_uop_prs1 : _GEN_3711; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_6_uop_pdst = slots_6_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3811 = issue_slots_6_grant ? issue_slots_6_uop_pdst : _GEN_3712; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_rxq_idx = slots_6_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3812 = issue_slots_6_grant ? issue_slots_6_uop_rxq_idx : _GEN_3713; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_6_uop_stq_idx = slots_6_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3813 = issue_slots_6_grant ? issue_slots_6_uop_stq_idx : _GEN_3714; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_6_uop_ldq_idx = slots_6_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3814 = issue_slots_6_grant ? issue_slots_6_uop_ldq_idx : _GEN_3715; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_6_uop_rob_idx = slots_6_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3815 = issue_slots_6_grant ? issue_slots_6_uop_rob_idx : _GEN_3716; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_6_uop_csr_addr = slots_6_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_3816 = issue_slots_6_grant ? issue_slots_6_uop_csr_addr : _GEN_3717; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_6_uop_imm_packed = slots_6_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_3817 = issue_slots_6_grant ? issue_slots_6_uop_imm_packed : _GEN_3718; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_taken = slots_6_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3818 = issue_slots_6_grant ? issue_slots_6_uop_taken : _GEN_3719; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_6_uop_pc_lob = slots_6_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3819 = issue_slots_6_grant ? issue_slots_6_uop_pc_lob : _GEN_3720; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_edge_inst = slots_6_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3820 = issue_slots_6_grant ? issue_slots_6_uop_edge_inst : _GEN_3721; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_6_uop_ftq_idx = slots_6_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3821 = issue_slots_6_grant ? issue_slots_6_uop_ftq_idx : _GEN_3722; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_6_uop_br_tag = slots_6_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3822 = issue_slots_6_grant ? issue_slots_6_uop_br_tag : _GEN_3723; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_6_uop_br_mask = slots_6_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_3823 = issue_slots_6_grant ? issue_slots_6_uop_br_mask : _GEN_3724; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_sfb = slots_6_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3824 = issue_slots_6_grant ? issue_slots_6_uop_is_sfb : _GEN_3725; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_jal = slots_6_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3825 = issue_slots_6_grant ? issue_slots_6_uop_is_jal : _GEN_3726; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_jalr = slots_6_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3826 = issue_slots_6_grant ? issue_slots_6_uop_is_jalr : _GEN_3727; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_br = slots_6_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3827 = issue_slots_6_grant ? issue_slots_6_uop_is_br : _GEN_3728; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_iw_p2_poisoned = slots_6_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3828 = issue_slots_6_grant ? issue_slots_6_uop_iw_p2_poisoned : _GEN_3729; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_iw_p1_poisoned = slots_6_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3829 = issue_slots_6_grant ? issue_slots_6_uop_iw_p1_poisoned : _GEN_3730; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_iw_state = slots_6_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3830 = issue_slots_6_grant ? issue_slots_6_uop_iw_state : _GEN_3731; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_ctrl_op3_sel = slots_6_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3831 = issue_slots_6_grant ? issue_slots_6_uop_ctrl_op3_sel : _GEN_3732; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_ctrl_is_std = slots_6_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3832 = issue_slots_6_grant ? issue_slots_6_uop_ctrl_is_std : _GEN_3733; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_ctrl_is_sta = slots_6_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3833 = issue_slots_6_grant ? issue_slots_6_uop_ctrl_is_sta : _GEN_3734; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_ctrl_is_load = slots_6_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3834 = issue_slots_6_grant ? issue_slots_6_uop_ctrl_is_load : _GEN_3735; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_6_uop_ctrl_csr_cmd = slots_6_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3835 = issue_slots_6_grant ? issue_slots_6_uop_ctrl_csr_cmd : _GEN_3736; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_ctrl_fcn_dw = slots_6_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3836 = issue_slots_6_grant ? issue_slots_6_uop_ctrl_fcn_dw : _GEN_3737; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_6_uop_ctrl_op_fcn = slots_6_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3837 = issue_slots_6_grant ? issue_slots_6_uop_ctrl_op_fcn : _GEN_3738; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_6_uop_ctrl_imm_sel = slots_6_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3838 = issue_slots_6_grant ? issue_slots_6_uop_ctrl_imm_sel : _GEN_3739; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_6_uop_ctrl_op2_sel = slots_6_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3839 = issue_slots_6_grant ? issue_slots_6_uop_ctrl_op2_sel : _GEN_3740; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_ctrl_op1_sel = slots_6_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3840 = issue_slots_6_grant ? issue_slots_6_uop_ctrl_op1_sel : _GEN_3741; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_6_uop_ctrl_br_type = slots_6_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3841 = issue_slots_6_grant ? issue_slots_6_uop_ctrl_br_type : _GEN_3742; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_3842 = issue_slots_6_grant ? issue_slots_6_uop_fu_code : _GEN_3743; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_6_uop_iq_type = slots_6_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3843 = issue_slots_6_grant ? issue_slots_6_uop_iq_type : _GEN_3744; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_6_uop_debug_pc = slots_6_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_3844 = issue_slots_6_grant ? issue_slots_6_uop_debug_pc : _GEN_3745; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_rvc = slots_6_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3845 = issue_slots_6_grant ? issue_slots_6_uop_is_rvc : _GEN_3746; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_6_uop_debug_inst = slots_6_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_3846 = issue_slots_6_grant ? issue_slots_6_uop_debug_inst : _GEN_3747; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_6_uop_inst = slots_6_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_3847 = issue_slots_6_grant ? issue_slots_6_uop_inst : _GEN_3748; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_6_uop_uopc = slots_6_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3848 = issue_slots_6_grant ? issue_slots_6_uop_uopc : _GEN_3749; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_6_uop_address_num = slots_6_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3849 = issue_slots_6_grant ? issue_slots_6_uop_address_num : _GEN_3750; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_6_uop_rob_inst_idx = slots_6_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3850 = issue_slots_6_grant ? issue_slots_6_uop_rob_inst_idx : _GEN_3751; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_6_uop_self_index = slots_6_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3851 = issue_slots_6_grant ? issue_slots_6_uop_self_index : _GEN_3752; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_6_uop_split_num = slots_6_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3852 = issue_slots_6_grant ? issue_slots_6_uop_split_num : _GEN_3753; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_6_uop_op2_sel = slots_6_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3853 = issue_slots_6_grant ? issue_slots_6_uop_op2_sel : _GEN_3754; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_6_uop_op1_sel = slots_6_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3854 = issue_slots_6_grant ? issue_slots_6_uop_op1_sel : _GEN_3755; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_6_uop_stale_pflag = slots_6_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3855 = issue_slots_6_grant ? issue_slots_6_uop_stale_pflag : _GEN_3756; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_pflag_busy = slots_6_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3856 = issue_slots_6_grant ? issue_slots_6_uop_pflag_busy : _GEN_3757; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_6_uop_pwflag = slots_6_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3857 = issue_slots_6_grant ? issue_slots_6_uop_pwflag : _GEN_3758; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_6_uop_prflag = slots_6_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3858 = issue_slots_6_grant ? issue_slots_6_uop_prflag : _GEN_3759; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_wflag = slots_6_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3859 = issue_slots_6_grant ? issue_slots_6_uop_wflag : _GEN_3760; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_rflag = slots_6_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3860 = issue_slots_6_grant ? issue_slots_6_uop_rflag : _GEN_3761; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_6_uop_lrs3_rtype = slots_6_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3861 = issue_slots_6_grant ? issue_slots_6_uop_lrs3_rtype : _GEN_3762; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_6_uop_shift = slots_6_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3862 = issue_slots_6_grant ? issue_slots_6_uop_shift : _GEN_3763; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_is_unicore = slots_6_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3863 = issue_slots_6_grant ? issue_slots_6_uop_is_unicore : _GEN_3764; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_switch_off = slots_6_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3864 = issue_slots_6_grant ? issue_slots_6_uop_switch_off : _GEN_3765; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_6_uop_switch = slots_6_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3865 = issue_slots_6_grant ? issue_slots_6_uop_switch : _GEN_3766; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_debug_tsrc = slots_7_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3868 = issue_slots_7_grant ? issue_slots_7_uop_debug_tsrc : _GEN_3769; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_debug_fsrc = slots_7_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3869 = issue_slots_7_grant ? issue_slots_7_uop_debug_fsrc : _GEN_3770; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_bp_xcpt_if = slots_7_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3870 = issue_slots_7_grant ? issue_slots_7_uop_bp_xcpt_if : _GEN_3771; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_bp_debug_if = slots_7_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3871 = issue_slots_7_grant ? issue_slots_7_uop_bp_debug_if : _GEN_3772; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_xcpt_ma_if = slots_7_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3872 = issue_slots_7_grant ? issue_slots_7_uop_xcpt_ma_if : _GEN_3773; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_xcpt_ae_if = slots_7_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3873 = issue_slots_7_grant ? issue_slots_7_uop_xcpt_ae_if : _GEN_3774; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_xcpt_pf_if = slots_7_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3874 = issue_slots_7_grant ? issue_slots_7_uop_xcpt_pf_if : _GEN_3775; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_fp_single = slots_7_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3875 = issue_slots_7_grant ? issue_slots_7_uop_fp_single : _GEN_3776; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_fp_val = slots_7_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3876 = issue_slots_7_grant ? issue_slots_7_uop_fp_val : _GEN_3777; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_frs3_en = slots_7_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3877 = issue_slots_7_grant ? issue_slots_7_uop_frs3_en : _GEN_3778; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_lrs2_rtype = slots_7_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3878 = issue_slots_7_grant ? issue_slots_7_uop_lrs2_rtype : _GEN_3779; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_lrs1_rtype = slots_7_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3879 = issue_slots_7_grant ? issue_slots_7_uop_lrs1_rtype : _GEN_3780; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_dst_rtype = slots_7_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3880 = issue_slots_7_grant ? issue_slots_7_uop_dst_rtype : _GEN_3781; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_ldst_val = slots_7_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3881 = issue_slots_7_grant ? issue_slots_7_uop_ldst_val : _GEN_3782; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_7_uop_lrs3 = slots_7_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3882 = issue_slots_7_grant ? issue_slots_7_uop_lrs3 : _GEN_3783; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_7_uop_lrs2 = slots_7_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3883 = issue_slots_7_grant ? issue_slots_7_uop_lrs2 : _GEN_3784; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_7_uop_lrs1 = slots_7_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3884 = issue_slots_7_grant ? issue_slots_7_uop_lrs1 : _GEN_3785; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_7_uop_ldst = slots_7_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3885 = issue_slots_7_grant ? issue_slots_7_uop_ldst : _GEN_3786; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_ldst_is_rs1 = slots_7_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3886 = issue_slots_7_grant ? issue_slots_7_uop_ldst_is_rs1 : _GEN_3787; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_flush_on_commit = slots_7_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3887 = issue_slots_7_grant ? issue_slots_7_uop_flush_on_commit : _GEN_3788; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_unique = slots_7_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3888 = issue_slots_7_grant ? issue_slots_7_uop_is_unique : _GEN_3789; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_sys_pc2epc = slots_7_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3889 = issue_slots_7_grant ? issue_slots_7_uop_is_sys_pc2epc : _GEN_3790; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_uses_stq = slots_7_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3890 = issue_slots_7_grant ? issue_slots_7_uop_uses_stq : _GEN_3791; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_uses_ldq = slots_7_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3891 = issue_slots_7_grant ? issue_slots_7_uop_uses_ldq : _GEN_3792; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_amo = slots_7_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3892 = issue_slots_7_grant ? issue_slots_7_uop_is_amo : _GEN_3793; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_fencei = slots_7_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3893 = issue_slots_7_grant ? issue_slots_7_uop_is_fencei : _GEN_3794; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_fence = slots_7_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3894 = issue_slots_7_grant ? issue_slots_7_uop_is_fence : _GEN_3795; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_mem_signed = slots_7_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3895 = issue_slots_7_grant ? issue_slots_7_uop_mem_signed : _GEN_3796; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_mem_size = slots_7_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3896 = issue_slots_7_grant ? issue_slots_7_uop_mem_size : _GEN_3797; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_7_uop_mem_cmd = slots_7_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3897 = issue_slots_7_grant ? issue_slots_7_uop_mem_cmd : _GEN_3798; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_bypassable = slots_7_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3898 = issue_slots_7_grant ? issue_slots_7_uop_bypassable : _GEN_3799; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_7_uop_exc_cause = slots_7_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_3899 = issue_slots_7_grant ? issue_slots_7_uop_exc_cause : _GEN_3800; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_exception = slots_7_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3900 = issue_slots_7_grant ? issue_slots_7_uop_exception : _GEN_3801; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_7_uop_stale_pdst = slots_7_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3901 = issue_slots_7_grant ? issue_slots_7_uop_stale_pdst : _GEN_3802; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_ppred_busy = slots_7_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3902 = issue_slots_7_grant ? issue_slots_7_uop_ppred_busy : _GEN_3803; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_prs3_busy = slots_7_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3903 = issue_slots_7_grant ? issue_slots_7_uop_prs3_busy : _GEN_3804; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_prs2_busy = slots_7_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3904 = issue_slots_7_grant ? issue_slots_7_uop_prs2_busy : _GEN_3805; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_prs1_busy = slots_7_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3905 = issue_slots_7_grant ? issue_slots_7_uop_prs1_busy : _GEN_3806; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_7_uop_ppred = slots_7_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3906 = issue_slots_7_grant ? issue_slots_7_uop_ppred : _GEN_3807; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_7_uop_prs3 = slots_7_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3907 = issue_slots_7_grant ? issue_slots_7_uop_prs3 : _GEN_3808; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_7_uop_prs2 = slots_7_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3908 = issue_slots_7_grant ? issue_slots_7_uop_prs2 : _GEN_3809; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_7_uop_prs1 = slots_7_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3909 = issue_slots_7_grant ? issue_slots_7_uop_prs1 : _GEN_3810; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_7_uop_pdst = slots_7_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3910 = issue_slots_7_grant ? issue_slots_7_uop_pdst : _GEN_3811; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_rxq_idx = slots_7_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3911 = issue_slots_7_grant ? issue_slots_7_uop_rxq_idx : _GEN_3812; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_7_uop_stq_idx = slots_7_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3912 = issue_slots_7_grant ? issue_slots_7_uop_stq_idx : _GEN_3813; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_7_uop_ldq_idx = slots_7_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3913 = issue_slots_7_grant ? issue_slots_7_uop_ldq_idx : _GEN_3814; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_7_uop_rob_idx = slots_7_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3914 = issue_slots_7_grant ? issue_slots_7_uop_rob_idx : _GEN_3815; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_7_uop_csr_addr = slots_7_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_3915 = issue_slots_7_grant ? issue_slots_7_uop_csr_addr : _GEN_3816; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_7_uop_imm_packed = slots_7_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_3916 = issue_slots_7_grant ? issue_slots_7_uop_imm_packed : _GEN_3817; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_taken = slots_7_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3917 = issue_slots_7_grant ? issue_slots_7_uop_taken : _GEN_3818; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_7_uop_pc_lob = slots_7_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3918 = issue_slots_7_grant ? issue_slots_7_uop_pc_lob : _GEN_3819; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_edge_inst = slots_7_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3919 = issue_slots_7_grant ? issue_slots_7_uop_edge_inst : _GEN_3820; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_7_uop_ftq_idx = slots_7_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3920 = issue_slots_7_grant ? issue_slots_7_uop_ftq_idx : _GEN_3821; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_7_uop_br_tag = slots_7_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3921 = issue_slots_7_grant ? issue_slots_7_uop_br_tag : _GEN_3822; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_7_uop_br_mask = slots_7_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_3922 = issue_slots_7_grant ? issue_slots_7_uop_br_mask : _GEN_3823; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_sfb = slots_7_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3923 = issue_slots_7_grant ? issue_slots_7_uop_is_sfb : _GEN_3824; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_jal = slots_7_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3924 = issue_slots_7_grant ? issue_slots_7_uop_is_jal : _GEN_3825; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_jalr = slots_7_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3925 = issue_slots_7_grant ? issue_slots_7_uop_is_jalr : _GEN_3826; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_br = slots_7_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3926 = issue_slots_7_grant ? issue_slots_7_uop_is_br : _GEN_3827; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_iw_p2_poisoned = slots_7_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3927 = issue_slots_7_grant ? issue_slots_7_uop_iw_p2_poisoned : _GEN_3828; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_iw_p1_poisoned = slots_7_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3928 = issue_slots_7_grant ? issue_slots_7_uop_iw_p1_poisoned : _GEN_3829; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_iw_state = slots_7_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3929 = issue_slots_7_grant ? issue_slots_7_uop_iw_state : _GEN_3830; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_ctrl_op3_sel = slots_7_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3930 = issue_slots_7_grant ? issue_slots_7_uop_ctrl_op3_sel : _GEN_3831; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_ctrl_is_std = slots_7_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3931 = issue_slots_7_grant ? issue_slots_7_uop_ctrl_is_std : _GEN_3832; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_ctrl_is_sta = slots_7_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3932 = issue_slots_7_grant ? issue_slots_7_uop_ctrl_is_sta : _GEN_3833; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_ctrl_is_load = slots_7_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3933 = issue_slots_7_grant ? issue_slots_7_uop_ctrl_is_load : _GEN_3834; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_7_uop_ctrl_csr_cmd = slots_7_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3934 = issue_slots_7_grant ? issue_slots_7_uop_ctrl_csr_cmd : _GEN_3835; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_ctrl_fcn_dw = slots_7_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3935 = issue_slots_7_grant ? issue_slots_7_uop_ctrl_fcn_dw : _GEN_3836; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_7_uop_ctrl_op_fcn = slots_7_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3936 = issue_slots_7_grant ? issue_slots_7_uop_ctrl_op_fcn : _GEN_3837; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_7_uop_ctrl_imm_sel = slots_7_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3937 = issue_slots_7_grant ? issue_slots_7_uop_ctrl_imm_sel : _GEN_3838; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_7_uop_ctrl_op2_sel = slots_7_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3938 = issue_slots_7_grant ? issue_slots_7_uop_ctrl_op2_sel : _GEN_3839; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_ctrl_op1_sel = slots_7_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3939 = issue_slots_7_grant ? issue_slots_7_uop_ctrl_op1_sel : _GEN_3840; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_7_uop_ctrl_br_type = slots_7_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3940 = issue_slots_7_grant ? issue_slots_7_uop_ctrl_br_type : _GEN_3841; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_3941 = issue_slots_7_grant ? issue_slots_7_uop_fu_code : _GEN_3842; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_7_uop_iq_type = slots_7_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3942 = issue_slots_7_grant ? issue_slots_7_uop_iq_type : _GEN_3843; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_7_uop_debug_pc = slots_7_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_3943 = issue_slots_7_grant ? issue_slots_7_uop_debug_pc : _GEN_3844; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_rvc = slots_7_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3944 = issue_slots_7_grant ? issue_slots_7_uop_is_rvc : _GEN_3845; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_7_uop_debug_inst = slots_7_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_3945 = issue_slots_7_grant ? issue_slots_7_uop_debug_inst : _GEN_3846; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_7_uop_inst = slots_7_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_3946 = issue_slots_7_grant ? issue_slots_7_uop_inst : _GEN_3847; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_7_uop_uopc = slots_7_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_3947 = issue_slots_7_grant ? issue_slots_7_uop_uopc : _GEN_3848; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_7_uop_address_num = slots_7_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3948 = issue_slots_7_grant ? issue_slots_7_uop_address_num : _GEN_3849; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_7_uop_rob_inst_idx = slots_7_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3949 = issue_slots_7_grant ? issue_slots_7_uop_rob_inst_idx : _GEN_3850; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_7_uop_self_index = slots_7_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3950 = issue_slots_7_grant ? issue_slots_7_uop_self_index : _GEN_3851; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_7_uop_split_num = slots_7_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3951 = issue_slots_7_grant ? issue_slots_7_uop_split_num : _GEN_3852; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_7_uop_op2_sel = slots_7_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3952 = issue_slots_7_grant ? issue_slots_7_uop_op2_sel : _GEN_3853; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_7_uop_op1_sel = slots_7_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3953 = issue_slots_7_grant ? issue_slots_7_uop_op1_sel : _GEN_3854; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_7_uop_stale_pflag = slots_7_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3954 = issue_slots_7_grant ? issue_slots_7_uop_stale_pflag : _GEN_3855; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_pflag_busy = slots_7_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3955 = issue_slots_7_grant ? issue_slots_7_uop_pflag_busy : _GEN_3856; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_7_uop_pwflag = slots_7_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3956 = issue_slots_7_grant ? issue_slots_7_uop_pwflag : _GEN_3857; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_7_uop_prflag = slots_7_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_3957 = issue_slots_7_grant ? issue_slots_7_uop_prflag : _GEN_3858; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_wflag = slots_7_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3958 = issue_slots_7_grant ? issue_slots_7_uop_wflag : _GEN_3859; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_rflag = slots_7_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3959 = issue_slots_7_grant ? issue_slots_7_uop_rflag : _GEN_3860; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_7_uop_lrs3_rtype = slots_7_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3960 = issue_slots_7_grant ? issue_slots_7_uop_lrs3_rtype : _GEN_3861; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_7_uop_shift = slots_7_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_3961 = issue_slots_7_grant ? issue_slots_7_uop_shift : _GEN_3862; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_is_unicore = slots_7_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3962 = issue_slots_7_grant ? issue_slots_7_uop_is_unicore : _GEN_3863; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_switch_off = slots_7_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3963 = issue_slots_7_grant ? issue_slots_7_uop_switch_off : _GEN_3864; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_7_uop_switch = slots_7_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3964 = issue_slots_7_grant ? issue_slots_7_uop_switch : _GEN_3865; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_debug_tsrc = slots_8_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3967 = issue_slots_8_grant ? issue_slots_8_uop_debug_tsrc : _GEN_3868; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_debug_fsrc = slots_8_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3968 = issue_slots_8_grant ? issue_slots_8_uop_debug_fsrc : _GEN_3869; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_bp_xcpt_if = slots_8_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3969 = issue_slots_8_grant ? issue_slots_8_uop_bp_xcpt_if : _GEN_3870; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_bp_debug_if = slots_8_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3970 = issue_slots_8_grant ? issue_slots_8_uop_bp_debug_if : _GEN_3871; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_xcpt_ma_if = slots_8_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3971 = issue_slots_8_grant ? issue_slots_8_uop_xcpt_ma_if : _GEN_3872; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_xcpt_ae_if = slots_8_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3972 = issue_slots_8_grant ? issue_slots_8_uop_xcpt_ae_if : _GEN_3873; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_xcpt_pf_if = slots_8_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3973 = issue_slots_8_grant ? issue_slots_8_uop_xcpt_pf_if : _GEN_3874; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_fp_single = slots_8_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3974 = issue_slots_8_grant ? issue_slots_8_uop_fp_single : _GEN_3875; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_fp_val = slots_8_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3975 = issue_slots_8_grant ? issue_slots_8_uop_fp_val : _GEN_3876; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_frs3_en = slots_8_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3976 = issue_slots_8_grant ? issue_slots_8_uop_frs3_en : _GEN_3877; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_lrs2_rtype = slots_8_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3977 = issue_slots_8_grant ? issue_slots_8_uop_lrs2_rtype : _GEN_3878; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_lrs1_rtype = slots_8_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3978 = issue_slots_8_grant ? issue_slots_8_uop_lrs1_rtype : _GEN_3879; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_dst_rtype = slots_8_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3979 = issue_slots_8_grant ? issue_slots_8_uop_dst_rtype : _GEN_3880; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_ldst_val = slots_8_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3980 = issue_slots_8_grant ? issue_slots_8_uop_ldst_val : _GEN_3881; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_8_uop_lrs3 = slots_8_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3981 = issue_slots_8_grant ? issue_slots_8_uop_lrs3 : _GEN_3882; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_8_uop_lrs2 = slots_8_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3982 = issue_slots_8_grant ? issue_slots_8_uop_lrs2 : _GEN_3883; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_8_uop_lrs1 = slots_8_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3983 = issue_slots_8_grant ? issue_slots_8_uop_lrs1 : _GEN_3884; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_8_uop_ldst = slots_8_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_3984 = issue_slots_8_grant ? issue_slots_8_uop_ldst : _GEN_3885; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_ldst_is_rs1 = slots_8_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3985 = issue_slots_8_grant ? issue_slots_8_uop_ldst_is_rs1 : _GEN_3886; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_flush_on_commit = slots_8_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3986 = issue_slots_8_grant ? issue_slots_8_uop_flush_on_commit : _GEN_3887; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_unique = slots_8_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3987 = issue_slots_8_grant ? issue_slots_8_uop_is_unique : _GEN_3888; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_sys_pc2epc = slots_8_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3988 = issue_slots_8_grant ? issue_slots_8_uop_is_sys_pc2epc : _GEN_3889; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_uses_stq = slots_8_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3989 = issue_slots_8_grant ? issue_slots_8_uop_uses_stq : _GEN_3890; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_uses_ldq = slots_8_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3990 = issue_slots_8_grant ? issue_slots_8_uop_uses_ldq : _GEN_3891; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_amo = slots_8_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3991 = issue_slots_8_grant ? issue_slots_8_uop_is_amo : _GEN_3892; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_fencei = slots_8_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3992 = issue_slots_8_grant ? issue_slots_8_uop_is_fencei : _GEN_3893; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_fence = slots_8_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3993 = issue_slots_8_grant ? issue_slots_8_uop_is_fence : _GEN_3894; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_mem_signed = slots_8_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3994 = issue_slots_8_grant ? issue_slots_8_uop_mem_signed : _GEN_3895; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_mem_size = slots_8_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_3995 = issue_slots_8_grant ? issue_slots_8_uop_mem_size : _GEN_3896; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_8_uop_mem_cmd = slots_8_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_3996 = issue_slots_8_grant ? issue_slots_8_uop_mem_cmd : _GEN_3897; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_bypassable = slots_8_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3997 = issue_slots_8_grant ? issue_slots_8_uop_bypassable : _GEN_3898; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_8_uop_exc_cause = slots_8_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_3998 = issue_slots_8_grant ? issue_slots_8_uop_exc_cause : _GEN_3899; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_exception = slots_8_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_3999 = issue_slots_8_grant ? issue_slots_8_uop_exception : _GEN_3900; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_8_uop_stale_pdst = slots_8_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4000 = issue_slots_8_grant ? issue_slots_8_uop_stale_pdst : _GEN_3901; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_ppred_busy = slots_8_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4001 = issue_slots_8_grant ? issue_slots_8_uop_ppred_busy : _GEN_3902; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_prs3_busy = slots_8_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4002 = issue_slots_8_grant ? issue_slots_8_uop_prs3_busy : _GEN_3903; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_prs2_busy = slots_8_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4003 = issue_slots_8_grant ? issue_slots_8_uop_prs2_busy : _GEN_3904; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_prs1_busy = slots_8_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4004 = issue_slots_8_grant ? issue_slots_8_uop_prs1_busy : _GEN_3905; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_8_uop_ppred = slots_8_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4005 = issue_slots_8_grant ? issue_slots_8_uop_ppred : _GEN_3906; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_8_uop_prs3 = slots_8_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4006 = issue_slots_8_grant ? issue_slots_8_uop_prs3 : _GEN_3907; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_8_uop_prs2 = slots_8_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4007 = issue_slots_8_grant ? issue_slots_8_uop_prs2 : _GEN_3908; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_8_uop_prs1 = slots_8_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4008 = issue_slots_8_grant ? issue_slots_8_uop_prs1 : _GEN_3909; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_8_uop_pdst = slots_8_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4009 = issue_slots_8_grant ? issue_slots_8_uop_pdst : _GEN_3910; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_rxq_idx = slots_8_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4010 = issue_slots_8_grant ? issue_slots_8_uop_rxq_idx : _GEN_3911; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_8_uop_stq_idx = slots_8_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4011 = issue_slots_8_grant ? issue_slots_8_uop_stq_idx : _GEN_3912; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_8_uop_ldq_idx = slots_8_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4012 = issue_slots_8_grant ? issue_slots_8_uop_ldq_idx : _GEN_3913; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_8_uop_rob_idx = slots_8_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4013 = issue_slots_8_grant ? issue_slots_8_uop_rob_idx : _GEN_3914; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_8_uop_csr_addr = slots_8_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4014 = issue_slots_8_grant ? issue_slots_8_uop_csr_addr : _GEN_3915; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_8_uop_imm_packed = slots_8_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_4015 = issue_slots_8_grant ? issue_slots_8_uop_imm_packed : _GEN_3916; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_taken = slots_8_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4016 = issue_slots_8_grant ? issue_slots_8_uop_taken : _GEN_3917; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_8_uop_pc_lob = slots_8_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4017 = issue_slots_8_grant ? issue_slots_8_uop_pc_lob : _GEN_3918; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_edge_inst = slots_8_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4018 = issue_slots_8_grant ? issue_slots_8_uop_edge_inst : _GEN_3919; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_8_uop_ftq_idx = slots_8_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4019 = issue_slots_8_grant ? issue_slots_8_uop_ftq_idx : _GEN_3920; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_8_uop_br_tag = slots_8_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4020 = issue_slots_8_grant ? issue_slots_8_uop_br_tag : _GEN_3921; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_8_uop_br_mask = slots_8_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4021 = issue_slots_8_grant ? issue_slots_8_uop_br_mask : _GEN_3922; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_sfb = slots_8_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4022 = issue_slots_8_grant ? issue_slots_8_uop_is_sfb : _GEN_3923; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_jal = slots_8_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4023 = issue_slots_8_grant ? issue_slots_8_uop_is_jal : _GEN_3924; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_jalr = slots_8_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4024 = issue_slots_8_grant ? issue_slots_8_uop_is_jalr : _GEN_3925; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_br = slots_8_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4025 = issue_slots_8_grant ? issue_slots_8_uop_is_br : _GEN_3926; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_iw_p2_poisoned = slots_8_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4026 = issue_slots_8_grant ? issue_slots_8_uop_iw_p2_poisoned : _GEN_3927; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_iw_p1_poisoned = slots_8_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4027 = issue_slots_8_grant ? issue_slots_8_uop_iw_p1_poisoned : _GEN_3928; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_iw_state = slots_8_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4028 = issue_slots_8_grant ? issue_slots_8_uop_iw_state : _GEN_3929; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_ctrl_op3_sel = slots_8_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4029 = issue_slots_8_grant ? issue_slots_8_uop_ctrl_op3_sel : _GEN_3930; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_ctrl_is_std = slots_8_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4030 = issue_slots_8_grant ? issue_slots_8_uop_ctrl_is_std : _GEN_3931; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_ctrl_is_sta = slots_8_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4031 = issue_slots_8_grant ? issue_slots_8_uop_ctrl_is_sta : _GEN_3932; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_ctrl_is_load = slots_8_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4032 = issue_slots_8_grant ? issue_slots_8_uop_ctrl_is_load : _GEN_3933; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_8_uop_ctrl_csr_cmd = slots_8_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4033 = issue_slots_8_grant ? issue_slots_8_uop_ctrl_csr_cmd : _GEN_3934; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_ctrl_fcn_dw = slots_8_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4034 = issue_slots_8_grant ? issue_slots_8_uop_ctrl_fcn_dw : _GEN_3935; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_8_uop_ctrl_op_fcn = slots_8_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4035 = issue_slots_8_grant ? issue_slots_8_uop_ctrl_op_fcn : _GEN_3936; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_8_uop_ctrl_imm_sel = slots_8_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4036 = issue_slots_8_grant ? issue_slots_8_uop_ctrl_imm_sel : _GEN_3937; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_8_uop_ctrl_op2_sel = slots_8_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4037 = issue_slots_8_grant ? issue_slots_8_uop_ctrl_op2_sel : _GEN_3938; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_ctrl_op1_sel = slots_8_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4038 = issue_slots_8_grant ? issue_slots_8_uop_ctrl_op1_sel : _GEN_3939; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_8_uop_ctrl_br_type = slots_8_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4039 = issue_slots_8_grant ? issue_slots_8_uop_ctrl_br_type : _GEN_3940; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_4040 = issue_slots_8_grant ? issue_slots_8_uop_fu_code : _GEN_3941; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_8_uop_iq_type = slots_8_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4041 = issue_slots_8_grant ? issue_slots_8_uop_iq_type : _GEN_3942; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_8_uop_debug_pc = slots_8_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_4042 = issue_slots_8_grant ? issue_slots_8_uop_debug_pc : _GEN_3943; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_rvc = slots_8_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4043 = issue_slots_8_grant ? issue_slots_8_uop_is_rvc : _GEN_3944; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_8_uop_debug_inst = slots_8_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4044 = issue_slots_8_grant ? issue_slots_8_uop_debug_inst : _GEN_3945; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_8_uop_inst = slots_8_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4045 = issue_slots_8_grant ? issue_slots_8_uop_inst : _GEN_3946; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_8_uop_uopc = slots_8_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4046 = issue_slots_8_grant ? issue_slots_8_uop_uopc : _GEN_3947; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_8_uop_address_num = slots_8_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4047 = issue_slots_8_grant ? issue_slots_8_uop_address_num : _GEN_3948; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_8_uop_rob_inst_idx = slots_8_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4048 = issue_slots_8_grant ? issue_slots_8_uop_rob_inst_idx : _GEN_3949; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_8_uop_self_index = slots_8_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4049 = issue_slots_8_grant ? issue_slots_8_uop_self_index : _GEN_3950; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_8_uop_split_num = slots_8_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4050 = issue_slots_8_grant ? issue_slots_8_uop_split_num : _GEN_3951; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_8_uop_op2_sel = slots_8_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4051 = issue_slots_8_grant ? issue_slots_8_uop_op2_sel : _GEN_3952; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_8_uop_op1_sel = slots_8_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4052 = issue_slots_8_grant ? issue_slots_8_uop_op1_sel : _GEN_3953; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_8_uop_stale_pflag = slots_8_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4053 = issue_slots_8_grant ? issue_slots_8_uop_stale_pflag : _GEN_3954; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_pflag_busy = slots_8_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4054 = issue_slots_8_grant ? issue_slots_8_uop_pflag_busy : _GEN_3955; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_8_uop_pwflag = slots_8_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4055 = issue_slots_8_grant ? issue_slots_8_uop_pwflag : _GEN_3956; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_8_uop_prflag = slots_8_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4056 = issue_slots_8_grant ? issue_slots_8_uop_prflag : _GEN_3957; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_wflag = slots_8_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4057 = issue_slots_8_grant ? issue_slots_8_uop_wflag : _GEN_3958; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_rflag = slots_8_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4058 = issue_slots_8_grant ? issue_slots_8_uop_rflag : _GEN_3959; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_8_uop_lrs3_rtype = slots_8_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4059 = issue_slots_8_grant ? issue_slots_8_uop_lrs3_rtype : _GEN_3960; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_8_uop_shift = slots_8_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4060 = issue_slots_8_grant ? issue_slots_8_uop_shift : _GEN_3961; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_is_unicore = slots_8_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4061 = issue_slots_8_grant ? issue_slots_8_uop_is_unicore : _GEN_3962; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_switch_off = slots_8_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4062 = issue_slots_8_grant ? issue_slots_8_uop_switch_off : _GEN_3963; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_8_uop_switch = slots_8_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4063 = issue_slots_8_grant ? issue_slots_8_uop_switch : _GEN_3964; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_debug_tsrc = slots_9_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4066 = issue_slots_9_grant ? issue_slots_9_uop_debug_tsrc : _GEN_3967; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_debug_fsrc = slots_9_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4067 = issue_slots_9_grant ? issue_slots_9_uop_debug_fsrc : _GEN_3968; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_bp_xcpt_if = slots_9_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4068 = issue_slots_9_grant ? issue_slots_9_uop_bp_xcpt_if : _GEN_3969; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_bp_debug_if = slots_9_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4069 = issue_slots_9_grant ? issue_slots_9_uop_bp_debug_if : _GEN_3970; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_xcpt_ma_if = slots_9_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4070 = issue_slots_9_grant ? issue_slots_9_uop_xcpt_ma_if : _GEN_3971; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_xcpt_ae_if = slots_9_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4071 = issue_slots_9_grant ? issue_slots_9_uop_xcpt_ae_if : _GEN_3972; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_xcpt_pf_if = slots_9_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4072 = issue_slots_9_grant ? issue_slots_9_uop_xcpt_pf_if : _GEN_3973; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_fp_single = slots_9_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4073 = issue_slots_9_grant ? issue_slots_9_uop_fp_single : _GEN_3974; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_fp_val = slots_9_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4074 = issue_slots_9_grant ? issue_slots_9_uop_fp_val : _GEN_3975; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_frs3_en = slots_9_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4075 = issue_slots_9_grant ? issue_slots_9_uop_frs3_en : _GEN_3976; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_lrs2_rtype = slots_9_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4076 = issue_slots_9_grant ? issue_slots_9_uop_lrs2_rtype : _GEN_3977; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_lrs1_rtype = slots_9_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4077 = issue_slots_9_grant ? issue_slots_9_uop_lrs1_rtype : _GEN_3978; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_dst_rtype = slots_9_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4078 = issue_slots_9_grant ? issue_slots_9_uop_dst_rtype : _GEN_3979; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_ldst_val = slots_9_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4079 = issue_slots_9_grant ? issue_slots_9_uop_ldst_val : _GEN_3980; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_9_uop_lrs3 = slots_9_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4080 = issue_slots_9_grant ? issue_slots_9_uop_lrs3 : _GEN_3981; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_9_uop_lrs2 = slots_9_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4081 = issue_slots_9_grant ? issue_slots_9_uop_lrs2 : _GEN_3982; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_9_uop_lrs1 = slots_9_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4082 = issue_slots_9_grant ? issue_slots_9_uop_lrs1 : _GEN_3983; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_9_uop_ldst = slots_9_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4083 = issue_slots_9_grant ? issue_slots_9_uop_ldst : _GEN_3984; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_ldst_is_rs1 = slots_9_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4084 = issue_slots_9_grant ? issue_slots_9_uop_ldst_is_rs1 : _GEN_3985; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_flush_on_commit = slots_9_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4085 = issue_slots_9_grant ? issue_slots_9_uop_flush_on_commit : _GEN_3986; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_unique = slots_9_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4086 = issue_slots_9_grant ? issue_slots_9_uop_is_unique : _GEN_3987; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_sys_pc2epc = slots_9_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4087 = issue_slots_9_grant ? issue_slots_9_uop_is_sys_pc2epc : _GEN_3988; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_uses_stq = slots_9_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4088 = issue_slots_9_grant ? issue_slots_9_uop_uses_stq : _GEN_3989; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_uses_ldq = slots_9_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4089 = issue_slots_9_grant ? issue_slots_9_uop_uses_ldq : _GEN_3990; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_amo = slots_9_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4090 = issue_slots_9_grant ? issue_slots_9_uop_is_amo : _GEN_3991; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_fencei = slots_9_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4091 = issue_slots_9_grant ? issue_slots_9_uop_is_fencei : _GEN_3992; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_fence = slots_9_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4092 = issue_slots_9_grant ? issue_slots_9_uop_is_fence : _GEN_3993; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_mem_signed = slots_9_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4093 = issue_slots_9_grant ? issue_slots_9_uop_mem_signed : _GEN_3994; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_mem_size = slots_9_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4094 = issue_slots_9_grant ? issue_slots_9_uop_mem_size : _GEN_3995; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_9_uop_mem_cmd = slots_9_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4095 = issue_slots_9_grant ? issue_slots_9_uop_mem_cmd : _GEN_3996; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_bypassable = slots_9_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4096 = issue_slots_9_grant ? issue_slots_9_uop_bypassable : _GEN_3997; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_9_uop_exc_cause = slots_9_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_4097 = issue_slots_9_grant ? issue_slots_9_uop_exc_cause : _GEN_3998; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_exception = slots_9_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4098 = issue_slots_9_grant ? issue_slots_9_uop_exception : _GEN_3999; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_9_uop_stale_pdst = slots_9_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4099 = issue_slots_9_grant ? issue_slots_9_uop_stale_pdst : _GEN_4000; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_ppred_busy = slots_9_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4100 = issue_slots_9_grant ? issue_slots_9_uop_ppred_busy : _GEN_4001; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_prs3_busy = slots_9_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4101 = issue_slots_9_grant ? issue_slots_9_uop_prs3_busy : _GEN_4002; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_prs2_busy = slots_9_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4102 = issue_slots_9_grant ? issue_slots_9_uop_prs2_busy : _GEN_4003; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_prs1_busy = slots_9_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4103 = issue_slots_9_grant ? issue_slots_9_uop_prs1_busy : _GEN_4004; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_9_uop_ppred = slots_9_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4104 = issue_slots_9_grant ? issue_slots_9_uop_ppred : _GEN_4005; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_9_uop_prs3 = slots_9_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4105 = issue_slots_9_grant ? issue_slots_9_uop_prs3 : _GEN_4006; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_9_uop_prs2 = slots_9_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4106 = issue_slots_9_grant ? issue_slots_9_uop_prs2 : _GEN_4007; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_9_uop_prs1 = slots_9_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4107 = issue_slots_9_grant ? issue_slots_9_uop_prs1 : _GEN_4008; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_9_uop_pdst = slots_9_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4108 = issue_slots_9_grant ? issue_slots_9_uop_pdst : _GEN_4009; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_rxq_idx = slots_9_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4109 = issue_slots_9_grant ? issue_slots_9_uop_rxq_idx : _GEN_4010; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_9_uop_stq_idx = slots_9_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4110 = issue_slots_9_grant ? issue_slots_9_uop_stq_idx : _GEN_4011; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_9_uop_ldq_idx = slots_9_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4111 = issue_slots_9_grant ? issue_slots_9_uop_ldq_idx : _GEN_4012; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_9_uop_rob_idx = slots_9_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4112 = issue_slots_9_grant ? issue_slots_9_uop_rob_idx : _GEN_4013; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_9_uop_csr_addr = slots_9_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4113 = issue_slots_9_grant ? issue_slots_9_uop_csr_addr : _GEN_4014; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_9_uop_imm_packed = slots_9_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_4114 = issue_slots_9_grant ? issue_slots_9_uop_imm_packed : _GEN_4015; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_taken = slots_9_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4115 = issue_slots_9_grant ? issue_slots_9_uop_taken : _GEN_4016; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_9_uop_pc_lob = slots_9_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4116 = issue_slots_9_grant ? issue_slots_9_uop_pc_lob : _GEN_4017; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_edge_inst = slots_9_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4117 = issue_slots_9_grant ? issue_slots_9_uop_edge_inst : _GEN_4018; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_9_uop_ftq_idx = slots_9_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4118 = issue_slots_9_grant ? issue_slots_9_uop_ftq_idx : _GEN_4019; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_9_uop_br_tag = slots_9_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4119 = issue_slots_9_grant ? issue_slots_9_uop_br_tag : _GEN_4020; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_9_uop_br_mask = slots_9_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4120 = issue_slots_9_grant ? issue_slots_9_uop_br_mask : _GEN_4021; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_sfb = slots_9_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4121 = issue_slots_9_grant ? issue_slots_9_uop_is_sfb : _GEN_4022; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_jal = slots_9_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4122 = issue_slots_9_grant ? issue_slots_9_uop_is_jal : _GEN_4023; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_jalr = slots_9_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4123 = issue_slots_9_grant ? issue_slots_9_uop_is_jalr : _GEN_4024; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_br = slots_9_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4124 = issue_slots_9_grant ? issue_slots_9_uop_is_br : _GEN_4025; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_iw_p2_poisoned = slots_9_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4125 = issue_slots_9_grant ? issue_slots_9_uop_iw_p2_poisoned : _GEN_4026; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_iw_p1_poisoned = slots_9_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4126 = issue_slots_9_grant ? issue_slots_9_uop_iw_p1_poisoned : _GEN_4027; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_iw_state = slots_9_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4127 = issue_slots_9_grant ? issue_slots_9_uop_iw_state : _GEN_4028; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_ctrl_op3_sel = slots_9_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4128 = issue_slots_9_grant ? issue_slots_9_uop_ctrl_op3_sel : _GEN_4029; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_ctrl_is_std = slots_9_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4129 = issue_slots_9_grant ? issue_slots_9_uop_ctrl_is_std : _GEN_4030; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_ctrl_is_sta = slots_9_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4130 = issue_slots_9_grant ? issue_slots_9_uop_ctrl_is_sta : _GEN_4031; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_ctrl_is_load = slots_9_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4131 = issue_slots_9_grant ? issue_slots_9_uop_ctrl_is_load : _GEN_4032; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_9_uop_ctrl_csr_cmd = slots_9_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4132 = issue_slots_9_grant ? issue_slots_9_uop_ctrl_csr_cmd : _GEN_4033; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_ctrl_fcn_dw = slots_9_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4133 = issue_slots_9_grant ? issue_slots_9_uop_ctrl_fcn_dw : _GEN_4034; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_9_uop_ctrl_op_fcn = slots_9_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4134 = issue_slots_9_grant ? issue_slots_9_uop_ctrl_op_fcn : _GEN_4035; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_9_uop_ctrl_imm_sel = slots_9_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4135 = issue_slots_9_grant ? issue_slots_9_uop_ctrl_imm_sel : _GEN_4036; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_9_uop_ctrl_op2_sel = slots_9_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4136 = issue_slots_9_grant ? issue_slots_9_uop_ctrl_op2_sel : _GEN_4037; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_ctrl_op1_sel = slots_9_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4137 = issue_slots_9_grant ? issue_slots_9_uop_ctrl_op1_sel : _GEN_4038; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_9_uop_ctrl_br_type = slots_9_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4138 = issue_slots_9_grant ? issue_slots_9_uop_ctrl_br_type : _GEN_4039; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_4139 = issue_slots_9_grant ? issue_slots_9_uop_fu_code : _GEN_4040; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_9_uop_iq_type = slots_9_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4140 = issue_slots_9_grant ? issue_slots_9_uop_iq_type : _GEN_4041; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_9_uop_debug_pc = slots_9_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_4141 = issue_slots_9_grant ? issue_slots_9_uop_debug_pc : _GEN_4042; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_rvc = slots_9_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4142 = issue_slots_9_grant ? issue_slots_9_uop_is_rvc : _GEN_4043; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_9_uop_debug_inst = slots_9_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4143 = issue_slots_9_grant ? issue_slots_9_uop_debug_inst : _GEN_4044; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_9_uop_inst = slots_9_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4144 = issue_slots_9_grant ? issue_slots_9_uop_inst : _GEN_4045; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_9_uop_uopc = slots_9_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4145 = issue_slots_9_grant ? issue_slots_9_uop_uopc : _GEN_4046; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_9_uop_address_num = slots_9_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4146 = issue_slots_9_grant ? issue_slots_9_uop_address_num : _GEN_4047; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_9_uop_rob_inst_idx = slots_9_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4147 = issue_slots_9_grant ? issue_slots_9_uop_rob_inst_idx : _GEN_4048; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_9_uop_self_index = slots_9_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4148 = issue_slots_9_grant ? issue_slots_9_uop_self_index : _GEN_4049; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_9_uop_split_num = slots_9_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4149 = issue_slots_9_grant ? issue_slots_9_uop_split_num : _GEN_4050; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_9_uop_op2_sel = slots_9_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4150 = issue_slots_9_grant ? issue_slots_9_uop_op2_sel : _GEN_4051; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_9_uop_op1_sel = slots_9_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4151 = issue_slots_9_grant ? issue_slots_9_uop_op1_sel : _GEN_4052; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_9_uop_stale_pflag = slots_9_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4152 = issue_slots_9_grant ? issue_slots_9_uop_stale_pflag : _GEN_4053; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_pflag_busy = slots_9_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4153 = issue_slots_9_grant ? issue_slots_9_uop_pflag_busy : _GEN_4054; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_9_uop_pwflag = slots_9_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4154 = issue_slots_9_grant ? issue_slots_9_uop_pwflag : _GEN_4055; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_9_uop_prflag = slots_9_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4155 = issue_slots_9_grant ? issue_slots_9_uop_prflag : _GEN_4056; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_wflag = slots_9_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4156 = issue_slots_9_grant ? issue_slots_9_uop_wflag : _GEN_4057; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_rflag = slots_9_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4157 = issue_slots_9_grant ? issue_slots_9_uop_rflag : _GEN_4058; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_9_uop_lrs3_rtype = slots_9_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4158 = issue_slots_9_grant ? issue_slots_9_uop_lrs3_rtype : _GEN_4059; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_9_uop_shift = slots_9_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4159 = issue_slots_9_grant ? issue_slots_9_uop_shift : _GEN_4060; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_is_unicore = slots_9_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4160 = issue_slots_9_grant ? issue_slots_9_uop_is_unicore : _GEN_4061; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_switch_off = slots_9_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4161 = issue_slots_9_grant ? issue_slots_9_uop_switch_off : _GEN_4062; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_9_uop_switch = slots_9_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4162 = issue_slots_9_grant ? issue_slots_9_uop_switch : _GEN_4063; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_debug_tsrc = slots_10_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4165 = issue_slots_10_grant ? issue_slots_10_uop_debug_tsrc : _GEN_4066; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_debug_fsrc = slots_10_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4166 = issue_slots_10_grant ? issue_slots_10_uop_debug_fsrc : _GEN_4067; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_bp_xcpt_if = slots_10_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4167 = issue_slots_10_grant ? issue_slots_10_uop_bp_xcpt_if : _GEN_4068; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_bp_debug_if = slots_10_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4168 = issue_slots_10_grant ? issue_slots_10_uop_bp_debug_if : _GEN_4069; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_xcpt_ma_if = slots_10_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4169 = issue_slots_10_grant ? issue_slots_10_uop_xcpt_ma_if : _GEN_4070; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_xcpt_ae_if = slots_10_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4170 = issue_slots_10_grant ? issue_slots_10_uop_xcpt_ae_if : _GEN_4071; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_xcpt_pf_if = slots_10_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4171 = issue_slots_10_grant ? issue_slots_10_uop_xcpt_pf_if : _GEN_4072; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_fp_single = slots_10_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4172 = issue_slots_10_grant ? issue_slots_10_uop_fp_single : _GEN_4073; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_fp_val = slots_10_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4173 = issue_slots_10_grant ? issue_slots_10_uop_fp_val : _GEN_4074; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_frs3_en = slots_10_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4174 = issue_slots_10_grant ? issue_slots_10_uop_frs3_en : _GEN_4075; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_lrs2_rtype = slots_10_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4175 = issue_slots_10_grant ? issue_slots_10_uop_lrs2_rtype : _GEN_4076; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_lrs1_rtype = slots_10_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4176 = issue_slots_10_grant ? issue_slots_10_uop_lrs1_rtype : _GEN_4077; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_dst_rtype = slots_10_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4177 = issue_slots_10_grant ? issue_slots_10_uop_dst_rtype : _GEN_4078; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_ldst_val = slots_10_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4178 = issue_slots_10_grant ? issue_slots_10_uop_ldst_val : _GEN_4079; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_10_uop_lrs3 = slots_10_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4179 = issue_slots_10_grant ? issue_slots_10_uop_lrs3 : _GEN_4080; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_10_uop_lrs2 = slots_10_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4180 = issue_slots_10_grant ? issue_slots_10_uop_lrs2 : _GEN_4081; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_10_uop_lrs1 = slots_10_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4181 = issue_slots_10_grant ? issue_slots_10_uop_lrs1 : _GEN_4082; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_10_uop_ldst = slots_10_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4182 = issue_slots_10_grant ? issue_slots_10_uop_ldst : _GEN_4083; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_ldst_is_rs1 = slots_10_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4183 = issue_slots_10_grant ? issue_slots_10_uop_ldst_is_rs1 : _GEN_4084; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_flush_on_commit = slots_10_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4184 = issue_slots_10_grant ? issue_slots_10_uop_flush_on_commit : _GEN_4085; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_unique = slots_10_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4185 = issue_slots_10_grant ? issue_slots_10_uop_is_unique : _GEN_4086; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_sys_pc2epc = slots_10_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4186 = issue_slots_10_grant ? issue_slots_10_uop_is_sys_pc2epc : _GEN_4087; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_uses_stq = slots_10_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4187 = issue_slots_10_grant ? issue_slots_10_uop_uses_stq : _GEN_4088; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_uses_ldq = slots_10_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4188 = issue_slots_10_grant ? issue_slots_10_uop_uses_ldq : _GEN_4089; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_amo = slots_10_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4189 = issue_slots_10_grant ? issue_slots_10_uop_is_amo : _GEN_4090; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_fencei = slots_10_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4190 = issue_slots_10_grant ? issue_slots_10_uop_is_fencei : _GEN_4091; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_fence = slots_10_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4191 = issue_slots_10_grant ? issue_slots_10_uop_is_fence : _GEN_4092; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_mem_signed = slots_10_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4192 = issue_slots_10_grant ? issue_slots_10_uop_mem_signed : _GEN_4093; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_mem_size = slots_10_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4193 = issue_slots_10_grant ? issue_slots_10_uop_mem_size : _GEN_4094; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_10_uop_mem_cmd = slots_10_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4194 = issue_slots_10_grant ? issue_slots_10_uop_mem_cmd : _GEN_4095; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_bypassable = slots_10_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4195 = issue_slots_10_grant ? issue_slots_10_uop_bypassable : _GEN_4096; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_10_uop_exc_cause = slots_10_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_4196 = issue_slots_10_grant ? issue_slots_10_uop_exc_cause : _GEN_4097; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_exception = slots_10_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4197 = issue_slots_10_grant ? issue_slots_10_uop_exception : _GEN_4098; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_10_uop_stale_pdst = slots_10_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4198 = issue_slots_10_grant ? issue_slots_10_uop_stale_pdst : _GEN_4099; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_ppred_busy = slots_10_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4199 = issue_slots_10_grant ? issue_slots_10_uop_ppred_busy : _GEN_4100; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_prs3_busy = slots_10_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4200 = issue_slots_10_grant ? issue_slots_10_uop_prs3_busy : _GEN_4101; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_prs2_busy = slots_10_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4201 = issue_slots_10_grant ? issue_slots_10_uop_prs2_busy : _GEN_4102; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_prs1_busy = slots_10_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4202 = issue_slots_10_grant ? issue_slots_10_uop_prs1_busy : _GEN_4103; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_10_uop_ppred = slots_10_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4203 = issue_slots_10_grant ? issue_slots_10_uop_ppred : _GEN_4104; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_10_uop_prs3 = slots_10_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4204 = issue_slots_10_grant ? issue_slots_10_uop_prs3 : _GEN_4105; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_10_uop_prs2 = slots_10_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4205 = issue_slots_10_grant ? issue_slots_10_uop_prs2 : _GEN_4106; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_10_uop_prs1 = slots_10_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4206 = issue_slots_10_grant ? issue_slots_10_uop_prs1 : _GEN_4107; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_10_uop_pdst = slots_10_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4207 = issue_slots_10_grant ? issue_slots_10_uop_pdst : _GEN_4108; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_rxq_idx = slots_10_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4208 = issue_slots_10_grant ? issue_slots_10_uop_rxq_idx : _GEN_4109; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_10_uop_stq_idx = slots_10_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4209 = issue_slots_10_grant ? issue_slots_10_uop_stq_idx : _GEN_4110; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_10_uop_ldq_idx = slots_10_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4210 = issue_slots_10_grant ? issue_slots_10_uop_ldq_idx : _GEN_4111; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_10_uop_rob_idx = slots_10_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4211 = issue_slots_10_grant ? issue_slots_10_uop_rob_idx : _GEN_4112; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_10_uop_csr_addr = slots_10_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4212 = issue_slots_10_grant ? issue_slots_10_uop_csr_addr : _GEN_4113; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_10_uop_imm_packed = slots_10_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_4213 = issue_slots_10_grant ? issue_slots_10_uop_imm_packed : _GEN_4114; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_taken = slots_10_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4214 = issue_slots_10_grant ? issue_slots_10_uop_taken : _GEN_4115; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_10_uop_pc_lob = slots_10_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4215 = issue_slots_10_grant ? issue_slots_10_uop_pc_lob : _GEN_4116; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_edge_inst = slots_10_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4216 = issue_slots_10_grant ? issue_slots_10_uop_edge_inst : _GEN_4117; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_10_uop_ftq_idx = slots_10_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4217 = issue_slots_10_grant ? issue_slots_10_uop_ftq_idx : _GEN_4118; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_10_uop_br_tag = slots_10_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4218 = issue_slots_10_grant ? issue_slots_10_uop_br_tag : _GEN_4119; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_10_uop_br_mask = slots_10_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4219 = issue_slots_10_grant ? issue_slots_10_uop_br_mask : _GEN_4120; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_sfb = slots_10_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4220 = issue_slots_10_grant ? issue_slots_10_uop_is_sfb : _GEN_4121; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_jal = slots_10_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4221 = issue_slots_10_grant ? issue_slots_10_uop_is_jal : _GEN_4122; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_jalr = slots_10_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4222 = issue_slots_10_grant ? issue_slots_10_uop_is_jalr : _GEN_4123; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_br = slots_10_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4223 = issue_slots_10_grant ? issue_slots_10_uop_is_br : _GEN_4124; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_iw_p2_poisoned = slots_10_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4224 = issue_slots_10_grant ? issue_slots_10_uop_iw_p2_poisoned : _GEN_4125; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_iw_p1_poisoned = slots_10_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4225 = issue_slots_10_grant ? issue_slots_10_uop_iw_p1_poisoned : _GEN_4126; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_iw_state = slots_10_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4226 = issue_slots_10_grant ? issue_slots_10_uop_iw_state : _GEN_4127; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_ctrl_op3_sel = slots_10_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4227 = issue_slots_10_grant ? issue_slots_10_uop_ctrl_op3_sel : _GEN_4128; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_ctrl_is_std = slots_10_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4228 = issue_slots_10_grant ? issue_slots_10_uop_ctrl_is_std : _GEN_4129; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_ctrl_is_sta = slots_10_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4229 = issue_slots_10_grant ? issue_slots_10_uop_ctrl_is_sta : _GEN_4130; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_ctrl_is_load = slots_10_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4230 = issue_slots_10_grant ? issue_slots_10_uop_ctrl_is_load : _GEN_4131; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_10_uop_ctrl_csr_cmd = slots_10_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4231 = issue_slots_10_grant ? issue_slots_10_uop_ctrl_csr_cmd : _GEN_4132; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_ctrl_fcn_dw = slots_10_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4232 = issue_slots_10_grant ? issue_slots_10_uop_ctrl_fcn_dw : _GEN_4133; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_10_uop_ctrl_op_fcn = slots_10_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4233 = issue_slots_10_grant ? issue_slots_10_uop_ctrl_op_fcn : _GEN_4134; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_10_uop_ctrl_imm_sel = slots_10_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4234 = issue_slots_10_grant ? issue_slots_10_uop_ctrl_imm_sel : _GEN_4135; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_10_uop_ctrl_op2_sel = slots_10_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4235 = issue_slots_10_grant ? issue_slots_10_uop_ctrl_op2_sel : _GEN_4136; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_ctrl_op1_sel = slots_10_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4236 = issue_slots_10_grant ? issue_slots_10_uop_ctrl_op1_sel : _GEN_4137; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_10_uop_ctrl_br_type = slots_10_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4237 = issue_slots_10_grant ? issue_slots_10_uop_ctrl_br_type : _GEN_4138; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_4238 = issue_slots_10_grant ? issue_slots_10_uop_fu_code : _GEN_4139; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_10_uop_iq_type = slots_10_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4239 = issue_slots_10_grant ? issue_slots_10_uop_iq_type : _GEN_4140; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_10_uop_debug_pc = slots_10_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_4240 = issue_slots_10_grant ? issue_slots_10_uop_debug_pc : _GEN_4141; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_rvc = slots_10_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4241 = issue_slots_10_grant ? issue_slots_10_uop_is_rvc : _GEN_4142; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_10_uop_debug_inst = slots_10_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4242 = issue_slots_10_grant ? issue_slots_10_uop_debug_inst : _GEN_4143; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_10_uop_inst = slots_10_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4243 = issue_slots_10_grant ? issue_slots_10_uop_inst : _GEN_4144; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_10_uop_uopc = slots_10_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4244 = issue_slots_10_grant ? issue_slots_10_uop_uopc : _GEN_4145; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_10_uop_address_num = slots_10_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4245 = issue_slots_10_grant ? issue_slots_10_uop_address_num : _GEN_4146; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_10_uop_rob_inst_idx = slots_10_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4246 = issue_slots_10_grant ? issue_slots_10_uop_rob_inst_idx : _GEN_4147; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_10_uop_self_index = slots_10_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4247 = issue_slots_10_grant ? issue_slots_10_uop_self_index : _GEN_4148; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_10_uop_split_num = slots_10_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4248 = issue_slots_10_grant ? issue_slots_10_uop_split_num : _GEN_4149; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_10_uop_op2_sel = slots_10_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4249 = issue_slots_10_grant ? issue_slots_10_uop_op2_sel : _GEN_4150; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_10_uop_op1_sel = slots_10_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4250 = issue_slots_10_grant ? issue_slots_10_uop_op1_sel : _GEN_4151; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_10_uop_stale_pflag = slots_10_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4251 = issue_slots_10_grant ? issue_slots_10_uop_stale_pflag : _GEN_4152; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_pflag_busy = slots_10_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4252 = issue_slots_10_grant ? issue_slots_10_uop_pflag_busy : _GEN_4153; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_10_uop_pwflag = slots_10_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4253 = issue_slots_10_grant ? issue_slots_10_uop_pwflag : _GEN_4154; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_10_uop_prflag = slots_10_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4254 = issue_slots_10_grant ? issue_slots_10_uop_prflag : _GEN_4155; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_wflag = slots_10_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4255 = issue_slots_10_grant ? issue_slots_10_uop_wflag : _GEN_4156; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_rflag = slots_10_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4256 = issue_slots_10_grant ? issue_slots_10_uop_rflag : _GEN_4157; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_10_uop_lrs3_rtype = slots_10_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4257 = issue_slots_10_grant ? issue_slots_10_uop_lrs3_rtype : _GEN_4158; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_10_uop_shift = slots_10_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4258 = issue_slots_10_grant ? issue_slots_10_uop_shift : _GEN_4159; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_is_unicore = slots_10_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4259 = issue_slots_10_grant ? issue_slots_10_uop_is_unicore : _GEN_4160; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_switch_off = slots_10_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4260 = issue_slots_10_grant ? issue_slots_10_uop_switch_off : _GEN_4161; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_10_uop_switch = slots_10_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4261 = issue_slots_10_grant ? issue_slots_10_uop_switch : _GEN_4162; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_debug_tsrc = slots_11_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4264 = issue_slots_11_grant ? issue_slots_11_uop_debug_tsrc : _GEN_4165; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_debug_fsrc = slots_11_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4265 = issue_slots_11_grant ? issue_slots_11_uop_debug_fsrc : _GEN_4166; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_bp_xcpt_if = slots_11_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4266 = issue_slots_11_grant ? issue_slots_11_uop_bp_xcpt_if : _GEN_4167; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_bp_debug_if = slots_11_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4267 = issue_slots_11_grant ? issue_slots_11_uop_bp_debug_if : _GEN_4168; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_xcpt_ma_if = slots_11_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4268 = issue_slots_11_grant ? issue_slots_11_uop_xcpt_ma_if : _GEN_4169; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_xcpt_ae_if = slots_11_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4269 = issue_slots_11_grant ? issue_slots_11_uop_xcpt_ae_if : _GEN_4170; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_xcpt_pf_if = slots_11_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4270 = issue_slots_11_grant ? issue_slots_11_uop_xcpt_pf_if : _GEN_4171; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_fp_single = slots_11_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4271 = issue_slots_11_grant ? issue_slots_11_uop_fp_single : _GEN_4172; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_fp_val = slots_11_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4272 = issue_slots_11_grant ? issue_slots_11_uop_fp_val : _GEN_4173; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_frs3_en = slots_11_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4273 = issue_slots_11_grant ? issue_slots_11_uop_frs3_en : _GEN_4174; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_lrs2_rtype = slots_11_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4274 = issue_slots_11_grant ? issue_slots_11_uop_lrs2_rtype : _GEN_4175; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_lrs1_rtype = slots_11_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4275 = issue_slots_11_grant ? issue_slots_11_uop_lrs1_rtype : _GEN_4176; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_dst_rtype = slots_11_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4276 = issue_slots_11_grant ? issue_slots_11_uop_dst_rtype : _GEN_4177; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_ldst_val = slots_11_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4277 = issue_slots_11_grant ? issue_slots_11_uop_ldst_val : _GEN_4178; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_11_uop_lrs3 = slots_11_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4278 = issue_slots_11_grant ? issue_slots_11_uop_lrs3 : _GEN_4179; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_11_uop_lrs2 = slots_11_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4279 = issue_slots_11_grant ? issue_slots_11_uop_lrs2 : _GEN_4180; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_11_uop_lrs1 = slots_11_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4280 = issue_slots_11_grant ? issue_slots_11_uop_lrs1 : _GEN_4181; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_11_uop_ldst = slots_11_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4281 = issue_slots_11_grant ? issue_slots_11_uop_ldst : _GEN_4182; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_ldst_is_rs1 = slots_11_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4282 = issue_slots_11_grant ? issue_slots_11_uop_ldst_is_rs1 : _GEN_4183; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_flush_on_commit = slots_11_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4283 = issue_slots_11_grant ? issue_slots_11_uop_flush_on_commit : _GEN_4184; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_unique = slots_11_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4284 = issue_slots_11_grant ? issue_slots_11_uop_is_unique : _GEN_4185; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_sys_pc2epc = slots_11_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4285 = issue_slots_11_grant ? issue_slots_11_uop_is_sys_pc2epc : _GEN_4186; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_uses_stq = slots_11_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4286 = issue_slots_11_grant ? issue_slots_11_uop_uses_stq : _GEN_4187; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_uses_ldq = slots_11_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4287 = issue_slots_11_grant ? issue_slots_11_uop_uses_ldq : _GEN_4188; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_amo = slots_11_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4288 = issue_slots_11_grant ? issue_slots_11_uop_is_amo : _GEN_4189; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_fencei = slots_11_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4289 = issue_slots_11_grant ? issue_slots_11_uop_is_fencei : _GEN_4190; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_fence = slots_11_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4290 = issue_slots_11_grant ? issue_slots_11_uop_is_fence : _GEN_4191; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_mem_signed = slots_11_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4291 = issue_slots_11_grant ? issue_slots_11_uop_mem_signed : _GEN_4192; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_mem_size = slots_11_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4292 = issue_slots_11_grant ? issue_slots_11_uop_mem_size : _GEN_4193; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_11_uop_mem_cmd = slots_11_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4293 = issue_slots_11_grant ? issue_slots_11_uop_mem_cmd : _GEN_4194; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_bypassable = slots_11_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4294 = issue_slots_11_grant ? issue_slots_11_uop_bypassable : _GEN_4195; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_11_uop_exc_cause = slots_11_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_4295 = issue_slots_11_grant ? issue_slots_11_uop_exc_cause : _GEN_4196; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_exception = slots_11_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4296 = issue_slots_11_grant ? issue_slots_11_uop_exception : _GEN_4197; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_11_uop_stale_pdst = slots_11_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4297 = issue_slots_11_grant ? issue_slots_11_uop_stale_pdst : _GEN_4198; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_ppred_busy = slots_11_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4298 = issue_slots_11_grant ? issue_slots_11_uop_ppred_busy : _GEN_4199; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_prs3_busy = slots_11_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4299 = issue_slots_11_grant ? issue_slots_11_uop_prs3_busy : _GEN_4200; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_prs2_busy = slots_11_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4300 = issue_slots_11_grant ? issue_slots_11_uop_prs2_busy : _GEN_4201; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_prs1_busy = slots_11_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4301 = issue_slots_11_grant ? issue_slots_11_uop_prs1_busy : _GEN_4202; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_11_uop_ppred = slots_11_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4302 = issue_slots_11_grant ? issue_slots_11_uop_ppred : _GEN_4203; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_11_uop_prs3 = slots_11_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4303 = issue_slots_11_grant ? issue_slots_11_uop_prs3 : _GEN_4204; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_11_uop_prs2 = slots_11_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4304 = issue_slots_11_grant ? issue_slots_11_uop_prs2 : _GEN_4205; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_11_uop_prs1 = slots_11_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4305 = issue_slots_11_grant ? issue_slots_11_uop_prs1 : _GEN_4206; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_11_uop_pdst = slots_11_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4306 = issue_slots_11_grant ? issue_slots_11_uop_pdst : _GEN_4207; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_rxq_idx = slots_11_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4307 = issue_slots_11_grant ? issue_slots_11_uop_rxq_idx : _GEN_4208; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_11_uop_stq_idx = slots_11_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4308 = issue_slots_11_grant ? issue_slots_11_uop_stq_idx : _GEN_4209; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_11_uop_ldq_idx = slots_11_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4309 = issue_slots_11_grant ? issue_slots_11_uop_ldq_idx : _GEN_4210; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_11_uop_rob_idx = slots_11_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4310 = issue_slots_11_grant ? issue_slots_11_uop_rob_idx : _GEN_4211; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_11_uop_csr_addr = slots_11_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4311 = issue_slots_11_grant ? issue_slots_11_uop_csr_addr : _GEN_4212; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_11_uop_imm_packed = slots_11_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_4312 = issue_slots_11_grant ? issue_slots_11_uop_imm_packed : _GEN_4213; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_taken = slots_11_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4313 = issue_slots_11_grant ? issue_slots_11_uop_taken : _GEN_4214; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_11_uop_pc_lob = slots_11_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4314 = issue_slots_11_grant ? issue_slots_11_uop_pc_lob : _GEN_4215; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_edge_inst = slots_11_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4315 = issue_slots_11_grant ? issue_slots_11_uop_edge_inst : _GEN_4216; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_11_uop_ftq_idx = slots_11_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4316 = issue_slots_11_grant ? issue_slots_11_uop_ftq_idx : _GEN_4217; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_11_uop_br_tag = slots_11_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4317 = issue_slots_11_grant ? issue_slots_11_uop_br_tag : _GEN_4218; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_11_uop_br_mask = slots_11_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4318 = issue_slots_11_grant ? issue_slots_11_uop_br_mask : _GEN_4219; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_sfb = slots_11_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4319 = issue_slots_11_grant ? issue_slots_11_uop_is_sfb : _GEN_4220; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_jal = slots_11_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4320 = issue_slots_11_grant ? issue_slots_11_uop_is_jal : _GEN_4221; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_jalr = slots_11_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4321 = issue_slots_11_grant ? issue_slots_11_uop_is_jalr : _GEN_4222; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_br = slots_11_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4322 = issue_slots_11_grant ? issue_slots_11_uop_is_br : _GEN_4223; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_iw_p2_poisoned = slots_11_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4323 = issue_slots_11_grant ? issue_slots_11_uop_iw_p2_poisoned : _GEN_4224; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_iw_p1_poisoned = slots_11_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4324 = issue_slots_11_grant ? issue_slots_11_uop_iw_p1_poisoned : _GEN_4225; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_iw_state = slots_11_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4325 = issue_slots_11_grant ? issue_slots_11_uop_iw_state : _GEN_4226; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_ctrl_op3_sel = slots_11_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4326 = issue_slots_11_grant ? issue_slots_11_uop_ctrl_op3_sel : _GEN_4227; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_ctrl_is_std = slots_11_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4327 = issue_slots_11_grant ? issue_slots_11_uop_ctrl_is_std : _GEN_4228; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_ctrl_is_sta = slots_11_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4328 = issue_slots_11_grant ? issue_slots_11_uop_ctrl_is_sta : _GEN_4229; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_ctrl_is_load = slots_11_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4329 = issue_slots_11_grant ? issue_slots_11_uop_ctrl_is_load : _GEN_4230; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_11_uop_ctrl_csr_cmd = slots_11_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4330 = issue_slots_11_grant ? issue_slots_11_uop_ctrl_csr_cmd : _GEN_4231; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_ctrl_fcn_dw = slots_11_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4331 = issue_slots_11_grant ? issue_slots_11_uop_ctrl_fcn_dw : _GEN_4232; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_11_uop_ctrl_op_fcn = slots_11_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4332 = issue_slots_11_grant ? issue_slots_11_uop_ctrl_op_fcn : _GEN_4233; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_11_uop_ctrl_imm_sel = slots_11_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4333 = issue_slots_11_grant ? issue_slots_11_uop_ctrl_imm_sel : _GEN_4234; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_11_uop_ctrl_op2_sel = slots_11_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4334 = issue_slots_11_grant ? issue_slots_11_uop_ctrl_op2_sel : _GEN_4235; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_ctrl_op1_sel = slots_11_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4335 = issue_slots_11_grant ? issue_slots_11_uop_ctrl_op1_sel : _GEN_4236; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_11_uop_ctrl_br_type = slots_11_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4336 = issue_slots_11_grant ? issue_slots_11_uop_ctrl_br_type : _GEN_4237; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_4337 = issue_slots_11_grant ? issue_slots_11_uop_fu_code : _GEN_4238; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_11_uop_iq_type = slots_11_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4338 = issue_slots_11_grant ? issue_slots_11_uop_iq_type : _GEN_4239; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_11_uop_debug_pc = slots_11_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_4339 = issue_slots_11_grant ? issue_slots_11_uop_debug_pc : _GEN_4240; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_rvc = slots_11_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4340 = issue_slots_11_grant ? issue_slots_11_uop_is_rvc : _GEN_4241; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_11_uop_debug_inst = slots_11_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4341 = issue_slots_11_grant ? issue_slots_11_uop_debug_inst : _GEN_4242; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_11_uop_inst = slots_11_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4342 = issue_slots_11_grant ? issue_slots_11_uop_inst : _GEN_4243; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_11_uop_uopc = slots_11_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4343 = issue_slots_11_grant ? issue_slots_11_uop_uopc : _GEN_4244; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_11_uop_address_num = slots_11_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4344 = issue_slots_11_grant ? issue_slots_11_uop_address_num : _GEN_4245; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_11_uop_rob_inst_idx = slots_11_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4345 = issue_slots_11_grant ? issue_slots_11_uop_rob_inst_idx : _GEN_4246; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_11_uop_self_index = slots_11_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4346 = issue_slots_11_grant ? issue_slots_11_uop_self_index : _GEN_4247; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_11_uop_split_num = slots_11_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4347 = issue_slots_11_grant ? issue_slots_11_uop_split_num : _GEN_4248; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_11_uop_op2_sel = slots_11_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4348 = issue_slots_11_grant ? issue_slots_11_uop_op2_sel : _GEN_4249; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_11_uop_op1_sel = slots_11_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4349 = issue_slots_11_grant ? issue_slots_11_uop_op1_sel : _GEN_4250; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_11_uop_stale_pflag = slots_11_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4350 = issue_slots_11_grant ? issue_slots_11_uop_stale_pflag : _GEN_4251; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_pflag_busy = slots_11_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4351 = issue_slots_11_grant ? issue_slots_11_uop_pflag_busy : _GEN_4252; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_11_uop_pwflag = slots_11_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4352 = issue_slots_11_grant ? issue_slots_11_uop_pwflag : _GEN_4253; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_11_uop_prflag = slots_11_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4353 = issue_slots_11_grant ? issue_slots_11_uop_prflag : _GEN_4254; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_wflag = slots_11_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4354 = issue_slots_11_grant ? issue_slots_11_uop_wflag : _GEN_4255; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_rflag = slots_11_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4355 = issue_slots_11_grant ? issue_slots_11_uop_rflag : _GEN_4256; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_11_uop_lrs3_rtype = slots_11_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4356 = issue_slots_11_grant ? issue_slots_11_uop_lrs3_rtype : _GEN_4257; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_11_uop_shift = slots_11_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4357 = issue_slots_11_grant ? issue_slots_11_uop_shift : _GEN_4258; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_is_unicore = slots_11_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4358 = issue_slots_11_grant ? issue_slots_11_uop_is_unicore : _GEN_4259; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_switch_off = slots_11_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4359 = issue_slots_11_grant ? issue_slots_11_uop_switch_off : _GEN_4260; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_11_uop_switch = slots_11_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4360 = issue_slots_11_grant ? issue_slots_11_uop_switch : _GEN_4261; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_debug_tsrc = slots_12_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4363 = issue_slots_12_grant ? issue_slots_12_uop_debug_tsrc : _GEN_4264; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_debug_fsrc = slots_12_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4364 = issue_slots_12_grant ? issue_slots_12_uop_debug_fsrc : _GEN_4265; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_bp_xcpt_if = slots_12_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4365 = issue_slots_12_grant ? issue_slots_12_uop_bp_xcpt_if : _GEN_4266; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_bp_debug_if = slots_12_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4366 = issue_slots_12_grant ? issue_slots_12_uop_bp_debug_if : _GEN_4267; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_xcpt_ma_if = slots_12_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4367 = issue_slots_12_grant ? issue_slots_12_uop_xcpt_ma_if : _GEN_4268; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_xcpt_ae_if = slots_12_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4368 = issue_slots_12_grant ? issue_slots_12_uop_xcpt_ae_if : _GEN_4269; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_xcpt_pf_if = slots_12_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4369 = issue_slots_12_grant ? issue_slots_12_uop_xcpt_pf_if : _GEN_4270; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_fp_single = slots_12_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4370 = issue_slots_12_grant ? issue_slots_12_uop_fp_single : _GEN_4271; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_fp_val = slots_12_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4371 = issue_slots_12_grant ? issue_slots_12_uop_fp_val : _GEN_4272; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_frs3_en = slots_12_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4372 = issue_slots_12_grant ? issue_slots_12_uop_frs3_en : _GEN_4273; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_lrs2_rtype = slots_12_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4373 = issue_slots_12_grant ? issue_slots_12_uop_lrs2_rtype : _GEN_4274; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_lrs1_rtype = slots_12_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4374 = issue_slots_12_grant ? issue_slots_12_uop_lrs1_rtype : _GEN_4275; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_dst_rtype = slots_12_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4375 = issue_slots_12_grant ? issue_slots_12_uop_dst_rtype : _GEN_4276; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_ldst_val = slots_12_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4376 = issue_slots_12_grant ? issue_slots_12_uop_ldst_val : _GEN_4277; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_12_uop_lrs3 = slots_12_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4377 = issue_slots_12_grant ? issue_slots_12_uop_lrs3 : _GEN_4278; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_12_uop_lrs2 = slots_12_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4378 = issue_slots_12_grant ? issue_slots_12_uop_lrs2 : _GEN_4279; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_12_uop_lrs1 = slots_12_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4379 = issue_slots_12_grant ? issue_slots_12_uop_lrs1 : _GEN_4280; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_12_uop_ldst = slots_12_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4380 = issue_slots_12_grant ? issue_slots_12_uop_ldst : _GEN_4281; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_ldst_is_rs1 = slots_12_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4381 = issue_slots_12_grant ? issue_slots_12_uop_ldst_is_rs1 : _GEN_4282; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_flush_on_commit = slots_12_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4382 = issue_slots_12_grant ? issue_slots_12_uop_flush_on_commit : _GEN_4283; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_unique = slots_12_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4383 = issue_slots_12_grant ? issue_slots_12_uop_is_unique : _GEN_4284; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_sys_pc2epc = slots_12_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4384 = issue_slots_12_grant ? issue_slots_12_uop_is_sys_pc2epc : _GEN_4285; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_uses_stq = slots_12_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4385 = issue_slots_12_grant ? issue_slots_12_uop_uses_stq : _GEN_4286; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_uses_ldq = slots_12_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4386 = issue_slots_12_grant ? issue_slots_12_uop_uses_ldq : _GEN_4287; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_amo = slots_12_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4387 = issue_slots_12_grant ? issue_slots_12_uop_is_amo : _GEN_4288; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_fencei = slots_12_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4388 = issue_slots_12_grant ? issue_slots_12_uop_is_fencei : _GEN_4289; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_fence = slots_12_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4389 = issue_slots_12_grant ? issue_slots_12_uop_is_fence : _GEN_4290; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_mem_signed = slots_12_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4390 = issue_slots_12_grant ? issue_slots_12_uop_mem_signed : _GEN_4291; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_mem_size = slots_12_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4391 = issue_slots_12_grant ? issue_slots_12_uop_mem_size : _GEN_4292; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_12_uop_mem_cmd = slots_12_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4392 = issue_slots_12_grant ? issue_slots_12_uop_mem_cmd : _GEN_4293; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_bypassable = slots_12_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4393 = issue_slots_12_grant ? issue_slots_12_uop_bypassable : _GEN_4294; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_12_uop_exc_cause = slots_12_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_4394 = issue_slots_12_grant ? issue_slots_12_uop_exc_cause : _GEN_4295; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_exception = slots_12_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4395 = issue_slots_12_grant ? issue_slots_12_uop_exception : _GEN_4296; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_12_uop_stale_pdst = slots_12_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4396 = issue_slots_12_grant ? issue_slots_12_uop_stale_pdst : _GEN_4297; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_ppred_busy = slots_12_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4397 = issue_slots_12_grant ? issue_slots_12_uop_ppred_busy : _GEN_4298; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_prs3_busy = slots_12_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4398 = issue_slots_12_grant ? issue_slots_12_uop_prs3_busy : _GEN_4299; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_prs2_busy = slots_12_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4399 = issue_slots_12_grant ? issue_slots_12_uop_prs2_busy : _GEN_4300; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_prs1_busy = slots_12_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4400 = issue_slots_12_grant ? issue_slots_12_uop_prs1_busy : _GEN_4301; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_12_uop_ppred = slots_12_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4401 = issue_slots_12_grant ? issue_slots_12_uop_ppred : _GEN_4302; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_12_uop_prs3 = slots_12_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4402 = issue_slots_12_grant ? issue_slots_12_uop_prs3 : _GEN_4303; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_12_uop_prs2 = slots_12_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4403 = issue_slots_12_grant ? issue_slots_12_uop_prs2 : _GEN_4304; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_12_uop_prs1 = slots_12_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4404 = issue_slots_12_grant ? issue_slots_12_uop_prs1 : _GEN_4305; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_12_uop_pdst = slots_12_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4405 = issue_slots_12_grant ? issue_slots_12_uop_pdst : _GEN_4306; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_rxq_idx = slots_12_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4406 = issue_slots_12_grant ? issue_slots_12_uop_rxq_idx : _GEN_4307; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_12_uop_stq_idx = slots_12_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4407 = issue_slots_12_grant ? issue_slots_12_uop_stq_idx : _GEN_4308; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_12_uop_ldq_idx = slots_12_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4408 = issue_slots_12_grant ? issue_slots_12_uop_ldq_idx : _GEN_4309; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_12_uop_rob_idx = slots_12_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4409 = issue_slots_12_grant ? issue_slots_12_uop_rob_idx : _GEN_4310; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_12_uop_csr_addr = slots_12_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4410 = issue_slots_12_grant ? issue_slots_12_uop_csr_addr : _GEN_4311; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_12_uop_imm_packed = slots_12_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_4411 = issue_slots_12_grant ? issue_slots_12_uop_imm_packed : _GEN_4312; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_taken = slots_12_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4412 = issue_slots_12_grant ? issue_slots_12_uop_taken : _GEN_4313; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_12_uop_pc_lob = slots_12_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4413 = issue_slots_12_grant ? issue_slots_12_uop_pc_lob : _GEN_4314; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_edge_inst = slots_12_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4414 = issue_slots_12_grant ? issue_slots_12_uop_edge_inst : _GEN_4315; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_12_uop_ftq_idx = slots_12_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4415 = issue_slots_12_grant ? issue_slots_12_uop_ftq_idx : _GEN_4316; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_12_uop_br_tag = slots_12_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4416 = issue_slots_12_grant ? issue_slots_12_uop_br_tag : _GEN_4317; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_12_uop_br_mask = slots_12_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4417 = issue_slots_12_grant ? issue_slots_12_uop_br_mask : _GEN_4318; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_sfb = slots_12_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4418 = issue_slots_12_grant ? issue_slots_12_uop_is_sfb : _GEN_4319; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_jal = slots_12_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4419 = issue_slots_12_grant ? issue_slots_12_uop_is_jal : _GEN_4320; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_jalr = slots_12_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4420 = issue_slots_12_grant ? issue_slots_12_uop_is_jalr : _GEN_4321; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_br = slots_12_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4421 = issue_slots_12_grant ? issue_slots_12_uop_is_br : _GEN_4322; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_iw_p2_poisoned = slots_12_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4422 = issue_slots_12_grant ? issue_slots_12_uop_iw_p2_poisoned : _GEN_4323; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_iw_p1_poisoned = slots_12_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4423 = issue_slots_12_grant ? issue_slots_12_uop_iw_p1_poisoned : _GEN_4324; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_iw_state = slots_12_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4424 = issue_slots_12_grant ? issue_slots_12_uop_iw_state : _GEN_4325; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_ctrl_op3_sel = slots_12_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4425 = issue_slots_12_grant ? issue_slots_12_uop_ctrl_op3_sel : _GEN_4326; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_ctrl_is_std = slots_12_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4426 = issue_slots_12_grant ? issue_slots_12_uop_ctrl_is_std : _GEN_4327; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_ctrl_is_sta = slots_12_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4427 = issue_slots_12_grant ? issue_slots_12_uop_ctrl_is_sta : _GEN_4328; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_ctrl_is_load = slots_12_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4428 = issue_slots_12_grant ? issue_slots_12_uop_ctrl_is_load : _GEN_4329; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_12_uop_ctrl_csr_cmd = slots_12_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4429 = issue_slots_12_grant ? issue_slots_12_uop_ctrl_csr_cmd : _GEN_4330; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_ctrl_fcn_dw = slots_12_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4430 = issue_slots_12_grant ? issue_slots_12_uop_ctrl_fcn_dw : _GEN_4331; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_12_uop_ctrl_op_fcn = slots_12_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4431 = issue_slots_12_grant ? issue_slots_12_uop_ctrl_op_fcn : _GEN_4332; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_12_uop_ctrl_imm_sel = slots_12_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4432 = issue_slots_12_grant ? issue_slots_12_uop_ctrl_imm_sel : _GEN_4333; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_12_uop_ctrl_op2_sel = slots_12_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4433 = issue_slots_12_grant ? issue_slots_12_uop_ctrl_op2_sel : _GEN_4334; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_ctrl_op1_sel = slots_12_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4434 = issue_slots_12_grant ? issue_slots_12_uop_ctrl_op1_sel : _GEN_4335; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_12_uop_ctrl_br_type = slots_12_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4435 = issue_slots_12_grant ? issue_slots_12_uop_ctrl_br_type : _GEN_4336; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_4436 = issue_slots_12_grant ? issue_slots_12_uop_fu_code : _GEN_4337; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_12_uop_iq_type = slots_12_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4437 = issue_slots_12_grant ? issue_slots_12_uop_iq_type : _GEN_4338; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_12_uop_debug_pc = slots_12_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_4438 = issue_slots_12_grant ? issue_slots_12_uop_debug_pc : _GEN_4339; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_rvc = slots_12_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4439 = issue_slots_12_grant ? issue_slots_12_uop_is_rvc : _GEN_4340; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_12_uop_debug_inst = slots_12_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4440 = issue_slots_12_grant ? issue_slots_12_uop_debug_inst : _GEN_4341; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_12_uop_inst = slots_12_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4441 = issue_slots_12_grant ? issue_slots_12_uop_inst : _GEN_4342; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_12_uop_uopc = slots_12_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4442 = issue_slots_12_grant ? issue_slots_12_uop_uopc : _GEN_4343; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_12_uop_address_num = slots_12_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4443 = issue_slots_12_grant ? issue_slots_12_uop_address_num : _GEN_4344; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_12_uop_rob_inst_idx = slots_12_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4444 = issue_slots_12_grant ? issue_slots_12_uop_rob_inst_idx : _GEN_4345; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_12_uop_self_index = slots_12_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4445 = issue_slots_12_grant ? issue_slots_12_uop_self_index : _GEN_4346; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_12_uop_split_num = slots_12_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4446 = issue_slots_12_grant ? issue_slots_12_uop_split_num : _GEN_4347; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_12_uop_op2_sel = slots_12_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4447 = issue_slots_12_grant ? issue_slots_12_uop_op2_sel : _GEN_4348; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_12_uop_op1_sel = slots_12_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4448 = issue_slots_12_grant ? issue_slots_12_uop_op1_sel : _GEN_4349; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_12_uop_stale_pflag = slots_12_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4449 = issue_slots_12_grant ? issue_slots_12_uop_stale_pflag : _GEN_4350; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_pflag_busy = slots_12_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4450 = issue_slots_12_grant ? issue_slots_12_uop_pflag_busy : _GEN_4351; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_12_uop_pwflag = slots_12_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4451 = issue_slots_12_grant ? issue_slots_12_uop_pwflag : _GEN_4352; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_12_uop_prflag = slots_12_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4452 = issue_slots_12_grant ? issue_slots_12_uop_prflag : _GEN_4353; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_wflag = slots_12_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4453 = issue_slots_12_grant ? issue_slots_12_uop_wflag : _GEN_4354; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_rflag = slots_12_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4454 = issue_slots_12_grant ? issue_slots_12_uop_rflag : _GEN_4355; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_12_uop_lrs3_rtype = slots_12_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4455 = issue_slots_12_grant ? issue_slots_12_uop_lrs3_rtype : _GEN_4356; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_12_uop_shift = slots_12_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4456 = issue_slots_12_grant ? issue_slots_12_uop_shift : _GEN_4357; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_is_unicore = slots_12_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4457 = issue_slots_12_grant ? issue_slots_12_uop_is_unicore : _GEN_4358; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_switch_off = slots_12_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4458 = issue_slots_12_grant ? issue_slots_12_uop_switch_off : _GEN_4359; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_12_uop_switch = slots_12_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4459 = issue_slots_12_grant ? issue_slots_12_uop_switch : _GEN_4360; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_debug_tsrc = slots_13_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4462 = issue_slots_13_grant ? issue_slots_13_uop_debug_tsrc : _GEN_4363; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_debug_fsrc = slots_13_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4463 = issue_slots_13_grant ? issue_slots_13_uop_debug_fsrc : _GEN_4364; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_bp_xcpt_if = slots_13_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4464 = issue_slots_13_grant ? issue_slots_13_uop_bp_xcpt_if : _GEN_4365; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_bp_debug_if = slots_13_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4465 = issue_slots_13_grant ? issue_slots_13_uop_bp_debug_if : _GEN_4366; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_xcpt_ma_if = slots_13_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4466 = issue_slots_13_grant ? issue_slots_13_uop_xcpt_ma_if : _GEN_4367; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_xcpt_ae_if = slots_13_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4467 = issue_slots_13_grant ? issue_slots_13_uop_xcpt_ae_if : _GEN_4368; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_xcpt_pf_if = slots_13_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4468 = issue_slots_13_grant ? issue_slots_13_uop_xcpt_pf_if : _GEN_4369; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_fp_single = slots_13_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4469 = issue_slots_13_grant ? issue_slots_13_uop_fp_single : _GEN_4370; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_fp_val = slots_13_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4470 = issue_slots_13_grant ? issue_slots_13_uop_fp_val : _GEN_4371; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_frs3_en = slots_13_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4471 = issue_slots_13_grant ? issue_slots_13_uop_frs3_en : _GEN_4372; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_lrs2_rtype = slots_13_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4472 = issue_slots_13_grant ? issue_slots_13_uop_lrs2_rtype : _GEN_4373; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_lrs1_rtype = slots_13_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4473 = issue_slots_13_grant ? issue_slots_13_uop_lrs1_rtype : _GEN_4374; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_dst_rtype = slots_13_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4474 = issue_slots_13_grant ? issue_slots_13_uop_dst_rtype : _GEN_4375; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_ldst_val = slots_13_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4475 = issue_slots_13_grant ? issue_slots_13_uop_ldst_val : _GEN_4376; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_13_uop_lrs3 = slots_13_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4476 = issue_slots_13_grant ? issue_slots_13_uop_lrs3 : _GEN_4377; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_13_uop_lrs2 = slots_13_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4477 = issue_slots_13_grant ? issue_slots_13_uop_lrs2 : _GEN_4378; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_13_uop_lrs1 = slots_13_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4478 = issue_slots_13_grant ? issue_slots_13_uop_lrs1 : _GEN_4379; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_13_uop_ldst = slots_13_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4479 = issue_slots_13_grant ? issue_slots_13_uop_ldst : _GEN_4380; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_ldst_is_rs1 = slots_13_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4480 = issue_slots_13_grant ? issue_slots_13_uop_ldst_is_rs1 : _GEN_4381; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_flush_on_commit = slots_13_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4481 = issue_slots_13_grant ? issue_slots_13_uop_flush_on_commit : _GEN_4382; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_unique = slots_13_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4482 = issue_slots_13_grant ? issue_slots_13_uop_is_unique : _GEN_4383; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_sys_pc2epc = slots_13_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4483 = issue_slots_13_grant ? issue_slots_13_uop_is_sys_pc2epc : _GEN_4384; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_uses_stq = slots_13_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4484 = issue_slots_13_grant ? issue_slots_13_uop_uses_stq : _GEN_4385; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_uses_ldq = slots_13_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4485 = issue_slots_13_grant ? issue_slots_13_uop_uses_ldq : _GEN_4386; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_amo = slots_13_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4486 = issue_slots_13_grant ? issue_slots_13_uop_is_amo : _GEN_4387; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_fencei = slots_13_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4487 = issue_slots_13_grant ? issue_slots_13_uop_is_fencei : _GEN_4388; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_fence = slots_13_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4488 = issue_slots_13_grant ? issue_slots_13_uop_is_fence : _GEN_4389; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_mem_signed = slots_13_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4489 = issue_slots_13_grant ? issue_slots_13_uop_mem_signed : _GEN_4390; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_mem_size = slots_13_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4490 = issue_slots_13_grant ? issue_slots_13_uop_mem_size : _GEN_4391; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_13_uop_mem_cmd = slots_13_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4491 = issue_slots_13_grant ? issue_slots_13_uop_mem_cmd : _GEN_4392; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_bypassable = slots_13_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4492 = issue_slots_13_grant ? issue_slots_13_uop_bypassable : _GEN_4393; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_13_uop_exc_cause = slots_13_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_4493 = issue_slots_13_grant ? issue_slots_13_uop_exc_cause : _GEN_4394; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_exception = slots_13_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4494 = issue_slots_13_grant ? issue_slots_13_uop_exception : _GEN_4395; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_13_uop_stale_pdst = slots_13_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4495 = issue_slots_13_grant ? issue_slots_13_uop_stale_pdst : _GEN_4396; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_ppred_busy = slots_13_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4496 = issue_slots_13_grant ? issue_slots_13_uop_ppred_busy : _GEN_4397; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_prs3_busy = slots_13_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4497 = issue_slots_13_grant ? issue_slots_13_uop_prs3_busy : _GEN_4398; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_prs2_busy = slots_13_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4498 = issue_slots_13_grant ? issue_slots_13_uop_prs2_busy : _GEN_4399; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_prs1_busy = slots_13_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4499 = issue_slots_13_grant ? issue_slots_13_uop_prs1_busy : _GEN_4400; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_13_uop_ppred = slots_13_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4500 = issue_slots_13_grant ? issue_slots_13_uop_ppred : _GEN_4401; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_13_uop_prs3 = slots_13_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4501 = issue_slots_13_grant ? issue_slots_13_uop_prs3 : _GEN_4402; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_13_uop_prs2 = slots_13_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4502 = issue_slots_13_grant ? issue_slots_13_uop_prs2 : _GEN_4403; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_13_uop_prs1 = slots_13_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4503 = issue_slots_13_grant ? issue_slots_13_uop_prs1 : _GEN_4404; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_13_uop_pdst = slots_13_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4504 = issue_slots_13_grant ? issue_slots_13_uop_pdst : _GEN_4405; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_rxq_idx = slots_13_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4505 = issue_slots_13_grant ? issue_slots_13_uop_rxq_idx : _GEN_4406; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_13_uop_stq_idx = slots_13_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4506 = issue_slots_13_grant ? issue_slots_13_uop_stq_idx : _GEN_4407; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_13_uop_ldq_idx = slots_13_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4507 = issue_slots_13_grant ? issue_slots_13_uop_ldq_idx : _GEN_4408; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_13_uop_rob_idx = slots_13_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4508 = issue_slots_13_grant ? issue_slots_13_uop_rob_idx : _GEN_4409; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_13_uop_csr_addr = slots_13_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4509 = issue_slots_13_grant ? issue_slots_13_uop_csr_addr : _GEN_4410; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_13_uop_imm_packed = slots_13_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_4510 = issue_slots_13_grant ? issue_slots_13_uop_imm_packed : _GEN_4411; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_taken = slots_13_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4511 = issue_slots_13_grant ? issue_slots_13_uop_taken : _GEN_4412; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_13_uop_pc_lob = slots_13_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4512 = issue_slots_13_grant ? issue_slots_13_uop_pc_lob : _GEN_4413; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_edge_inst = slots_13_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4513 = issue_slots_13_grant ? issue_slots_13_uop_edge_inst : _GEN_4414; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_13_uop_ftq_idx = slots_13_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4514 = issue_slots_13_grant ? issue_slots_13_uop_ftq_idx : _GEN_4415; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_13_uop_br_tag = slots_13_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4515 = issue_slots_13_grant ? issue_slots_13_uop_br_tag : _GEN_4416; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_13_uop_br_mask = slots_13_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4516 = issue_slots_13_grant ? issue_slots_13_uop_br_mask : _GEN_4417; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_sfb = slots_13_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4517 = issue_slots_13_grant ? issue_slots_13_uop_is_sfb : _GEN_4418; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_jal = slots_13_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4518 = issue_slots_13_grant ? issue_slots_13_uop_is_jal : _GEN_4419; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_jalr = slots_13_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4519 = issue_slots_13_grant ? issue_slots_13_uop_is_jalr : _GEN_4420; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_br = slots_13_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4520 = issue_slots_13_grant ? issue_slots_13_uop_is_br : _GEN_4421; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_iw_p2_poisoned = slots_13_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4521 = issue_slots_13_grant ? issue_slots_13_uop_iw_p2_poisoned : _GEN_4422; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_iw_p1_poisoned = slots_13_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4522 = issue_slots_13_grant ? issue_slots_13_uop_iw_p1_poisoned : _GEN_4423; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_iw_state = slots_13_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4523 = issue_slots_13_grant ? issue_slots_13_uop_iw_state : _GEN_4424; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_ctrl_op3_sel = slots_13_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4524 = issue_slots_13_grant ? issue_slots_13_uop_ctrl_op3_sel : _GEN_4425; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_ctrl_is_std = slots_13_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4525 = issue_slots_13_grant ? issue_slots_13_uop_ctrl_is_std : _GEN_4426; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_ctrl_is_sta = slots_13_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4526 = issue_slots_13_grant ? issue_slots_13_uop_ctrl_is_sta : _GEN_4427; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_ctrl_is_load = slots_13_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4527 = issue_slots_13_grant ? issue_slots_13_uop_ctrl_is_load : _GEN_4428; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_13_uop_ctrl_csr_cmd = slots_13_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4528 = issue_slots_13_grant ? issue_slots_13_uop_ctrl_csr_cmd : _GEN_4429; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_ctrl_fcn_dw = slots_13_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4529 = issue_slots_13_grant ? issue_slots_13_uop_ctrl_fcn_dw : _GEN_4430; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_13_uop_ctrl_op_fcn = slots_13_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4530 = issue_slots_13_grant ? issue_slots_13_uop_ctrl_op_fcn : _GEN_4431; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_13_uop_ctrl_imm_sel = slots_13_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4531 = issue_slots_13_grant ? issue_slots_13_uop_ctrl_imm_sel : _GEN_4432; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_13_uop_ctrl_op2_sel = slots_13_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4532 = issue_slots_13_grant ? issue_slots_13_uop_ctrl_op2_sel : _GEN_4433; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_ctrl_op1_sel = slots_13_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4533 = issue_slots_13_grant ? issue_slots_13_uop_ctrl_op1_sel : _GEN_4434; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_13_uop_ctrl_br_type = slots_13_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4534 = issue_slots_13_grant ? issue_slots_13_uop_ctrl_br_type : _GEN_4435; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_4535 = issue_slots_13_grant ? issue_slots_13_uop_fu_code : _GEN_4436; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_13_uop_iq_type = slots_13_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4536 = issue_slots_13_grant ? issue_slots_13_uop_iq_type : _GEN_4437; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_13_uop_debug_pc = slots_13_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_4537 = issue_slots_13_grant ? issue_slots_13_uop_debug_pc : _GEN_4438; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_rvc = slots_13_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4538 = issue_slots_13_grant ? issue_slots_13_uop_is_rvc : _GEN_4439; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_13_uop_debug_inst = slots_13_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4539 = issue_slots_13_grant ? issue_slots_13_uop_debug_inst : _GEN_4440; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_13_uop_inst = slots_13_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4540 = issue_slots_13_grant ? issue_slots_13_uop_inst : _GEN_4441; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_13_uop_uopc = slots_13_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4541 = issue_slots_13_grant ? issue_slots_13_uop_uopc : _GEN_4442; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_13_uop_address_num = slots_13_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4542 = issue_slots_13_grant ? issue_slots_13_uop_address_num : _GEN_4443; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_13_uop_rob_inst_idx = slots_13_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4543 = issue_slots_13_grant ? issue_slots_13_uop_rob_inst_idx : _GEN_4444; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_13_uop_self_index = slots_13_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4544 = issue_slots_13_grant ? issue_slots_13_uop_self_index : _GEN_4445; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_13_uop_split_num = slots_13_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4545 = issue_slots_13_grant ? issue_slots_13_uop_split_num : _GEN_4446; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_13_uop_op2_sel = slots_13_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4546 = issue_slots_13_grant ? issue_slots_13_uop_op2_sel : _GEN_4447; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_13_uop_op1_sel = slots_13_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4547 = issue_slots_13_grant ? issue_slots_13_uop_op1_sel : _GEN_4448; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_13_uop_stale_pflag = slots_13_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4548 = issue_slots_13_grant ? issue_slots_13_uop_stale_pflag : _GEN_4449; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_pflag_busy = slots_13_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4549 = issue_slots_13_grant ? issue_slots_13_uop_pflag_busy : _GEN_4450; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_13_uop_pwflag = slots_13_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4550 = issue_slots_13_grant ? issue_slots_13_uop_pwflag : _GEN_4451; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_13_uop_prflag = slots_13_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4551 = issue_slots_13_grant ? issue_slots_13_uop_prflag : _GEN_4452; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_wflag = slots_13_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4552 = issue_slots_13_grant ? issue_slots_13_uop_wflag : _GEN_4453; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_rflag = slots_13_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4553 = issue_slots_13_grant ? issue_slots_13_uop_rflag : _GEN_4454; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_13_uop_lrs3_rtype = slots_13_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4554 = issue_slots_13_grant ? issue_slots_13_uop_lrs3_rtype : _GEN_4455; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_13_uop_shift = slots_13_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4555 = issue_slots_13_grant ? issue_slots_13_uop_shift : _GEN_4456; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_is_unicore = slots_13_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4556 = issue_slots_13_grant ? issue_slots_13_uop_is_unicore : _GEN_4457; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_switch_off = slots_13_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4557 = issue_slots_13_grant ? issue_slots_13_uop_switch_off : _GEN_4458; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_13_uop_switch = slots_13_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4558 = issue_slots_13_grant ? issue_slots_13_uop_switch : _GEN_4459; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_debug_tsrc = slots_14_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4561 = issue_slots_14_grant ? issue_slots_14_uop_debug_tsrc : _GEN_4462; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_debug_fsrc = slots_14_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4562 = issue_slots_14_grant ? issue_slots_14_uop_debug_fsrc : _GEN_4463; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_bp_xcpt_if = slots_14_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4563 = issue_slots_14_grant ? issue_slots_14_uop_bp_xcpt_if : _GEN_4464; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_bp_debug_if = slots_14_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4564 = issue_slots_14_grant ? issue_slots_14_uop_bp_debug_if : _GEN_4465; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_xcpt_ma_if = slots_14_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4565 = issue_slots_14_grant ? issue_slots_14_uop_xcpt_ma_if : _GEN_4466; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_xcpt_ae_if = slots_14_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4566 = issue_slots_14_grant ? issue_slots_14_uop_xcpt_ae_if : _GEN_4467; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_xcpt_pf_if = slots_14_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4567 = issue_slots_14_grant ? issue_slots_14_uop_xcpt_pf_if : _GEN_4468; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_fp_single = slots_14_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4568 = issue_slots_14_grant ? issue_slots_14_uop_fp_single : _GEN_4469; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_fp_val = slots_14_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4569 = issue_slots_14_grant ? issue_slots_14_uop_fp_val : _GEN_4470; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_frs3_en = slots_14_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4570 = issue_slots_14_grant ? issue_slots_14_uop_frs3_en : _GEN_4471; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_lrs2_rtype = slots_14_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4571 = issue_slots_14_grant ? issue_slots_14_uop_lrs2_rtype : _GEN_4472; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_lrs1_rtype = slots_14_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4572 = issue_slots_14_grant ? issue_slots_14_uop_lrs1_rtype : _GEN_4473; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_dst_rtype = slots_14_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4573 = issue_slots_14_grant ? issue_slots_14_uop_dst_rtype : _GEN_4474; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_ldst_val = slots_14_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4574 = issue_slots_14_grant ? issue_slots_14_uop_ldst_val : _GEN_4475; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_14_uop_lrs3 = slots_14_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4575 = issue_slots_14_grant ? issue_slots_14_uop_lrs3 : _GEN_4476; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_14_uop_lrs2 = slots_14_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4576 = issue_slots_14_grant ? issue_slots_14_uop_lrs2 : _GEN_4477; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_14_uop_lrs1 = slots_14_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4577 = issue_slots_14_grant ? issue_slots_14_uop_lrs1 : _GEN_4478; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_14_uop_ldst = slots_14_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4578 = issue_slots_14_grant ? issue_slots_14_uop_ldst : _GEN_4479; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_ldst_is_rs1 = slots_14_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4579 = issue_slots_14_grant ? issue_slots_14_uop_ldst_is_rs1 : _GEN_4480; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_flush_on_commit = slots_14_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4580 = issue_slots_14_grant ? issue_slots_14_uop_flush_on_commit : _GEN_4481; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_unique = slots_14_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4581 = issue_slots_14_grant ? issue_slots_14_uop_is_unique : _GEN_4482; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_sys_pc2epc = slots_14_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4582 = issue_slots_14_grant ? issue_slots_14_uop_is_sys_pc2epc : _GEN_4483; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_uses_stq = slots_14_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4583 = issue_slots_14_grant ? issue_slots_14_uop_uses_stq : _GEN_4484; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_uses_ldq = slots_14_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4584 = issue_slots_14_grant ? issue_slots_14_uop_uses_ldq : _GEN_4485; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_amo = slots_14_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4585 = issue_slots_14_grant ? issue_slots_14_uop_is_amo : _GEN_4486; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_fencei = slots_14_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4586 = issue_slots_14_grant ? issue_slots_14_uop_is_fencei : _GEN_4487; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_fence = slots_14_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4587 = issue_slots_14_grant ? issue_slots_14_uop_is_fence : _GEN_4488; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_mem_signed = slots_14_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4588 = issue_slots_14_grant ? issue_slots_14_uop_mem_signed : _GEN_4489; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_mem_size = slots_14_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4589 = issue_slots_14_grant ? issue_slots_14_uop_mem_size : _GEN_4490; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_14_uop_mem_cmd = slots_14_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4590 = issue_slots_14_grant ? issue_slots_14_uop_mem_cmd : _GEN_4491; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_bypassable = slots_14_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4591 = issue_slots_14_grant ? issue_slots_14_uop_bypassable : _GEN_4492; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [63:0] issue_slots_14_uop_exc_cause = slots_14_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] _GEN_4592 = issue_slots_14_grant ? issue_slots_14_uop_exc_cause : _GEN_4493; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_exception = slots_14_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4593 = issue_slots_14_grant ? issue_slots_14_uop_exception : _GEN_4494; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_14_uop_stale_pdst = slots_14_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4594 = issue_slots_14_grant ? issue_slots_14_uop_stale_pdst : _GEN_4495; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_ppred_busy = slots_14_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4595 = issue_slots_14_grant ? issue_slots_14_uop_ppred_busy : _GEN_4496; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_prs3_busy = slots_14_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4596 = issue_slots_14_grant ? issue_slots_14_uop_prs3_busy : _GEN_4497; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_prs2_busy = slots_14_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4597 = issue_slots_14_grant ? issue_slots_14_uop_prs2_busy : _GEN_4498; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_prs1_busy = slots_14_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4598 = issue_slots_14_grant ? issue_slots_14_uop_prs1_busy : _GEN_4499; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_14_uop_ppred = slots_14_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4599 = issue_slots_14_grant ? issue_slots_14_uop_ppred : _GEN_4500; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_14_uop_prs3 = slots_14_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4600 = issue_slots_14_grant ? issue_slots_14_uop_prs3 : _GEN_4501; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_14_uop_prs2 = slots_14_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4601 = issue_slots_14_grant ? issue_slots_14_uop_prs2 : _GEN_4502; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_14_uop_prs1 = slots_14_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4602 = issue_slots_14_grant ? issue_slots_14_uop_prs1 : _GEN_4503; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_14_uop_pdst = slots_14_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4603 = issue_slots_14_grant ? issue_slots_14_uop_pdst : _GEN_4504; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_rxq_idx = slots_14_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4604 = issue_slots_14_grant ? issue_slots_14_uop_rxq_idx : _GEN_4505; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_14_uop_stq_idx = slots_14_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4605 = issue_slots_14_grant ? issue_slots_14_uop_stq_idx : _GEN_4506; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_14_uop_ldq_idx = slots_14_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4606 = issue_slots_14_grant ? issue_slots_14_uop_ldq_idx : _GEN_4507; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_14_uop_rob_idx = slots_14_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4607 = issue_slots_14_grant ? issue_slots_14_uop_rob_idx : _GEN_4508; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_14_uop_csr_addr = slots_14_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4608 = issue_slots_14_grant ? issue_slots_14_uop_csr_addr : _GEN_4509; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [19:0] issue_slots_14_uop_imm_packed = slots_14_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] _GEN_4609 = issue_slots_14_grant ? issue_slots_14_uop_imm_packed : _GEN_4510; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_taken = slots_14_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4610 = issue_slots_14_grant ? issue_slots_14_uop_taken : _GEN_4511; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_14_uop_pc_lob = slots_14_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4611 = issue_slots_14_grant ? issue_slots_14_uop_pc_lob : _GEN_4512; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_edge_inst = slots_14_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4612 = issue_slots_14_grant ? issue_slots_14_uop_edge_inst : _GEN_4513; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [4:0] issue_slots_14_uop_ftq_idx = slots_14_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] _GEN_4613 = issue_slots_14_grant ? issue_slots_14_uop_ftq_idx : _GEN_4514; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_14_uop_br_tag = slots_14_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4614 = issue_slots_14_grant ? issue_slots_14_uop_br_tag : _GEN_4515; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [11:0] issue_slots_14_uop_br_mask = slots_14_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] _GEN_4615 = issue_slots_14_grant ? issue_slots_14_uop_br_mask : _GEN_4516; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_sfb = slots_14_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4616 = issue_slots_14_grant ? issue_slots_14_uop_is_sfb : _GEN_4517; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_jal = slots_14_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4617 = issue_slots_14_grant ? issue_slots_14_uop_is_jal : _GEN_4518; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_jalr = slots_14_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4618 = issue_slots_14_grant ? issue_slots_14_uop_is_jalr : _GEN_4519; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_br = slots_14_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4619 = issue_slots_14_grant ? issue_slots_14_uop_is_br : _GEN_4520; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_iw_p2_poisoned = slots_14_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4620 = issue_slots_14_grant ? issue_slots_14_uop_iw_p2_poisoned : _GEN_4521; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_iw_p1_poisoned = slots_14_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4621 = issue_slots_14_grant ? issue_slots_14_uop_iw_p1_poisoned : _GEN_4522; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_iw_state = slots_14_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4622 = issue_slots_14_grant ? issue_slots_14_uop_iw_state : _GEN_4523; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_ctrl_op3_sel = slots_14_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4623 = issue_slots_14_grant ? issue_slots_14_uop_ctrl_op3_sel : _GEN_4524; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_ctrl_is_std = slots_14_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4624 = issue_slots_14_grant ? issue_slots_14_uop_ctrl_is_std : _GEN_4525; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_ctrl_is_sta = slots_14_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4625 = issue_slots_14_grant ? issue_slots_14_uop_ctrl_is_sta : _GEN_4526; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_ctrl_is_load = slots_14_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4626 = issue_slots_14_grant ? issue_slots_14_uop_ctrl_is_load : _GEN_4527; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_14_uop_ctrl_csr_cmd = slots_14_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4627 = issue_slots_14_grant ? issue_slots_14_uop_ctrl_csr_cmd : _GEN_4528; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_ctrl_fcn_dw = slots_14_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4628 = issue_slots_14_grant ? issue_slots_14_uop_ctrl_fcn_dw : _GEN_4529; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_14_uop_ctrl_op_fcn = slots_14_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4629 = issue_slots_14_grant ? issue_slots_14_uop_ctrl_op_fcn : _GEN_4530; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_14_uop_ctrl_imm_sel = slots_14_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4630 = issue_slots_14_grant ? issue_slots_14_uop_ctrl_imm_sel : _GEN_4531; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_14_uop_ctrl_op2_sel = slots_14_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4631 = issue_slots_14_grant ? issue_slots_14_uop_ctrl_op2_sel : _GEN_4532; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_ctrl_op1_sel = slots_14_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4632 = issue_slots_14_grant ? issue_slots_14_uop_ctrl_op1_sel : _GEN_4533; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_14_uop_ctrl_br_type = slots_14_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4633 = issue_slots_14_grant ? issue_slots_14_uop_ctrl_br_type : _GEN_4534; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [9:0] _GEN_4634 = issue_slots_14_grant ? issue_slots_14_uop_fu_code : _GEN_4535; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_14_uop_iq_type = slots_14_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4635 = issue_slots_14_grant ? issue_slots_14_uop_iq_type : _GEN_4536; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [39:0] issue_slots_14_uop_debug_pc = slots_14_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] _GEN_4636 = issue_slots_14_grant ? issue_slots_14_uop_debug_pc : _GEN_4537; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_rvc = slots_14_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4637 = issue_slots_14_grant ? issue_slots_14_uop_is_rvc : _GEN_4538; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_14_uop_debug_inst = slots_14_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4638 = issue_slots_14_grant ? issue_slots_14_uop_debug_inst : _GEN_4539; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [31:0] issue_slots_14_uop_inst = slots_14_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] _GEN_4639 = issue_slots_14_grant ? issue_slots_14_uop_inst : _GEN_4540; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [6:0] issue_slots_14_uop_uopc = slots_14_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] _GEN_4640 = issue_slots_14_grant ? issue_slots_14_uop_uopc : _GEN_4541; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_14_uop_address_num = slots_14_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4641 = issue_slots_14_grant ? issue_slots_14_uop_address_num : _GEN_4542; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_14_uop_rob_inst_idx = slots_14_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4642 = issue_slots_14_grant ? issue_slots_14_uop_rob_inst_idx : _GEN_4543; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_14_uop_self_index = slots_14_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4643 = issue_slots_14_grant ? issue_slots_14_uop_self_index : _GEN_4544; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [5:0] issue_slots_14_uop_split_num = slots_14_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] _GEN_4644 = issue_slots_14_grant ? issue_slots_14_uop_split_num : _GEN_4545; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_14_uop_op2_sel = slots_14_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4645 = issue_slots_14_grant ? issue_slots_14_uop_op2_sel : _GEN_4546; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_14_uop_op1_sel = slots_14_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4646 = issue_slots_14_grant ? issue_slots_14_uop_op1_sel : _GEN_4547; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_14_uop_stale_pflag = slots_14_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4647 = issue_slots_14_grant ? issue_slots_14_uop_stale_pflag : _GEN_4548; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_pflag_busy = slots_14_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4648 = issue_slots_14_grant ? issue_slots_14_uop_pflag_busy : _GEN_4549; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_14_uop_pwflag = slots_14_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4649 = issue_slots_14_grant ? issue_slots_14_uop_pwflag : _GEN_4550; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [3:0] issue_slots_14_uop_prflag = slots_14_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] _GEN_4650 = issue_slots_14_grant ? issue_slots_14_uop_prflag : _GEN_4551; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_wflag = slots_14_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4651 = issue_slots_14_grant ? issue_slots_14_uop_wflag : _GEN_4552; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_rflag = slots_14_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4652 = issue_slots_14_grant ? issue_slots_14_uop_rflag : _GEN_4553; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_14_uop_lrs3_rtype = slots_14_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] _GEN_4653 = issue_slots_14_grant ? issue_slots_14_uop_lrs3_rtype : _GEN_4554; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [2:0] issue_slots_14_uop_shift = slots_14_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] _GEN_4654 = issue_slots_14_grant ? issue_slots_14_uop_shift : _GEN_4555; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_is_unicore = slots_14_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4655 = issue_slots_14_grant ? issue_slots_14_uop_is_unicore : _GEN_4556; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_switch_off = slots_14_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4656 = issue_slots_14_grant ? issue_slots_14_uop_switch_off : _GEN_4557; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire  issue_slots_14_uop_switch = slots_14_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  _GEN_4657 = issue_slots_14_grant ? issue_slots_14_uop_switch : _GEN_4558; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  wire [1:0] issue_slots_15_uop_debug_tsrc = slots_15_io_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_uop_debug_fsrc = slots_15_io_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_bp_xcpt_if = slots_15_io_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_bp_debug_if = slots_15_io_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_xcpt_ma_if = slots_15_io_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_xcpt_ae_if = slots_15_io_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_xcpt_pf_if = slots_15_io_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_fp_single = slots_15_io_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_fp_val = slots_15_io_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_frs3_en = slots_15_io_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_uop_lrs2_rtype = slots_15_io_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_uop_lrs1_rtype = slots_15_io_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_uop_dst_rtype = slots_15_io_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_ldst_val = slots_15_io_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_uop_lrs3 = slots_15_io_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_uop_lrs2 = slots_15_io_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_uop_lrs1 = slots_15_io_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_uop_ldst = slots_15_io_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_ldst_is_rs1 = slots_15_io_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_flush_on_commit = slots_15_io_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_is_unique = slots_15_io_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_is_sys_pc2epc = slots_15_io_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_uses_stq = slots_15_io_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_uses_ldq = slots_15_io_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_is_amo = slots_15_io_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_is_fencei = slots_15_io_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_is_fence = slots_15_io_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_mem_signed = slots_15_io_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_uop_mem_size = slots_15_io_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_15_uop_mem_cmd = slots_15_io_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_bypassable = slots_15_io_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [63:0] issue_slots_15_uop_exc_cause = slots_15_io_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_exception = slots_15_io_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_15_uop_stale_pdst = slots_15_io_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_ppred_busy = slots_15_io_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_prs3_busy = slots_15_io_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_prs2_busy = slots_15_io_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_prs1_busy = slots_15_io_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_15_uop_ppred = slots_15_io_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_15_uop_prs3 = slots_15_io_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_15_uop_prs2 = slots_15_io_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_15_uop_prs1 = slots_15_io_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_15_uop_pdst = slots_15_io_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_uop_rxq_idx = slots_15_io_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_15_uop_stq_idx = slots_15_io_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_15_uop_ldq_idx = slots_15_io_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_uop_rob_idx = slots_15_io_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_15_uop_csr_addr = slots_15_io_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [19:0] issue_slots_15_uop_imm_packed = slots_15_io_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_taken = slots_15_io_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_uop_pc_lob = slots_15_io_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_edge_inst = slots_15_io_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [4:0] issue_slots_15_uop_ftq_idx = slots_15_io_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_uop_br_tag = slots_15_io_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [11:0] issue_slots_15_uop_br_mask = slots_15_io_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_is_sfb = slots_15_io_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_is_jal = slots_15_io_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_is_jalr = slots_15_io_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_is_br = slots_15_io_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_iw_p2_poisoned = slots_15_io_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_iw_p1_poisoned = slots_15_io_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_uop_iw_state = slots_15_io_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_uop_ctrl_op3_sel = slots_15_io_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_ctrl_is_std = slots_15_io_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_ctrl_is_sta = slots_15_io_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_ctrl_is_load = slots_15_io_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_15_uop_ctrl_csr_cmd = slots_15_io_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_ctrl_fcn_dw = slots_15_io_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_uop_ctrl_op_fcn = slots_15_io_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_15_uop_ctrl_imm_sel = slots_15_io_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_15_uop_ctrl_op2_sel = slots_15_io_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_uop_ctrl_op1_sel = slots_15_io_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_uop_ctrl_br_type = slots_15_io_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_15_uop_iq_type = slots_15_io_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [39:0] issue_slots_15_uop_debug_pc = slots_15_io_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_is_rvc = slots_15_io_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_15_uop_debug_inst = slots_15_io_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [31:0] issue_slots_15_uop_inst = slots_15_io_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [6:0] issue_slots_15_uop_uopc = slots_15_io_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_uop_address_num = slots_15_io_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_uop_rob_inst_idx = slots_15_io_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_uop_self_index = slots_15_io_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [5:0] issue_slots_15_uop_split_num = slots_15_io_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_uop_op2_sel = slots_15_io_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_uop_op1_sel = slots_15_io_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_uop_stale_pflag = slots_15_io_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_pflag_busy = slots_15_io_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_uop_pwflag = slots_15_io_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [3:0] issue_slots_15_uop_prflag = slots_15_io_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_wflag = slots_15_io_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_rflag = slots_15_io_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [1:0] issue_slots_15_uop_lrs3_rtype = slots_15_io_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire [2:0] issue_slots_15_uop_shift = slots_15_io_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_is_unicore = slots_15_io_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_switch_off = slots_15_io_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  wire  issue_slots_15_uop_switch = slots_15_io_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 158:28]
  IssueSlot slots_0 ( // @[issue-unit.scala 157:73]
    .clock(slots_0_clock),
    .reset(slots_0_reset),
    .io_valid(slots_0_io_valid),
    .io_will_be_valid(slots_0_io_will_be_valid),
    .io_request(slots_0_io_request),
    .io_request_hp(slots_0_io_request_hp),
    .io_grant(slots_0_io_grant),
    .io_brupdate_b1_resolve_mask(slots_0_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_0_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_0_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_0_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_0_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_0_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_0_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_0_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_0_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_0_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_0_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_0_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_0_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_0_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_0_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_0_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_0_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_0_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_0_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_0_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_0_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_0_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_0_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_0_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_0_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_0_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_0_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_0_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_0_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_0_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_0_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_0_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_0_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_0_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_0_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_0_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_0_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_0_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_0_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_0_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_0_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_0_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_0_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_0_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_0_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_0_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_0_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_0_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_0_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_0_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_0_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_0_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_0_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_0_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_0_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_0_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_0_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_0_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_0_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_0_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_0_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_0_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_0_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_0_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_0_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_0_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_0_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_0_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_0_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_0_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_0_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_0_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_0_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_0_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_0_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_0_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_0_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_0_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_0_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_0_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_0_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_0_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_0_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_0_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_0_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_0_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_0_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_0_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_0_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_0_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_0_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_0_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_0_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_0_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_0_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_0_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_0_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_0_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_0_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_0_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_0_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_0_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_0_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_0_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_0_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_0_io_brupdate_b2_target_offset),
    .io_kill(slots_0_io_kill),
    .io_clear(slots_0_io_clear),
    .io_ldspec_miss(slots_0_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_0_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_0_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_0_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_0_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_0_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_0_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_0_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_0_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_0_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_0_io_wakeup_ports_1_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_0_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_0_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_0_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_0_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_0_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_0_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_0_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_0_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_0_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_0_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_0_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_0_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_0_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_0_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_0_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_0_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_0_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_0_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_0_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_0_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_0_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_0_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_0_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_0_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_0_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_0_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_0_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_0_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_0_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_0_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_0_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_0_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_0_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_0_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_0_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_0_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_0_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_0_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_0_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_0_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_0_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_0_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_0_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_0_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_0_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_0_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_0_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_0_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_0_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_0_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_0_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_0_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_0_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_0_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_0_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_0_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_0_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_0_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_0_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_0_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_0_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_0_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_0_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_0_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_0_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_0_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_0_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_0_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_0_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_0_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_0_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_0_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_0_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_0_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_0_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_0_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_0_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_0_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_0_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_0_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_0_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_0_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_0_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_0_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_0_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_0_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_0_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_0_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_0_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_0_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_0_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_0_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_0_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_0_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_0_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_0_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_0_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_0_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_0_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_0_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_0_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_0_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_0_io_out_uop_switch),
    .io_out_uop_switch_off(slots_0_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_0_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_0_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_0_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_0_io_out_uop_rflag),
    .io_out_uop_wflag(slots_0_io_out_uop_wflag),
    .io_out_uop_prflag(slots_0_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_0_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_0_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_0_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_0_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_0_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_0_io_out_uop_split_num),
    .io_out_uop_self_index(slots_0_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_0_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_0_io_out_uop_address_num),
    .io_out_uop_uopc(slots_0_io_out_uop_uopc),
    .io_out_uop_inst(slots_0_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_0_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_0_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_0_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_0_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_0_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_0_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_0_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_0_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_0_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_0_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_0_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_0_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_0_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_0_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_0_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_0_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_0_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_0_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_0_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_0_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_0_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_0_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_0_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_0_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_0_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_0_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_0_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_0_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_0_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_0_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_0_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_0_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_0_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_0_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_0_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_0_io_out_uop_pdst),
    .io_out_uop_prs1(slots_0_io_out_uop_prs1),
    .io_out_uop_prs2(slots_0_io_out_uop_prs2),
    .io_out_uop_prs3(slots_0_io_out_uop_prs3),
    .io_out_uop_ppred(slots_0_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_0_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_0_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_0_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_0_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_0_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_0_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_0_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_0_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_0_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_0_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_0_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_0_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_0_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_0_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_0_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_0_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_0_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_0_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_0_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_0_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_0_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_0_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_0_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_0_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_0_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_0_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_0_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_0_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_0_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_0_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_0_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_0_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_0_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_0_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_0_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_0_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_0_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_0_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_0_io_uop_switch),
    .io_uop_switch_off(slots_0_io_uop_switch_off),
    .io_uop_is_unicore(slots_0_io_uop_is_unicore),
    .io_uop_shift(slots_0_io_uop_shift),
    .io_uop_lrs3_rtype(slots_0_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_0_io_uop_rflag),
    .io_uop_wflag(slots_0_io_uop_wflag),
    .io_uop_prflag(slots_0_io_uop_prflag),
    .io_uop_pwflag(slots_0_io_uop_pwflag),
    .io_uop_pflag_busy(slots_0_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_0_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_0_io_uop_op1_sel),
    .io_uop_op2_sel(slots_0_io_uop_op2_sel),
    .io_uop_split_num(slots_0_io_uop_split_num),
    .io_uop_self_index(slots_0_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_0_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_0_io_uop_address_num),
    .io_uop_uopc(slots_0_io_uop_uopc),
    .io_uop_inst(slots_0_io_uop_inst),
    .io_uop_debug_inst(slots_0_io_uop_debug_inst),
    .io_uop_is_rvc(slots_0_io_uop_is_rvc),
    .io_uop_debug_pc(slots_0_io_uop_debug_pc),
    .io_uop_iq_type(slots_0_io_uop_iq_type),
    .io_uop_fu_code(slots_0_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_0_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_0_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_0_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_0_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_0_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_0_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_0_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_0_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_0_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_0_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_0_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_0_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_0_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_0_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_0_io_uop_is_br),
    .io_uop_is_jalr(slots_0_io_uop_is_jalr),
    .io_uop_is_jal(slots_0_io_uop_is_jal),
    .io_uop_is_sfb(slots_0_io_uop_is_sfb),
    .io_uop_br_mask(slots_0_io_uop_br_mask),
    .io_uop_br_tag(slots_0_io_uop_br_tag),
    .io_uop_ftq_idx(slots_0_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_0_io_uop_edge_inst),
    .io_uop_pc_lob(slots_0_io_uop_pc_lob),
    .io_uop_taken(slots_0_io_uop_taken),
    .io_uop_imm_packed(slots_0_io_uop_imm_packed),
    .io_uop_csr_addr(slots_0_io_uop_csr_addr),
    .io_uop_rob_idx(slots_0_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_0_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_0_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_0_io_uop_rxq_idx),
    .io_uop_pdst(slots_0_io_uop_pdst),
    .io_uop_prs1(slots_0_io_uop_prs1),
    .io_uop_prs2(slots_0_io_uop_prs2),
    .io_uop_prs3(slots_0_io_uop_prs3),
    .io_uop_ppred(slots_0_io_uop_ppred),
    .io_uop_prs1_busy(slots_0_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_0_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_0_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_0_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_0_io_uop_stale_pdst),
    .io_uop_exception(slots_0_io_uop_exception),
    .io_uop_exc_cause(slots_0_io_uop_exc_cause),
    .io_uop_bypassable(slots_0_io_uop_bypassable),
    .io_uop_mem_cmd(slots_0_io_uop_mem_cmd),
    .io_uop_mem_size(slots_0_io_uop_mem_size),
    .io_uop_mem_signed(slots_0_io_uop_mem_signed),
    .io_uop_is_fence(slots_0_io_uop_is_fence),
    .io_uop_is_fencei(slots_0_io_uop_is_fencei),
    .io_uop_is_amo(slots_0_io_uop_is_amo),
    .io_uop_uses_ldq(slots_0_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_0_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_0_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_0_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_0_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_0_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_0_io_uop_ldst),
    .io_uop_lrs1(slots_0_io_uop_lrs1),
    .io_uop_lrs2(slots_0_io_uop_lrs2),
    .io_uop_lrs3(slots_0_io_uop_lrs3),
    .io_uop_ldst_val(slots_0_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_0_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_0_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_0_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_0_io_uop_frs3_en),
    .io_uop_fp_val(slots_0_io_uop_fp_val),
    .io_uop_fp_single(slots_0_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_0_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_0_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_0_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_0_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_0_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_0_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_0_io_uop_debug_tsrc),
    .io_debug_p1(slots_0_io_debug_p1),
    .io_debug_p2(slots_0_io_debug_p2),
    .io_debug_p3(slots_0_io_debug_p3),
    .io_debug_ppred(slots_0_io_debug_ppred),
    .io_debug_state(slots_0_io_debug_state)
  );
  IssueSlot slots_1 ( // @[issue-unit.scala 157:73]
    .clock(slots_1_clock),
    .reset(slots_1_reset),
    .io_valid(slots_1_io_valid),
    .io_will_be_valid(slots_1_io_will_be_valid),
    .io_request(slots_1_io_request),
    .io_request_hp(slots_1_io_request_hp),
    .io_grant(slots_1_io_grant),
    .io_brupdate_b1_resolve_mask(slots_1_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_1_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_1_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_1_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_1_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_1_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_1_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_1_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_1_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_1_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_1_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_1_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_1_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_1_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_1_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_1_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_1_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_1_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_1_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_1_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_1_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_1_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_1_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_1_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_1_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_1_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_1_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_1_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_1_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_1_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_1_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_1_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_1_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_1_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_1_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_1_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_1_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_1_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_1_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_1_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_1_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_1_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_1_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_1_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_1_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_1_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_1_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_1_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_1_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_1_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_1_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_1_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_1_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_1_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_1_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_1_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_1_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_1_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_1_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_1_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_1_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_1_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_1_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_1_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_1_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_1_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_1_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_1_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_1_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_1_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_1_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_1_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_1_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_1_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_1_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_1_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_1_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_1_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_1_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_1_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_1_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_1_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_1_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_1_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_1_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_1_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_1_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_1_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_1_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_1_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_1_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_1_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_1_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_1_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_1_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_1_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_1_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_1_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_1_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_1_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_1_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_1_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_1_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_1_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_1_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_1_io_brupdate_b2_target_offset),
    .io_kill(slots_1_io_kill),
    .io_clear(slots_1_io_clear),
    .io_ldspec_miss(slots_1_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_1_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_1_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_1_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_1_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_1_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_1_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_1_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_1_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_1_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_1_io_wakeup_ports_1_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_1_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_1_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_1_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_1_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_1_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_1_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_1_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_1_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_1_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_1_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_1_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_1_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_1_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_1_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_1_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_1_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_1_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_1_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_1_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_1_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_1_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_1_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_1_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_1_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_1_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_1_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_1_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_1_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_1_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_1_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_1_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_1_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_1_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_1_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_1_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_1_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_1_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_1_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_1_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_1_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_1_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_1_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_1_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_1_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_1_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_1_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_1_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_1_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_1_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_1_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_1_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_1_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_1_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_1_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_1_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_1_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_1_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_1_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_1_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_1_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_1_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_1_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_1_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_1_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_1_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_1_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_1_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_1_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_1_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_1_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_1_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_1_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_1_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_1_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_1_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_1_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_1_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_1_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_1_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_1_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_1_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_1_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_1_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_1_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_1_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_1_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_1_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_1_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_1_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_1_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_1_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_1_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_1_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_1_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_1_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_1_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_1_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_1_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_1_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_1_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_1_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_1_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_1_io_out_uop_switch),
    .io_out_uop_switch_off(slots_1_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_1_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_1_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_1_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_1_io_out_uop_rflag),
    .io_out_uop_wflag(slots_1_io_out_uop_wflag),
    .io_out_uop_prflag(slots_1_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_1_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_1_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_1_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_1_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_1_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_1_io_out_uop_split_num),
    .io_out_uop_self_index(slots_1_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_1_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_1_io_out_uop_address_num),
    .io_out_uop_uopc(slots_1_io_out_uop_uopc),
    .io_out_uop_inst(slots_1_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_1_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_1_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_1_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_1_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_1_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_1_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_1_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_1_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_1_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_1_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_1_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_1_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_1_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_1_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_1_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_1_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_1_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_1_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_1_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_1_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_1_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_1_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_1_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_1_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_1_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_1_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_1_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_1_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_1_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_1_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_1_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_1_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_1_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_1_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_1_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_1_io_out_uop_pdst),
    .io_out_uop_prs1(slots_1_io_out_uop_prs1),
    .io_out_uop_prs2(slots_1_io_out_uop_prs2),
    .io_out_uop_prs3(slots_1_io_out_uop_prs3),
    .io_out_uop_ppred(slots_1_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_1_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_1_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_1_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_1_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_1_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_1_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_1_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_1_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_1_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_1_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_1_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_1_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_1_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_1_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_1_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_1_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_1_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_1_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_1_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_1_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_1_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_1_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_1_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_1_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_1_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_1_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_1_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_1_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_1_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_1_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_1_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_1_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_1_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_1_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_1_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_1_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_1_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_1_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_1_io_uop_switch),
    .io_uop_switch_off(slots_1_io_uop_switch_off),
    .io_uop_is_unicore(slots_1_io_uop_is_unicore),
    .io_uop_shift(slots_1_io_uop_shift),
    .io_uop_lrs3_rtype(slots_1_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_1_io_uop_rflag),
    .io_uop_wflag(slots_1_io_uop_wflag),
    .io_uop_prflag(slots_1_io_uop_prflag),
    .io_uop_pwflag(slots_1_io_uop_pwflag),
    .io_uop_pflag_busy(slots_1_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_1_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_1_io_uop_op1_sel),
    .io_uop_op2_sel(slots_1_io_uop_op2_sel),
    .io_uop_split_num(slots_1_io_uop_split_num),
    .io_uop_self_index(slots_1_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_1_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_1_io_uop_address_num),
    .io_uop_uopc(slots_1_io_uop_uopc),
    .io_uop_inst(slots_1_io_uop_inst),
    .io_uop_debug_inst(slots_1_io_uop_debug_inst),
    .io_uop_is_rvc(slots_1_io_uop_is_rvc),
    .io_uop_debug_pc(slots_1_io_uop_debug_pc),
    .io_uop_iq_type(slots_1_io_uop_iq_type),
    .io_uop_fu_code(slots_1_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_1_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_1_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_1_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_1_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_1_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_1_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_1_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_1_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_1_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_1_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_1_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_1_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_1_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_1_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_1_io_uop_is_br),
    .io_uop_is_jalr(slots_1_io_uop_is_jalr),
    .io_uop_is_jal(slots_1_io_uop_is_jal),
    .io_uop_is_sfb(slots_1_io_uop_is_sfb),
    .io_uop_br_mask(slots_1_io_uop_br_mask),
    .io_uop_br_tag(slots_1_io_uop_br_tag),
    .io_uop_ftq_idx(slots_1_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_1_io_uop_edge_inst),
    .io_uop_pc_lob(slots_1_io_uop_pc_lob),
    .io_uop_taken(slots_1_io_uop_taken),
    .io_uop_imm_packed(slots_1_io_uop_imm_packed),
    .io_uop_csr_addr(slots_1_io_uop_csr_addr),
    .io_uop_rob_idx(slots_1_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_1_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_1_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_1_io_uop_rxq_idx),
    .io_uop_pdst(slots_1_io_uop_pdst),
    .io_uop_prs1(slots_1_io_uop_prs1),
    .io_uop_prs2(slots_1_io_uop_prs2),
    .io_uop_prs3(slots_1_io_uop_prs3),
    .io_uop_ppred(slots_1_io_uop_ppred),
    .io_uop_prs1_busy(slots_1_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_1_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_1_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_1_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_1_io_uop_stale_pdst),
    .io_uop_exception(slots_1_io_uop_exception),
    .io_uop_exc_cause(slots_1_io_uop_exc_cause),
    .io_uop_bypassable(slots_1_io_uop_bypassable),
    .io_uop_mem_cmd(slots_1_io_uop_mem_cmd),
    .io_uop_mem_size(slots_1_io_uop_mem_size),
    .io_uop_mem_signed(slots_1_io_uop_mem_signed),
    .io_uop_is_fence(slots_1_io_uop_is_fence),
    .io_uop_is_fencei(slots_1_io_uop_is_fencei),
    .io_uop_is_amo(slots_1_io_uop_is_amo),
    .io_uop_uses_ldq(slots_1_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_1_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_1_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_1_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_1_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_1_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_1_io_uop_ldst),
    .io_uop_lrs1(slots_1_io_uop_lrs1),
    .io_uop_lrs2(slots_1_io_uop_lrs2),
    .io_uop_lrs3(slots_1_io_uop_lrs3),
    .io_uop_ldst_val(slots_1_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_1_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_1_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_1_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_1_io_uop_frs3_en),
    .io_uop_fp_val(slots_1_io_uop_fp_val),
    .io_uop_fp_single(slots_1_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_1_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_1_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_1_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_1_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_1_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_1_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_1_io_uop_debug_tsrc),
    .io_debug_p1(slots_1_io_debug_p1),
    .io_debug_p2(slots_1_io_debug_p2),
    .io_debug_p3(slots_1_io_debug_p3),
    .io_debug_ppred(slots_1_io_debug_ppred),
    .io_debug_state(slots_1_io_debug_state)
  );
  IssueSlot slots_2 ( // @[issue-unit.scala 157:73]
    .clock(slots_2_clock),
    .reset(slots_2_reset),
    .io_valid(slots_2_io_valid),
    .io_will_be_valid(slots_2_io_will_be_valid),
    .io_request(slots_2_io_request),
    .io_request_hp(slots_2_io_request_hp),
    .io_grant(slots_2_io_grant),
    .io_brupdate_b1_resolve_mask(slots_2_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_2_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_2_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_2_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_2_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_2_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_2_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_2_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_2_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_2_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_2_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_2_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_2_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_2_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_2_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_2_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_2_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_2_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_2_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_2_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_2_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_2_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_2_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_2_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_2_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_2_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_2_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_2_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_2_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_2_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_2_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_2_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_2_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_2_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_2_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_2_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_2_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_2_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_2_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_2_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_2_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_2_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_2_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_2_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_2_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_2_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_2_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_2_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_2_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_2_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_2_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_2_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_2_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_2_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_2_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_2_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_2_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_2_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_2_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_2_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_2_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_2_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_2_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_2_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_2_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_2_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_2_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_2_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_2_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_2_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_2_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_2_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_2_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_2_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_2_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_2_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_2_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_2_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_2_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_2_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_2_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_2_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_2_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_2_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_2_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_2_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_2_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_2_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_2_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_2_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_2_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_2_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_2_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_2_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_2_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_2_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_2_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_2_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_2_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_2_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_2_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_2_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_2_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_2_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_2_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_2_io_brupdate_b2_target_offset),
    .io_kill(slots_2_io_kill),
    .io_clear(slots_2_io_clear),
    .io_ldspec_miss(slots_2_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_2_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_2_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_2_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_2_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_2_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_2_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_2_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_2_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_2_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_2_io_wakeup_ports_1_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_2_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_2_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_2_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_2_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_2_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_2_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_2_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_2_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_2_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_2_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_2_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_2_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_2_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_2_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_2_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_2_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_2_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_2_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_2_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_2_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_2_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_2_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_2_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_2_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_2_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_2_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_2_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_2_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_2_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_2_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_2_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_2_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_2_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_2_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_2_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_2_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_2_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_2_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_2_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_2_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_2_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_2_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_2_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_2_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_2_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_2_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_2_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_2_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_2_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_2_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_2_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_2_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_2_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_2_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_2_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_2_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_2_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_2_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_2_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_2_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_2_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_2_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_2_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_2_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_2_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_2_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_2_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_2_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_2_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_2_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_2_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_2_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_2_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_2_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_2_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_2_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_2_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_2_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_2_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_2_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_2_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_2_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_2_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_2_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_2_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_2_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_2_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_2_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_2_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_2_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_2_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_2_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_2_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_2_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_2_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_2_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_2_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_2_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_2_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_2_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_2_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_2_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_2_io_out_uop_switch),
    .io_out_uop_switch_off(slots_2_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_2_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_2_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_2_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_2_io_out_uop_rflag),
    .io_out_uop_wflag(slots_2_io_out_uop_wflag),
    .io_out_uop_prflag(slots_2_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_2_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_2_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_2_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_2_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_2_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_2_io_out_uop_split_num),
    .io_out_uop_self_index(slots_2_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_2_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_2_io_out_uop_address_num),
    .io_out_uop_uopc(slots_2_io_out_uop_uopc),
    .io_out_uop_inst(slots_2_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_2_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_2_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_2_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_2_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_2_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_2_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_2_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_2_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_2_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_2_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_2_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_2_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_2_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_2_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_2_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_2_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_2_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_2_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_2_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_2_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_2_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_2_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_2_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_2_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_2_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_2_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_2_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_2_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_2_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_2_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_2_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_2_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_2_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_2_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_2_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_2_io_out_uop_pdst),
    .io_out_uop_prs1(slots_2_io_out_uop_prs1),
    .io_out_uop_prs2(slots_2_io_out_uop_prs2),
    .io_out_uop_prs3(slots_2_io_out_uop_prs3),
    .io_out_uop_ppred(slots_2_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_2_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_2_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_2_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_2_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_2_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_2_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_2_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_2_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_2_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_2_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_2_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_2_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_2_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_2_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_2_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_2_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_2_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_2_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_2_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_2_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_2_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_2_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_2_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_2_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_2_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_2_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_2_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_2_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_2_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_2_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_2_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_2_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_2_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_2_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_2_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_2_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_2_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_2_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_2_io_uop_switch),
    .io_uop_switch_off(slots_2_io_uop_switch_off),
    .io_uop_is_unicore(slots_2_io_uop_is_unicore),
    .io_uop_shift(slots_2_io_uop_shift),
    .io_uop_lrs3_rtype(slots_2_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_2_io_uop_rflag),
    .io_uop_wflag(slots_2_io_uop_wflag),
    .io_uop_prflag(slots_2_io_uop_prflag),
    .io_uop_pwflag(slots_2_io_uop_pwflag),
    .io_uop_pflag_busy(slots_2_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_2_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_2_io_uop_op1_sel),
    .io_uop_op2_sel(slots_2_io_uop_op2_sel),
    .io_uop_split_num(slots_2_io_uop_split_num),
    .io_uop_self_index(slots_2_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_2_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_2_io_uop_address_num),
    .io_uop_uopc(slots_2_io_uop_uopc),
    .io_uop_inst(slots_2_io_uop_inst),
    .io_uop_debug_inst(slots_2_io_uop_debug_inst),
    .io_uop_is_rvc(slots_2_io_uop_is_rvc),
    .io_uop_debug_pc(slots_2_io_uop_debug_pc),
    .io_uop_iq_type(slots_2_io_uop_iq_type),
    .io_uop_fu_code(slots_2_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_2_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_2_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_2_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_2_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_2_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_2_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_2_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_2_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_2_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_2_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_2_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_2_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_2_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_2_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_2_io_uop_is_br),
    .io_uop_is_jalr(slots_2_io_uop_is_jalr),
    .io_uop_is_jal(slots_2_io_uop_is_jal),
    .io_uop_is_sfb(slots_2_io_uop_is_sfb),
    .io_uop_br_mask(slots_2_io_uop_br_mask),
    .io_uop_br_tag(slots_2_io_uop_br_tag),
    .io_uop_ftq_idx(slots_2_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_2_io_uop_edge_inst),
    .io_uop_pc_lob(slots_2_io_uop_pc_lob),
    .io_uop_taken(slots_2_io_uop_taken),
    .io_uop_imm_packed(slots_2_io_uop_imm_packed),
    .io_uop_csr_addr(slots_2_io_uop_csr_addr),
    .io_uop_rob_idx(slots_2_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_2_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_2_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_2_io_uop_rxq_idx),
    .io_uop_pdst(slots_2_io_uop_pdst),
    .io_uop_prs1(slots_2_io_uop_prs1),
    .io_uop_prs2(slots_2_io_uop_prs2),
    .io_uop_prs3(slots_2_io_uop_prs3),
    .io_uop_ppred(slots_2_io_uop_ppred),
    .io_uop_prs1_busy(slots_2_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_2_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_2_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_2_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_2_io_uop_stale_pdst),
    .io_uop_exception(slots_2_io_uop_exception),
    .io_uop_exc_cause(slots_2_io_uop_exc_cause),
    .io_uop_bypassable(slots_2_io_uop_bypassable),
    .io_uop_mem_cmd(slots_2_io_uop_mem_cmd),
    .io_uop_mem_size(slots_2_io_uop_mem_size),
    .io_uop_mem_signed(slots_2_io_uop_mem_signed),
    .io_uop_is_fence(slots_2_io_uop_is_fence),
    .io_uop_is_fencei(slots_2_io_uop_is_fencei),
    .io_uop_is_amo(slots_2_io_uop_is_amo),
    .io_uop_uses_ldq(slots_2_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_2_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_2_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_2_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_2_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_2_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_2_io_uop_ldst),
    .io_uop_lrs1(slots_2_io_uop_lrs1),
    .io_uop_lrs2(slots_2_io_uop_lrs2),
    .io_uop_lrs3(slots_2_io_uop_lrs3),
    .io_uop_ldst_val(slots_2_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_2_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_2_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_2_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_2_io_uop_frs3_en),
    .io_uop_fp_val(slots_2_io_uop_fp_val),
    .io_uop_fp_single(slots_2_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_2_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_2_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_2_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_2_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_2_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_2_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_2_io_uop_debug_tsrc),
    .io_debug_p1(slots_2_io_debug_p1),
    .io_debug_p2(slots_2_io_debug_p2),
    .io_debug_p3(slots_2_io_debug_p3),
    .io_debug_ppred(slots_2_io_debug_ppred),
    .io_debug_state(slots_2_io_debug_state)
  );
  IssueSlot slots_3 ( // @[issue-unit.scala 157:73]
    .clock(slots_3_clock),
    .reset(slots_3_reset),
    .io_valid(slots_3_io_valid),
    .io_will_be_valid(slots_3_io_will_be_valid),
    .io_request(slots_3_io_request),
    .io_request_hp(slots_3_io_request_hp),
    .io_grant(slots_3_io_grant),
    .io_brupdate_b1_resolve_mask(slots_3_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_3_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_3_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_3_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_3_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_3_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_3_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_3_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_3_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_3_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_3_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_3_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_3_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_3_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_3_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_3_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_3_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_3_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_3_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_3_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_3_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_3_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_3_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_3_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_3_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_3_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_3_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_3_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_3_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_3_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_3_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_3_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_3_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_3_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_3_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_3_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_3_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_3_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_3_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_3_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_3_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_3_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_3_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_3_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_3_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_3_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_3_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_3_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_3_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_3_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_3_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_3_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_3_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_3_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_3_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_3_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_3_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_3_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_3_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_3_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_3_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_3_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_3_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_3_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_3_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_3_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_3_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_3_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_3_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_3_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_3_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_3_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_3_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_3_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_3_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_3_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_3_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_3_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_3_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_3_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_3_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_3_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_3_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_3_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_3_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_3_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_3_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_3_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_3_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_3_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_3_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_3_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_3_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_3_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_3_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_3_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_3_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_3_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_3_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_3_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_3_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_3_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_3_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_3_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_3_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_3_io_brupdate_b2_target_offset),
    .io_kill(slots_3_io_kill),
    .io_clear(slots_3_io_clear),
    .io_ldspec_miss(slots_3_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_3_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_3_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_3_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_3_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_3_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_3_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_3_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_3_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_3_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_3_io_wakeup_ports_1_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_3_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_3_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_3_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_3_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_3_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_3_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_3_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_3_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_3_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_3_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_3_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_3_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_3_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_3_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_3_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_3_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_3_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_3_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_3_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_3_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_3_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_3_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_3_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_3_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_3_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_3_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_3_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_3_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_3_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_3_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_3_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_3_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_3_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_3_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_3_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_3_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_3_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_3_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_3_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_3_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_3_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_3_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_3_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_3_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_3_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_3_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_3_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_3_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_3_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_3_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_3_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_3_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_3_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_3_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_3_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_3_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_3_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_3_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_3_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_3_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_3_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_3_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_3_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_3_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_3_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_3_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_3_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_3_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_3_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_3_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_3_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_3_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_3_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_3_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_3_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_3_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_3_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_3_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_3_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_3_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_3_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_3_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_3_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_3_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_3_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_3_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_3_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_3_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_3_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_3_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_3_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_3_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_3_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_3_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_3_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_3_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_3_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_3_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_3_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_3_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_3_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_3_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_3_io_out_uop_switch),
    .io_out_uop_switch_off(slots_3_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_3_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_3_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_3_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_3_io_out_uop_rflag),
    .io_out_uop_wflag(slots_3_io_out_uop_wflag),
    .io_out_uop_prflag(slots_3_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_3_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_3_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_3_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_3_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_3_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_3_io_out_uop_split_num),
    .io_out_uop_self_index(slots_3_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_3_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_3_io_out_uop_address_num),
    .io_out_uop_uopc(slots_3_io_out_uop_uopc),
    .io_out_uop_inst(slots_3_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_3_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_3_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_3_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_3_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_3_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_3_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_3_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_3_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_3_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_3_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_3_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_3_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_3_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_3_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_3_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_3_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_3_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_3_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_3_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_3_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_3_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_3_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_3_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_3_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_3_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_3_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_3_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_3_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_3_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_3_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_3_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_3_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_3_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_3_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_3_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_3_io_out_uop_pdst),
    .io_out_uop_prs1(slots_3_io_out_uop_prs1),
    .io_out_uop_prs2(slots_3_io_out_uop_prs2),
    .io_out_uop_prs3(slots_3_io_out_uop_prs3),
    .io_out_uop_ppred(slots_3_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_3_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_3_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_3_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_3_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_3_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_3_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_3_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_3_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_3_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_3_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_3_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_3_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_3_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_3_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_3_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_3_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_3_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_3_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_3_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_3_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_3_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_3_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_3_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_3_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_3_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_3_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_3_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_3_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_3_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_3_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_3_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_3_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_3_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_3_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_3_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_3_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_3_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_3_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_3_io_uop_switch),
    .io_uop_switch_off(slots_3_io_uop_switch_off),
    .io_uop_is_unicore(slots_3_io_uop_is_unicore),
    .io_uop_shift(slots_3_io_uop_shift),
    .io_uop_lrs3_rtype(slots_3_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_3_io_uop_rflag),
    .io_uop_wflag(slots_3_io_uop_wflag),
    .io_uop_prflag(slots_3_io_uop_prflag),
    .io_uop_pwflag(slots_3_io_uop_pwflag),
    .io_uop_pflag_busy(slots_3_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_3_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_3_io_uop_op1_sel),
    .io_uop_op2_sel(slots_3_io_uop_op2_sel),
    .io_uop_split_num(slots_3_io_uop_split_num),
    .io_uop_self_index(slots_3_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_3_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_3_io_uop_address_num),
    .io_uop_uopc(slots_3_io_uop_uopc),
    .io_uop_inst(slots_3_io_uop_inst),
    .io_uop_debug_inst(slots_3_io_uop_debug_inst),
    .io_uop_is_rvc(slots_3_io_uop_is_rvc),
    .io_uop_debug_pc(slots_3_io_uop_debug_pc),
    .io_uop_iq_type(slots_3_io_uop_iq_type),
    .io_uop_fu_code(slots_3_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_3_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_3_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_3_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_3_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_3_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_3_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_3_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_3_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_3_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_3_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_3_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_3_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_3_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_3_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_3_io_uop_is_br),
    .io_uop_is_jalr(slots_3_io_uop_is_jalr),
    .io_uop_is_jal(slots_3_io_uop_is_jal),
    .io_uop_is_sfb(slots_3_io_uop_is_sfb),
    .io_uop_br_mask(slots_3_io_uop_br_mask),
    .io_uop_br_tag(slots_3_io_uop_br_tag),
    .io_uop_ftq_idx(slots_3_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_3_io_uop_edge_inst),
    .io_uop_pc_lob(slots_3_io_uop_pc_lob),
    .io_uop_taken(slots_3_io_uop_taken),
    .io_uop_imm_packed(slots_3_io_uop_imm_packed),
    .io_uop_csr_addr(slots_3_io_uop_csr_addr),
    .io_uop_rob_idx(slots_3_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_3_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_3_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_3_io_uop_rxq_idx),
    .io_uop_pdst(slots_3_io_uop_pdst),
    .io_uop_prs1(slots_3_io_uop_prs1),
    .io_uop_prs2(slots_3_io_uop_prs2),
    .io_uop_prs3(slots_3_io_uop_prs3),
    .io_uop_ppred(slots_3_io_uop_ppred),
    .io_uop_prs1_busy(slots_3_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_3_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_3_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_3_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_3_io_uop_stale_pdst),
    .io_uop_exception(slots_3_io_uop_exception),
    .io_uop_exc_cause(slots_3_io_uop_exc_cause),
    .io_uop_bypassable(slots_3_io_uop_bypassable),
    .io_uop_mem_cmd(slots_3_io_uop_mem_cmd),
    .io_uop_mem_size(slots_3_io_uop_mem_size),
    .io_uop_mem_signed(slots_3_io_uop_mem_signed),
    .io_uop_is_fence(slots_3_io_uop_is_fence),
    .io_uop_is_fencei(slots_3_io_uop_is_fencei),
    .io_uop_is_amo(slots_3_io_uop_is_amo),
    .io_uop_uses_ldq(slots_3_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_3_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_3_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_3_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_3_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_3_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_3_io_uop_ldst),
    .io_uop_lrs1(slots_3_io_uop_lrs1),
    .io_uop_lrs2(slots_3_io_uop_lrs2),
    .io_uop_lrs3(slots_3_io_uop_lrs3),
    .io_uop_ldst_val(slots_3_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_3_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_3_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_3_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_3_io_uop_frs3_en),
    .io_uop_fp_val(slots_3_io_uop_fp_val),
    .io_uop_fp_single(slots_3_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_3_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_3_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_3_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_3_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_3_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_3_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_3_io_uop_debug_tsrc),
    .io_debug_p1(slots_3_io_debug_p1),
    .io_debug_p2(slots_3_io_debug_p2),
    .io_debug_p3(slots_3_io_debug_p3),
    .io_debug_ppred(slots_3_io_debug_ppred),
    .io_debug_state(slots_3_io_debug_state)
  );
  IssueSlot slots_4 ( // @[issue-unit.scala 157:73]
    .clock(slots_4_clock),
    .reset(slots_4_reset),
    .io_valid(slots_4_io_valid),
    .io_will_be_valid(slots_4_io_will_be_valid),
    .io_request(slots_4_io_request),
    .io_request_hp(slots_4_io_request_hp),
    .io_grant(slots_4_io_grant),
    .io_brupdate_b1_resolve_mask(slots_4_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_4_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_4_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_4_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_4_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_4_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_4_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_4_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_4_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_4_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_4_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_4_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_4_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_4_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_4_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_4_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_4_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_4_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_4_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_4_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_4_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_4_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_4_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_4_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_4_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_4_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_4_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_4_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_4_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_4_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_4_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_4_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_4_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_4_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_4_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_4_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_4_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_4_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_4_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_4_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_4_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_4_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_4_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_4_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_4_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_4_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_4_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_4_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_4_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_4_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_4_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_4_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_4_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_4_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_4_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_4_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_4_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_4_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_4_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_4_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_4_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_4_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_4_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_4_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_4_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_4_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_4_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_4_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_4_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_4_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_4_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_4_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_4_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_4_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_4_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_4_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_4_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_4_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_4_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_4_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_4_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_4_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_4_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_4_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_4_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_4_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_4_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_4_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_4_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_4_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_4_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_4_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_4_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_4_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_4_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_4_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_4_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_4_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_4_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_4_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_4_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_4_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_4_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_4_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_4_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_4_io_brupdate_b2_target_offset),
    .io_kill(slots_4_io_kill),
    .io_clear(slots_4_io_clear),
    .io_ldspec_miss(slots_4_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_4_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_4_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_4_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_4_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_4_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_4_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_4_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_4_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_4_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_4_io_wakeup_ports_1_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_4_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_4_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_4_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_4_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_4_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_4_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_4_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_4_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_4_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_4_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_4_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_4_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_4_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_4_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_4_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_4_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_4_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_4_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_4_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_4_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_4_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_4_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_4_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_4_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_4_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_4_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_4_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_4_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_4_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_4_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_4_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_4_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_4_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_4_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_4_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_4_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_4_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_4_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_4_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_4_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_4_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_4_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_4_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_4_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_4_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_4_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_4_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_4_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_4_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_4_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_4_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_4_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_4_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_4_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_4_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_4_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_4_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_4_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_4_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_4_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_4_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_4_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_4_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_4_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_4_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_4_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_4_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_4_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_4_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_4_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_4_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_4_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_4_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_4_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_4_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_4_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_4_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_4_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_4_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_4_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_4_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_4_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_4_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_4_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_4_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_4_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_4_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_4_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_4_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_4_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_4_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_4_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_4_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_4_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_4_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_4_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_4_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_4_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_4_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_4_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_4_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_4_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_4_io_out_uop_switch),
    .io_out_uop_switch_off(slots_4_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_4_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_4_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_4_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_4_io_out_uop_rflag),
    .io_out_uop_wflag(slots_4_io_out_uop_wflag),
    .io_out_uop_prflag(slots_4_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_4_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_4_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_4_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_4_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_4_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_4_io_out_uop_split_num),
    .io_out_uop_self_index(slots_4_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_4_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_4_io_out_uop_address_num),
    .io_out_uop_uopc(slots_4_io_out_uop_uopc),
    .io_out_uop_inst(slots_4_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_4_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_4_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_4_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_4_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_4_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_4_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_4_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_4_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_4_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_4_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_4_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_4_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_4_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_4_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_4_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_4_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_4_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_4_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_4_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_4_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_4_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_4_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_4_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_4_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_4_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_4_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_4_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_4_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_4_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_4_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_4_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_4_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_4_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_4_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_4_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_4_io_out_uop_pdst),
    .io_out_uop_prs1(slots_4_io_out_uop_prs1),
    .io_out_uop_prs2(slots_4_io_out_uop_prs2),
    .io_out_uop_prs3(slots_4_io_out_uop_prs3),
    .io_out_uop_ppred(slots_4_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_4_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_4_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_4_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_4_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_4_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_4_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_4_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_4_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_4_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_4_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_4_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_4_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_4_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_4_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_4_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_4_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_4_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_4_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_4_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_4_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_4_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_4_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_4_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_4_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_4_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_4_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_4_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_4_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_4_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_4_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_4_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_4_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_4_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_4_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_4_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_4_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_4_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_4_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_4_io_uop_switch),
    .io_uop_switch_off(slots_4_io_uop_switch_off),
    .io_uop_is_unicore(slots_4_io_uop_is_unicore),
    .io_uop_shift(slots_4_io_uop_shift),
    .io_uop_lrs3_rtype(slots_4_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_4_io_uop_rflag),
    .io_uop_wflag(slots_4_io_uop_wflag),
    .io_uop_prflag(slots_4_io_uop_prflag),
    .io_uop_pwflag(slots_4_io_uop_pwflag),
    .io_uop_pflag_busy(slots_4_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_4_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_4_io_uop_op1_sel),
    .io_uop_op2_sel(slots_4_io_uop_op2_sel),
    .io_uop_split_num(slots_4_io_uop_split_num),
    .io_uop_self_index(slots_4_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_4_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_4_io_uop_address_num),
    .io_uop_uopc(slots_4_io_uop_uopc),
    .io_uop_inst(slots_4_io_uop_inst),
    .io_uop_debug_inst(slots_4_io_uop_debug_inst),
    .io_uop_is_rvc(slots_4_io_uop_is_rvc),
    .io_uop_debug_pc(slots_4_io_uop_debug_pc),
    .io_uop_iq_type(slots_4_io_uop_iq_type),
    .io_uop_fu_code(slots_4_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_4_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_4_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_4_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_4_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_4_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_4_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_4_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_4_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_4_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_4_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_4_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_4_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_4_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_4_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_4_io_uop_is_br),
    .io_uop_is_jalr(slots_4_io_uop_is_jalr),
    .io_uop_is_jal(slots_4_io_uop_is_jal),
    .io_uop_is_sfb(slots_4_io_uop_is_sfb),
    .io_uop_br_mask(slots_4_io_uop_br_mask),
    .io_uop_br_tag(slots_4_io_uop_br_tag),
    .io_uop_ftq_idx(slots_4_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_4_io_uop_edge_inst),
    .io_uop_pc_lob(slots_4_io_uop_pc_lob),
    .io_uop_taken(slots_4_io_uop_taken),
    .io_uop_imm_packed(slots_4_io_uop_imm_packed),
    .io_uop_csr_addr(slots_4_io_uop_csr_addr),
    .io_uop_rob_idx(slots_4_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_4_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_4_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_4_io_uop_rxq_idx),
    .io_uop_pdst(slots_4_io_uop_pdst),
    .io_uop_prs1(slots_4_io_uop_prs1),
    .io_uop_prs2(slots_4_io_uop_prs2),
    .io_uop_prs3(slots_4_io_uop_prs3),
    .io_uop_ppred(slots_4_io_uop_ppred),
    .io_uop_prs1_busy(slots_4_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_4_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_4_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_4_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_4_io_uop_stale_pdst),
    .io_uop_exception(slots_4_io_uop_exception),
    .io_uop_exc_cause(slots_4_io_uop_exc_cause),
    .io_uop_bypassable(slots_4_io_uop_bypassable),
    .io_uop_mem_cmd(slots_4_io_uop_mem_cmd),
    .io_uop_mem_size(slots_4_io_uop_mem_size),
    .io_uop_mem_signed(slots_4_io_uop_mem_signed),
    .io_uop_is_fence(slots_4_io_uop_is_fence),
    .io_uop_is_fencei(slots_4_io_uop_is_fencei),
    .io_uop_is_amo(slots_4_io_uop_is_amo),
    .io_uop_uses_ldq(slots_4_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_4_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_4_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_4_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_4_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_4_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_4_io_uop_ldst),
    .io_uop_lrs1(slots_4_io_uop_lrs1),
    .io_uop_lrs2(slots_4_io_uop_lrs2),
    .io_uop_lrs3(slots_4_io_uop_lrs3),
    .io_uop_ldst_val(slots_4_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_4_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_4_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_4_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_4_io_uop_frs3_en),
    .io_uop_fp_val(slots_4_io_uop_fp_val),
    .io_uop_fp_single(slots_4_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_4_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_4_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_4_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_4_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_4_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_4_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_4_io_uop_debug_tsrc),
    .io_debug_p1(slots_4_io_debug_p1),
    .io_debug_p2(slots_4_io_debug_p2),
    .io_debug_p3(slots_4_io_debug_p3),
    .io_debug_ppred(slots_4_io_debug_ppred),
    .io_debug_state(slots_4_io_debug_state)
  );
  IssueSlot slots_5 ( // @[issue-unit.scala 157:73]
    .clock(slots_5_clock),
    .reset(slots_5_reset),
    .io_valid(slots_5_io_valid),
    .io_will_be_valid(slots_5_io_will_be_valid),
    .io_request(slots_5_io_request),
    .io_request_hp(slots_5_io_request_hp),
    .io_grant(slots_5_io_grant),
    .io_brupdate_b1_resolve_mask(slots_5_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_5_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_5_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_5_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_5_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_5_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_5_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_5_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_5_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_5_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_5_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_5_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_5_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_5_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_5_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_5_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_5_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_5_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_5_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_5_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_5_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_5_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_5_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_5_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_5_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_5_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_5_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_5_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_5_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_5_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_5_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_5_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_5_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_5_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_5_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_5_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_5_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_5_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_5_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_5_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_5_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_5_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_5_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_5_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_5_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_5_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_5_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_5_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_5_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_5_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_5_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_5_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_5_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_5_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_5_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_5_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_5_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_5_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_5_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_5_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_5_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_5_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_5_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_5_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_5_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_5_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_5_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_5_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_5_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_5_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_5_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_5_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_5_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_5_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_5_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_5_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_5_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_5_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_5_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_5_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_5_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_5_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_5_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_5_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_5_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_5_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_5_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_5_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_5_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_5_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_5_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_5_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_5_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_5_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_5_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_5_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_5_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_5_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_5_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_5_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_5_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_5_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_5_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_5_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_5_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_5_io_brupdate_b2_target_offset),
    .io_kill(slots_5_io_kill),
    .io_clear(slots_5_io_clear),
    .io_ldspec_miss(slots_5_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_5_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_5_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_5_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_5_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_5_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_5_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_5_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_5_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_5_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_5_io_wakeup_ports_1_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_5_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_5_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_5_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_5_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_5_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_5_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_5_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_5_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_5_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_5_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_5_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_5_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_5_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_5_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_5_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_5_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_5_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_5_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_5_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_5_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_5_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_5_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_5_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_5_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_5_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_5_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_5_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_5_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_5_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_5_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_5_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_5_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_5_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_5_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_5_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_5_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_5_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_5_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_5_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_5_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_5_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_5_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_5_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_5_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_5_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_5_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_5_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_5_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_5_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_5_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_5_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_5_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_5_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_5_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_5_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_5_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_5_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_5_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_5_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_5_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_5_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_5_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_5_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_5_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_5_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_5_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_5_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_5_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_5_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_5_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_5_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_5_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_5_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_5_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_5_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_5_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_5_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_5_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_5_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_5_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_5_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_5_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_5_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_5_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_5_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_5_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_5_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_5_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_5_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_5_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_5_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_5_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_5_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_5_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_5_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_5_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_5_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_5_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_5_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_5_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_5_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_5_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_5_io_out_uop_switch),
    .io_out_uop_switch_off(slots_5_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_5_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_5_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_5_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_5_io_out_uop_rflag),
    .io_out_uop_wflag(slots_5_io_out_uop_wflag),
    .io_out_uop_prflag(slots_5_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_5_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_5_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_5_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_5_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_5_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_5_io_out_uop_split_num),
    .io_out_uop_self_index(slots_5_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_5_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_5_io_out_uop_address_num),
    .io_out_uop_uopc(slots_5_io_out_uop_uopc),
    .io_out_uop_inst(slots_5_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_5_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_5_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_5_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_5_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_5_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_5_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_5_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_5_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_5_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_5_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_5_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_5_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_5_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_5_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_5_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_5_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_5_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_5_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_5_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_5_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_5_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_5_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_5_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_5_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_5_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_5_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_5_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_5_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_5_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_5_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_5_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_5_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_5_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_5_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_5_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_5_io_out_uop_pdst),
    .io_out_uop_prs1(slots_5_io_out_uop_prs1),
    .io_out_uop_prs2(slots_5_io_out_uop_prs2),
    .io_out_uop_prs3(slots_5_io_out_uop_prs3),
    .io_out_uop_ppred(slots_5_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_5_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_5_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_5_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_5_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_5_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_5_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_5_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_5_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_5_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_5_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_5_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_5_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_5_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_5_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_5_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_5_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_5_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_5_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_5_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_5_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_5_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_5_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_5_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_5_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_5_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_5_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_5_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_5_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_5_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_5_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_5_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_5_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_5_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_5_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_5_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_5_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_5_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_5_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_5_io_uop_switch),
    .io_uop_switch_off(slots_5_io_uop_switch_off),
    .io_uop_is_unicore(slots_5_io_uop_is_unicore),
    .io_uop_shift(slots_5_io_uop_shift),
    .io_uop_lrs3_rtype(slots_5_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_5_io_uop_rflag),
    .io_uop_wflag(slots_5_io_uop_wflag),
    .io_uop_prflag(slots_5_io_uop_prflag),
    .io_uop_pwflag(slots_5_io_uop_pwflag),
    .io_uop_pflag_busy(slots_5_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_5_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_5_io_uop_op1_sel),
    .io_uop_op2_sel(slots_5_io_uop_op2_sel),
    .io_uop_split_num(slots_5_io_uop_split_num),
    .io_uop_self_index(slots_5_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_5_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_5_io_uop_address_num),
    .io_uop_uopc(slots_5_io_uop_uopc),
    .io_uop_inst(slots_5_io_uop_inst),
    .io_uop_debug_inst(slots_5_io_uop_debug_inst),
    .io_uop_is_rvc(slots_5_io_uop_is_rvc),
    .io_uop_debug_pc(slots_5_io_uop_debug_pc),
    .io_uop_iq_type(slots_5_io_uop_iq_type),
    .io_uop_fu_code(slots_5_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_5_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_5_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_5_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_5_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_5_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_5_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_5_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_5_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_5_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_5_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_5_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_5_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_5_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_5_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_5_io_uop_is_br),
    .io_uop_is_jalr(slots_5_io_uop_is_jalr),
    .io_uop_is_jal(slots_5_io_uop_is_jal),
    .io_uop_is_sfb(slots_5_io_uop_is_sfb),
    .io_uop_br_mask(slots_5_io_uop_br_mask),
    .io_uop_br_tag(slots_5_io_uop_br_tag),
    .io_uop_ftq_idx(slots_5_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_5_io_uop_edge_inst),
    .io_uop_pc_lob(slots_5_io_uop_pc_lob),
    .io_uop_taken(slots_5_io_uop_taken),
    .io_uop_imm_packed(slots_5_io_uop_imm_packed),
    .io_uop_csr_addr(slots_5_io_uop_csr_addr),
    .io_uop_rob_idx(slots_5_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_5_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_5_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_5_io_uop_rxq_idx),
    .io_uop_pdst(slots_5_io_uop_pdst),
    .io_uop_prs1(slots_5_io_uop_prs1),
    .io_uop_prs2(slots_5_io_uop_prs2),
    .io_uop_prs3(slots_5_io_uop_prs3),
    .io_uop_ppred(slots_5_io_uop_ppred),
    .io_uop_prs1_busy(slots_5_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_5_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_5_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_5_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_5_io_uop_stale_pdst),
    .io_uop_exception(slots_5_io_uop_exception),
    .io_uop_exc_cause(slots_5_io_uop_exc_cause),
    .io_uop_bypassable(slots_5_io_uop_bypassable),
    .io_uop_mem_cmd(slots_5_io_uop_mem_cmd),
    .io_uop_mem_size(slots_5_io_uop_mem_size),
    .io_uop_mem_signed(slots_5_io_uop_mem_signed),
    .io_uop_is_fence(slots_5_io_uop_is_fence),
    .io_uop_is_fencei(slots_5_io_uop_is_fencei),
    .io_uop_is_amo(slots_5_io_uop_is_amo),
    .io_uop_uses_ldq(slots_5_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_5_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_5_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_5_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_5_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_5_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_5_io_uop_ldst),
    .io_uop_lrs1(slots_5_io_uop_lrs1),
    .io_uop_lrs2(slots_5_io_uop_lrs2),
    .io_uop_lrs3(slots_5_io_uop_lrs3),
    .io_uop_ldst_val(slots_5_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_5_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_5_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_5_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_5_io_uop_frs3_en),
    .io_uop_fp_val(slots_5_io_uop_fp_val),
    .io_uop_fp_single(slots_5_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_5_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_5_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_5_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_5_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_5_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_5_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_5_io_uop_debug_tsrc),
    .io_debug_p1(slots_5_io_debug_p1),
    .io_debug_p2(slots_5_io_debug_p2),
    .io_debug_p3(slots_5_io_debug_p3),
    .io_debug_ppred(slots_5_io_debug_ppred),
    .io_debug_state(slots_5_io_debug_state)
  );
  IssueSlot slots_6 ( // @[issue-unit.scala 157:73]
    .clock(slots_6_clock),
    .reset(slots_6_reset),
    .io_valid(slots_6_io_valid),
    .io_will_be_valid(slots_6_io_will_be_valid),
    .io_request(slots_6_io_request),
    .io_request_hp(slots_6_io_request_hp),
    .io_grant(slots_6_io_grant),
    .io_brupdate_b1_resolve_mask(slots_6_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_6_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_6_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_6_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_6_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_6_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_6_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_6_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_6_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_6_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_6_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_6_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_6_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_6_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_6_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_6_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_6_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_6_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_6_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_6_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_6_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_6_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_6_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_6_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_6_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_6_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_6_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_6_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_6_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_6_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_6_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_6_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_6_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_6_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_6_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_6_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_6_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_6_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_6_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_6_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_6_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_6_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_6_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_6_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_6_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_6_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_6_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_6_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_6_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_6_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_6_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_6_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_6_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_6_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_6_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_6_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_6_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_6_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_6_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_6_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_6_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_6_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_6_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_6_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_6_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_6_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_6_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_6_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_6_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_6_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_6_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_6_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_6_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_6_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_6_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_6_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_6_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_6_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_6_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_6_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_6_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_6_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_6_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_6_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_6_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_6_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_6_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_6_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_6_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_6_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_6_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_6_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_6_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_6_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_6_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_6_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_6_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_6_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_6_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_6_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_6_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_6_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_6_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_6_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_6_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_6_io_brupdate_b2_target_offset),
    .io_kill(slots_6_io_kill),
    .io_clear(slots_6_io_clear),
    .io_ldspec_miss(slots_6_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_6_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_6_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_6_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_6_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_6_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_6_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_6_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_6_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_6_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_6_io_wakeup_ports_1_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_6_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_6_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_6_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_6_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_6_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_6_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_6_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_6_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_6_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_6_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_6_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_6_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_6_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_6_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_6_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_6_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_6_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_6_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_6_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_6_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_6_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_6_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_6_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_6_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_6_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_6_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_6_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_6_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_6_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_6_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_6_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_6_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_6_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_6_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_6_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_6_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_6_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_6_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_6_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_6_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_6_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_6_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_6_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_6_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_6_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_6_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_6_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_6_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_6_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_6_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_6_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_6_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_6_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_6_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_6_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_6_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_6_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_6_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_6_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_6_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_6_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_6_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_6_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_6_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_6_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_6_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_6_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_6_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_6_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_6_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_6_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_6_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_6_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_6_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_6_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_6_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_6_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_6_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_6_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_6_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_6_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_6_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_6_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_6_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_6_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_6_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_6_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_6_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_6_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_6_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_6_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_6_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_6_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_6_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_6_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_6_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_6_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_6_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_6_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_6_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_6_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_6_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_6_io_out_uop_switch),
    .io_out_uop_switch_off(slots_6_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_6_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_6_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_6_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_6_io_out_uop_rflag),
    .io_out_uop_wflag(slots_6_io_out_uop_wflag),
    .io_out_uop_prflag(slots_6_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_6_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_6_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_6_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_6_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_6_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_6_io_out_uop_split_num),
    .io_out_uop_self_index(slots_6_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_6_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_6_io_out_uop_address_num),
    .io_out_uop_uopc(slots_6_io_out_uop_uopc),
    .io_out_uop_inst(slots_6_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_6_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_6_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_6_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_6_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_6_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_6_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_6_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_6_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_6_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_6_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_6_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_6_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_6_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_6_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_6_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_6_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_6_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_6_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_6_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_6_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_6_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_6_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_6_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_6_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_6_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_6_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_6_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_6_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_6_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_6_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_6_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_6_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_6_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_6_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_6_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_6_io_out_uop_pdst),
    .io_out_uop_prs1(slots_6_io_out_uop_prs1),
    .io_out_uop_prs2(slots_6_io_out_uop_prs2),
    .io_out_uop_prs3(slots_6_io_out_uop_prs3),
    .io_out_uop_ppred(slots_6_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_6_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_6_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_6_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_6_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_6_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_6_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_6_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_6_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_6_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_6_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_6_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_6_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_6_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_6_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_6_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_6_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_6_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_6_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_6_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_6_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_6_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_6_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_6_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_6_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_6_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_6_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_6_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_6_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_6_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_6_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_6_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_6_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_6_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_6_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_6_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_6_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_6_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_6_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_6_io_uop_switch),
    .io_uop_switch_off(slots_6_io_uop_switch_off),
    .io_uop_is_unicore(slots_6_io_uop_is_unicore),
    .io_uop_shift(slots_6_io_uop_shift),
    .io_uop_lrs3_rtype(slots_6_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_6_io_uop_rflag),
    .io_uop_wflag(slots_6_io_uop_wflag),
    .io_uop_prflag(slots_6_io_uop_prflag),
    .io_uop_pwflag(slots_6_io_uop_pwflag),
    .io_uop_pflag_busy(slots_6_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_6_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_6_io_uop_op1_sel),
    .io_uop_op2_sel(slots_6_io_uop_op2_sel),
    .io_uop_split_num(slots_6_io_uop_split_num),
    .io_uop_self_index(slots_6_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_6_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_6_io_uop_address_num),
    .io_uop_uopc(slots_6_io_uop_uopc),
    .io_uop_inst(slots_6_io_uop_inst),
    .io_uop_debug_inst(slots_6_io_uop_debug_inst),
    .io_uop_is_rvc(slots_6_io_uop_is_rvc),
    .io_uop_debug_pc(slots_6_io_uop_debug_pc),
    .io_uop_iq_type(slots_6_io_uop_iq_type),
    .io_uop_fu_code(slots_6_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_6_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_6_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_6_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_6_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_6_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_6_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_6_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_6_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_6_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_6_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_6_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_6_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_6_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_6_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_6_io_uop_is_br),
    .io_uop_is_jalr(slots_6_io_uop_is_jalr),
    .io_uop_is_jal(slots_6_io_uop_is_jal),
    .io_uop_is_sfb(slots_6_io_uop_is_sfb),
    .io_uop_br_mask(slots_6_io_uop_br_mask),
    .io_uop_br_tag(slots_6_io_uop_br_tag),
    .io_uop_ftq_idx(slots_6_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_6_io_uop_edge_inst),
    .io_uop_pc_lob(slots_6_io_uop_pc_lob),
    .io_uop_taken(slots_6_io_uop_taken),
    .io_uop_imm_packed(slots_6_io_uop_imm_packed),
    .io_uop_csr_addr(slots_6_io_uop_csr_addr),
    .io_uop_rob_idx(slots_6_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_6_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_6_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_6_io_uop_rxq_idx),
    .io_uop_pdst(slots_6_io_uop_pdst),
    .io_uop_prs1(slots_6_io_uop_prs1),
    .io_uop_prs2(slots_6_io_uop_prs2),
    .io_uop_prs3(slots_6_io_uop_prs3),
    .io_uop_ppred(slots_6_io_uop_ppred),
    .io_uop_prs1_busy(slots_6_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_6_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_6_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_6_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_6_io_uop_stale_pdst),
    .io_uop_exception(slots_6_io_uop_exception),
    .io_uop_exc_cause(slots_6_io_uop_exc_cause),
    .io_uop_bypassable(slots_6_io_uop_bypassable),
    .io_uop_mem_cmd(slots_6_io_uop_mem_cmd),
    .io_uop_mem_size(slots_6_io_uop_mem_size),
    .io_uop_mem_signed(slots_6_io_uop_mem_signed),
    .io_uop_is_fence(slots_6_io_uop_is_fence),
    .io_uop_is_fencei(slots_6_io_uop_is_fencei),
    .io_uop_is_amo(slots_6_io_uop_is_amo),
    .io_uop_uses_ldq(slots_6_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_6_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_6_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_6_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_6_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_6_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_6_io_uop_ldst),
    .io_uop_lrs1(slots_6_io_uop_lrs1),
    .io_uop_lrs2(slots_6_io_uop_lrs2),
    .io_uop_lrs3(slots_6_io_uop_lrs3),
    .io_uop_ldst_val(slots_6_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_6_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_6_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_6_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_6_io_uop_frs3_en),
    .io_uop_fp_val(slots_6_io_uop_fp_val),
    .io_uop_fp_single(slots_6_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_6_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_6_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_6_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_6_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_6_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_6_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_6_io_uop_debug_tsrc),
    .io_debug_p1(slots_6_io_debug_p1),
    .io_debug_p2(slots_6_io_debug_p2),
    .io_debug_p3(slots_6_io_debug_p3),
    .io_debug_ppred(slots_6_io_debug_ppred),
    .io_debug_state(slots_6_io_debug_state)
  );
  IssueSlot slots_7 ( // @[issue-unit.scala 157:73]
    .clock(slots_7_clock),
    .reset(slots_7_reset),
    .io_valid(slots_7_io_valid),
    .io_will_be_valid(slots_7_io_will_be_valid),
    .io_request(slots_7_io_request),
    .io_request_hp(slots_7_io_request_hp),
    .io_grant(slots_7_io_grant),
    .io_brupdate_b1_resolve_mask(slots_7_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_7_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_7_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_7_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_7_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_7_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_7_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_7_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_7_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_7_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_7_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_7_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_7_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_7_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_7_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_7_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_7_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_7_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_7_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_7_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_7_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_7_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_7_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_7_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_7_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_7_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_7_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_7_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_7_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_7_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_7_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_7_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_7_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_7_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_7_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_7_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_7_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_7_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_7_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_7_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_7_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_7_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_7_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_7_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_7_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_7_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_7_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_7_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_7_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_7_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_7_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_7_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_7_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_7_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_7_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_7_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_7_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_7_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_7_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_7_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_7_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_7_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_7_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_7_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_7_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_7_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_7_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_7_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_7_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_7_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_7_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_7_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_7_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_7_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_7_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_7_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_7_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_7_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_7_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_7_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_7_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_7_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_7_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_7_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_7_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_7_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_7_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_7_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_7_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_7_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_7_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_7_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_7_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_7_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_7_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_7_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_7_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_7_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_7_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_7_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_7_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_7_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_7_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_7_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_7_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_7_io_brupdate_b2_target_offset),
    .io_kill(slots_7_io_kill),
    .io_clear(slots_7_io_clear),
    .io_ldspec_miss(slots_7_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_7_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_7_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_7_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_7_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_7_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_7_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_7_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_7_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_7_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_7_io_wakeup_ports_1_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_7_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_7_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_7_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_7_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_7_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_7_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_7_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_7_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_7_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_7_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_7_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_7_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_7_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_7_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_7_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_7_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_7_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_7_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_7_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_7_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_7_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_7_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_7_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_7_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_7_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_7_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_7_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_7_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_7_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_7_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_7_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_7_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_7_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_7_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_7_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_7_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_7_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_7_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_7_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_7_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_7_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_7_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_7_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_7_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_7_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_7_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_7_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_7_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_7_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_7_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_7_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_7_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_7_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_7_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_7_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_7_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_7_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_7_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_7_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_7_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_7_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_7_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_7_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_7_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_7_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_7_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_7_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_7_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_7_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_7_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_7_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_7_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_7_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_7_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_7_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_7_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_7_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_7_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_7_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_7_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_7_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_7_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_7_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_7_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_7_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_7_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_7_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_7_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_7_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_7_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_7_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_7_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_7_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_7_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_7_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_7_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_7_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_7_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_7_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_7_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_7_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_7_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_7_io_out_uop_switch),
    .io_out_uop_switch_off(slots_7_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_7_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_7_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_7_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_7_io_out_uop_rflag),
    .io_out_uop_wflag(slots_7_io_out_uop_wflag),
    .io_out_uop_prflag(slots_7_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_7_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_7_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_7_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_7_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_7_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_7_io_out_uop_split_num),
    .io_out_uop_self_index(slots_7_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_7_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_7_io_out_uop_address_num),
    .io_out_uop_uopc(slots_7_io_out_uop_uopc),
    .io_out_uop_inst(slots_7_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_7_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_7_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_7_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_7_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_7_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_7_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_7_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_7_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_7_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_7_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_7_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_7_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_7_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_7_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_7_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_7_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_7_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_7_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_7_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_7_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_7_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_7_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_7_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_7_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_7_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_7_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_7_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_7_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_7_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_7_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_7_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_7_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_7_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_7_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_7_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_7_io_out_uop_pdst),
    .io_out_uop_prs1(slots_7_io_out_uop_prs1),
    .io_out_uop_prs2(slots_7_io_out_uop_prs2),
    .io_out_uop_prs3(slots_7_io_out_uop_prs3),
    .io_out_uop_ppred(slots_7_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_7_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_7_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_7_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_7_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_7_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_7_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_7_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_7_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_7_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_7_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_7_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_7_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_7_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_7_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_7_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_7_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_7_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_7_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_7_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_7_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_7_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_7_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_7_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_7_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_7_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_7_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_7_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_7_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_7_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_7_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_7_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_7_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_7_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_7_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_7_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_7_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_7_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_7_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_7_io_uop_switch),
    .io_uop_switch_off(slots_7_io_uop_switch_off),
    .io_uop_is_unicore(slots_7_io_uop_is_unicore),
    .io_uop_shift(slots_7_io_uop_shift),
    .io_uop_lrs3_rtype(slots_7_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_7_io_uop_rflag),
    .io_uop_wflag(slots_7_io_uop_wflag),
    .io_uop_prflag(slots_7_io_uop_prflag),
    .io_uop_pwflag(slots_7_io_uop_pwflag),
    .io_uop_pflag_busy(slots_7_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_7_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_7_io_uop_op1_sel),
    .io_uop_op2_sel(slots_7_io_uop_op2_sel),
    .io_uop_split_num(slots_7_io_uop_split_num),
    .io_uop_self_index(slots_7_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_7_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_7_io_uop_address_num),
    .io_uop_uopc(slots_7_io_uop_uopc),
    .io_uop_inst(slots_7_io_uop_inst),
    .io_uop_debug_inst(slots_7_io_uop_debug_inst),
    .io_uop_is_rvc(slots_7_io_uop_is_rvc),
    .io_uop_debug_pc(slots_7_io_uop_debug_pc),
    .io_uop_iq_type(slots_7_io_uop_iq_type),
    .io_uop_fu_code(slots_7_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_7_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_7_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_7_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_7_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_7_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_7_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_7_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_7_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_7_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_7_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_7_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_7_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_7_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_7_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_7_io_uop_is_br),
    .io_uop_is_jalr(slots_7_io_uop_is_jalr),
    .io_uop_is_jal(slots_7_io_uop_is_jal),
    .io_uop_is_sfb(slots_7_io_uop_is_sfb),
    .io_uop_br_mask(slots_7_io_uop_br_mask),
    .io_uop_br_tag(slots_7_io_uop_br_tag),
    .io_uop_ftq_idx(slots_7_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_7_io_uop_edge_inst),
    .io_uop_pc_lob(slots_7_io_uop_pc_lob),
    .io_uop_taken(slots_7_io_uop_taken),
    .io_uop_imm_packed(slots_7_io_uop_imm_packed),
    .io_uop_csr_addr(slots_7_io_uop_csr_addr),
    .io_uop_rob_idx(slots_7_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_7_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_7_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_7_io_uop_rxq_idx),
    .io_uop_pdst(slots_7_io_uop_pdst),
    .io_uop_prs1(slots_7_io_uop_prs1),
    .io_uop_prs2(slots_7_io_uop_prs2),
    .io_uop_prs3(slots_7_io_uop_prs3),
    .io_uop_ppred(slots_7_io_uop_ppred),
    .io_uop_prs1_busy(slots_7_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_7_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_7_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_7_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_7_io_uop_stale_pdst),
    .io_uop_exception(slots_7_io_uop_exception),
    .io_uop_exc_cause(slots_7_io_uop_exc_cause),
    .io_uop_bypassable(slots_7_io_uop_bypassable),
    .io_uop_mem_cmd(slots_7_io_uop_mem_cmd),
    .io_uop_mem_size(slots_7_io_uop_mem_size),
    .io_uop_mem_signed(slots_7_io_uop_mem_signed),
    .io_uop_is_fence(slots_7_io_uop_is_fence),
    .io_uop_is_fencei(slots_7_io_uop_is_fencei),
    .io_uop_is_amo(slots_7_io_uop_is_amo),
    .io_uop_uses_ldq(slots_7_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_7_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_7_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_7_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_7_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_7_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_7_io_uop_ldst),
    .io_uop_lrs1(slots_7_io_uop_lrs1),
    .io_uop_lrs2(slots_7_io_uop_lrs2),
    .io_uop_lrs3(slots_7_io_uop_lrs3),
    .io_uop_ldst_val(slots_7_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_7_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_7_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_7_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_7_io_uop_frs3_en),
    .io_uop_fp_val(slots_7_io_uop_fp_val),
    .io_uop_fp_single(slots_7_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_7_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_7_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_7_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_7_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_7_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_7_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_7_io_uop_debug_tsrc),
    .io_debug_p1(slots_7_io_debug_p1),
    .io_debug_p2(slots_7_io_debug_p2),
    .io_debug_p3(slots_7_io_debug_p3),
    .io_debug_ppred(slots_7_io_debug_ppred),
    .io_debug_state(slots_7_io_debug_state)
  );
  IssueSlot slots_8 ( // @[issue-unit.scala 157:73]
    .clock(slots_8_clock),
    .reset(slots_8_reset),
    .io_valid(slots_8_io_valid),
    .io_will_be_valid(slots_8_io_will_be_valid),
    .io_request(slots_8_io_request),
    .io_request_hp(slots_8_io_request_hp),
    .io_grant(slots_8_io_grant),
    .io_brupdate_b1_resolve_mask(slots_8_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_8_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_8_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_8_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_8_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_8_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_8_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_8_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_8_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_8_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_8_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_8_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_8_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_8_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_8_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_8_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_8_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_8_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_8_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_8_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_8_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_8_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_8_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_8_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_8_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_8_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_8_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_8_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_8_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_8_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_8_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_8_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_8_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_8_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_8_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_8_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_8_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_8_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_8_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_8_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_8_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_8_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_8_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_8_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_8_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_8_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_8_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_8_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_8_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_8_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_8_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_8_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_8_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_8_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_8_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_8_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_8_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_8_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_8_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_8_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_8_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_8_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_8_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_8_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_8_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_8_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_8_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_8_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_8_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_8_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_8_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_8_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_8_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_8_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_8_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_8_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_8_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_8_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_8_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_8_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_8_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_8_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_8_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_8_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_8_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_8_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_8_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_8_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_8_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_8_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_8_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_8_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_8_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_8_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_8_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_8_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_8_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_8_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_8_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_8_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_8_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_8_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_8_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_8_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_8_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_8_io_brupdate_b2_target_offset),
    .io_kill(slots_8_io_kill),
    .io_clear(slots_8_io_clear),
    .io_ldspec_miss(slots_8_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_8_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_8_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_8_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_8_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_8_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_8_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_8_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_8_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_8_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_8_io_wakeup_ports_1_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_8_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_8_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_8_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_8_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_8_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_8_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_8_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_8_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_8_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_8_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_8_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_8_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_8_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_8_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_8_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_8_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_8_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_8_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_8_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_8_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_8_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_8_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_8_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_8_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_8_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_8_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_8_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_8_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_8_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_8_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_8_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_8_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_8_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_8_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_8_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_8_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_8_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_8_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_8_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_8_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_8_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_8_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_8_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_8_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_8_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_8_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_8_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_8_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_8_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_8_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_8_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_8_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_8_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_8_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_8_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_8_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_8_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_8_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_8_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_8_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_8_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_8_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_8_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_8_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_8_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_8_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_8_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_8_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_8_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_8_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_8_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_8_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_8_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_8_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_8_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_8_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_8_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_8_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_8_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_8_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_8_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_8_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_8_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_8_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_8_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_8_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_8_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_8_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_8_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_8_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_8_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_8_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_8_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_8_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_8_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_8_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_8_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_8_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_8_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_8_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_8_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_8_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_8_io_out_uop_switch),
    .io_out_uop_switch_off(slots_8_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_8_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_8_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_8_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_8_io_out_uop_rflag),
    .io_out_uop_wflag(slots_8_io_out_uop_wflag),
    .io_out_uop_prflag(slots_8_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_8_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_8_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_8_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_8_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_8_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_8_io_out_uop_split_num),
    .io_out_uop_self_index(slots_8_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_8_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_8_io_out_uop_address_num),
    .io_out_uop_uopc(slots_8_io_out_uop_uopc),
    .io_out_uop_inst(slots_8_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_8_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_8_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_8_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_8_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_8_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_8_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_8_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_8_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_8_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_8_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_8_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_8_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_8_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_8_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_8_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_8_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_8_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_8_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_8_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_8_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_8_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_8_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_8_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_8_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_8_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_8_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_8_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_8_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_8_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_8_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_8_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_8_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_8_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_8_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_8_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_8_io_out_uop_pdst),
    .io_out_uop_prs1(slots_8_io_out_uop_prs1),
    .io_out_uop_prs2(slots_8_io_out_uop_prs2),
    .io_out_uop_prs3(slots_8_io_out_uop_prs3),
    .io_out_uop_ppred(slots_8_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_8_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_8_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_8_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_8_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_8_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_8_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_8_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_8_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_8_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_8_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_8_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_8_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_8_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_8_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_8_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_8_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_8_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_8_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_8_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_8_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_8_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_8_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_8_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_8_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_8_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_8_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_8_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_8_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_8_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_8_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_8_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_8_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_8_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_8_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_8_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_8_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_8_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_8_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_8_io_uop_switch),
    .io_uop_switch_off(slots_8_io_uop_switch_off),
    .io_uop_is_unicore(slots_8_io_uop_is_unicore),
    .io_uop_shift(slots_8_io_uop_shift),
    .io_uop_lrs3_rtype(slots_8_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_8_io_uop_rflag),
    .io_uop_wflag(slots_8_io_uop_wflag),
    .io_uop_prflag(slots_8_io_uop_prflag),
    .io_uop_pwflag(slots_8_io_uop_pwflag),
    .io_uop_pflag_busy(slots_8_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_8_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_8_io_uop_op1_sel),
    .io_uop_op2_sel(slots_8_io_uop_op2_sel),
    .io_uop_split_num(slots_8_io_uop_split_num),
    .io_uop_self_index(slots_8_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_8_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_8_io_uop_address_num),
    .io_uop_uopc(slots_8_io_uop_uopc),
    .io_uop_inst(slots_8_io_uop_inst),
    .io_uop_debug_inst(slots_8_io_uop_debug_inst),
    .io_uop_is_rvc(slots_8_io_uop_is_rvc),
    .io_uop_debug_pc(slots_8_io_uop_debug_pc),
    .io_uop_iq_type(slots_8_io_uop_iq_type),
    .io_uop_fu_code(slots_8_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_8_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_8_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_8_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_8_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_8_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_8_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_8_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_8_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_8_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_8_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_8_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_8_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_8_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_8_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_8_io_uop_is_br),
    .io_uop_is_jalr(slots_8_io_uop_is_jalr),
    .io_uop_is_jal(slots_8_io_uop_is_jal),
    .io_uop_is_sfb(slots_8_io_uop_is_sfb),
    .io_uop_br_mask(slots_8_io_uop_br_mask),
    .io_uop_br_tag(slots_8_io_uop_br_tag),
    .io_uop_ftq_idx(slots_8_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_8_io_uop_edge_inst),
    .io_uop_pc_lob(slots_8_io_uop_pc_lob),
    .io_uop_taken(slots_8_io_uop_taken),
    .io_uop_imm_packed(slots_8_io_uop_imm_packed),
    .io_uop_csr_addr(slots_8_io_uop_csr_addr),
    .io_uop_rob_idx(slots_8_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_8_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_8_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_8_io_uop_rxq_idx),
    .io_uop_pdst(slots_8_io_uop_pdst),
    .io_uop_prs1(slots_8_io_uop_prs1),
    .io_uop_prs2(slots_8_io_uop_prs2),
    .io_uop_prs3(slots_8_io_uop_prs3),
    .io_uop_ppred(slots_8_io_uop_ppred),
    .io_uop_prs1_busy(slots_8_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_8_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_8_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_8_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_8_io_uop_stale_pdst),
    .io_uop_exception(slots_8_io_uop_exception),
    .io_uop_exc_cause(slots_8_io_uop_exc_cause),
    .io_uop_bypassable(slots_8_io_uop_bypassable),
    .io_uop_mem_cmd(slots_8_io_uop_mem_cmd),
    .io_uop_mem_size(slots_8_io_uop_mem_size),
    .io_uop_mem_signed(slots_8_io_uop_mem_signed),
    .io_uop_is_fence(slots_8_io_uop_is_fence),
    .io_uop_is_fencei(slots_8_io_uop_is_fencei),
    .io_uop_is_amo(slots_8_io_uop_is_amo),
    .io_uop_uses_ldq(slots_8_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_8_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_8_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_8_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_8_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_8_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_8_io_uop_ldst),
    .io_uop_lrs1(slots_8_io_uop_lrs1),
    .io_uop_lrs2(slots_8_io_uop_lrs2),
    .io_uop_lrs3(slots_8_io_uop_lrs3),
    .io_uop_ldst_val(slots_8_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_8_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_8_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_8_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_8_io_uop_frs3_en),
    .io_uop_fp_val(slots_8_io_uop_fp_val),
    .io_uop_fp_single(slots_8_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_8_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_8_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_8_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_8_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_8_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_8_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_8_io_uop_debug_tsrc),
    .io_debug_p1(slots_8_io_debug_p1),
    .io_debug_p2(slots_8_io_debug_p2),
    .io_debug_p3(slots_8_io_debug_p3),
    .io_debug_ppred(slots_8_io_debug_ppred),
    .io_debug_state(slots_8_io_debug_state)
  );
  IssueSlot slots_9 ( // @[issue-unit.scala 157:73]
    .clock(slots_9_clock),
    .reset(slots_9_reset),
    .io_valid(slots_9_io_valid),
    .io_will_be_valid(slots_9_io_will_be_valid),
    .io_request(slots_9_io_request),
    .io_request_hp(slots_9_io_request_hp),
    .io_grant(slots_9_io_grant),
    .io_brupdate_b1_resolve_mask(slots_9_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_9_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_9_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_9_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_9_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_9_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_9_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_9_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_9_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_9_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_9_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_9_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_9_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_9_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_9_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_9_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_9_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_9_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_9_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_9_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_9_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_9_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_9_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_9_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_9_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_9_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_9_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_9_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_9_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_9_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_9_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_9_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_9_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_9_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_9_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_9_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_9_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_9_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_9_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_9_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_9_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_9_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_9_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_9_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_9_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_9_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_9_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_9_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_9_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_9_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_9_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_9_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_9_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_9_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_9_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_9_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_9_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_9_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_9_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_9_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_9_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_9_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_9_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_9_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_9_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_9_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_9_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_9_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_9_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_9_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_9_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_9_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_9_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_9_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_9_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_9_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_9_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_9_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_9_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_9_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_9_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_9_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_9_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_9_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_9_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_9_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_9_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_9_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_9_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_9_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_9_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_9_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_9_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_9_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_9_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_9_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_9_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_9_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_9_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_9_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_9_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_9_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_9_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_9_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_9_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_9_io_brupdate_b2_target_offset),
    .io_kill(slots_9_io_kill),
    .io_clear(slots_9_io_clear),
    .io_ldspec_miss(slots_9_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_9_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_9_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_9_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_9_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_9_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_9_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_9_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_9_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_9_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_9_io_wakeup_ports_1_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_9_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_9_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_9_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_9_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_9_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_9_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_9_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_9_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_9_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_9_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_9_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_9_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_9_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_9_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_9_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_9_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_9_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_9_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_9_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_9_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_9_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_9_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_9_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_9_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_9_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_9_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_9_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_9_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_9_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_9_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_9_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_9_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_9_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_9_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_9_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_9_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_9_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_9_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_9_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_9_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_9_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_9_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_9_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_9_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_9_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_9_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_9_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_9_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_9_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_9_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_9_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_9_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_9_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_9_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_9_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_9_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_9_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_9_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_9_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_9_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_9_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_9_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_9_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_9_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_9_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_9_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_9_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_9_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_9_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_9_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_9_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_9_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_9_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_9_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_9_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_9_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_9_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_9_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_9_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_9_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_9_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_9_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_9_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_9_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_9_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_9_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_9_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_9_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_9_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_9_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_9_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_9_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_9_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_9_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_9_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_9_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_9_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_9_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_9_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_9_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_9_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_9_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_9_io_out_uop_switch),
    .io_out_uop_switch_off(slots_9_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_9_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_9_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_9_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_9_io_out_uop_rflag),
    .io_out_uop_wflag(slots_9_io_out_uop_wflag),
    .io_out_uop_prflag(slots_9_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_9_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_9_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_9_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_9_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_9_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_9_io_out_uop_split_num),
    .io_out_uop_self_index(slots_9_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_9_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_9_io_out_uop_address_num),
    .io_out_uop_uopc(slots_9_io_out_uop_uopc),
    .io_out_uop_inst(slots_9_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_9_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_9_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_9_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_9_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_9_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_9_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_9_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_9_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_9_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_9_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_9_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_9_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_9_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_9_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_9_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_9_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_9_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_9_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_9_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_9_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_9_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_9_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_9_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_9_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_9_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_9_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_9_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_9_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_9_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_9_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_9_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_9_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_9_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_9_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_9_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_9_io_out_uop_pdst),
    .io_out_uop_prs1(slots_9_io_out_uop_prs1),
    .io_out_uop_prs2(slots_9_io_out_uop_prs2),
    .io_out_uop_prs3(slots_9_io_out_uop_prs3),
    .io_out_uop_ppred(slots_9_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_9_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_9_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_9_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_9_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_9_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_9_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_9_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_9_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_9_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_9_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_9_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_9_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_9_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_9_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_9_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_9_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_9_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_9_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_9_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_9_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_9_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_9_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_9_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_9_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_9_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_9_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_9_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_9_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_9_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_9_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_9_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_9_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_9_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_9_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_9_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_9_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_9_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_9_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_9_io_uop_switch),
    .io_uop_switch_off(slots_9_io_uop_switch_off),
    .io_uop_is_unicore(slots_9_io_uop_is_unicore),
    .io_uop_shift(slots_9_io_uop_shift),
    .io_uop_lrs3_rtype(slots_9_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_9_io_uop_rflag),
    .io_uop_wflag(slots_9_io_uop_wflag),
    .io_uop_prflag(slots_9_io_uop_prflag),
    .io_uop_pwflag(slots_9_io_uop_pwflag),
    .io_uop_pflag_busy(slots_9_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_9_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_9_io_uop_op1_sel),
    .io_uop_op2_sel(slots_9_io_uop_op2_sel),
    .io_uop_split_num(slots_9_io_uop_split_num),
    .io_uop_self_index(slots_9_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_9_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_9_io_uop_address_num),
    .io_uop_uopc(slots_9_io_uop_uopc),
    .io_uop_inst(slots_9_io_uop_inst),
    .io_uop_debug_inst(slots_9_io_uop_debug_inst),
    .io_uop_is_rvc(slots_9_io_uop_is_rvc),
    .io_uop_debug_pc(slots_9_io_uop_debug_pc),
    .io_uop_iq_type(slots_9_io_uop_iq_type),
    .io_uop_fu_code(slots_9_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_9_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_9_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_9_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_9_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_9_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_9_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_9_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_9_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_9_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_9_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_9_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_9_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_9_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_9_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_9_io_uop_is_br),
    .io_uop_is_jalr(slots_9_io_uop_is_jalr),
    .io_uop_is_jal(slots_9_io_uop_is_jal),
    .io_uop_is_sfb(slots_9_io_uop_is_sfb),
    .io_uop_br_mask(slots_9_io_uop_br_mask),
    .io_uop_br_tag(slots_9_io_uop_br_tag),
    .io_uop_ftq_idx(slots_9_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_9_io_uop_edge_inst),
    .io_uop_pc_lob(slots_9_io_uop_pc_lob),
    .io_uop_taken(slots_9_io_uop_taken),
    .io_uop_imm_packed(slots_9_io_uop_imm_packed),
    .io_uop_csr_addr(slots_9_io_uop_csr_addr),
    .io_uop_rob_idx(slots_9_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_9_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_9_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_9_io_uop_rxq_idx),
    .io_uop_pdst(slots_9_io_uop_pdst),
    .io_uop_prs1(slots_9_io_uop_prs1),
    .io_uop_prs2(slots_9_io_uop_prs2),
    .io_uop_prs3(slots_9_io_uop_prs3),
    .io_uop_ppred(slots_9_io_uop_ppred),
    .io_uop_prs1_busy(slots_9_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_9_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_9_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_9_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_9_io_uop_stale_pdst),
    .io_uop_exception(slots_9_io_uop_exception),
    .io_uop_exc_cause(slots_9_io_uop_exc_cause),
    .io_uop_bypassable(slots_9_io_uop_bypassable),
    .io_uop_mem_cmd(slots_9_io_uop_mem_cmd),
    .io_uop_mem_size(slots_9_io_uop_mem_size),
    .io_uop_mem_signed(slots_9_io_uop_mem_signed),
    .io_uop_is_fence(slots_9_io_uop_is_fence),
    .io_uop_is_fencei(slots_9_io_uop_is_fencei),
    .io_uop_is_amo(slots_9_io_uop_is_amo),
    .io_uop_uses_ldq(slots_9_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_9_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_9_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_9_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_9_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_9_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_9_io_uop_ldst),
    .io_uop_lrs1(slots_9_io_uop_lrs1),
    .io_uop_lrs2(slots_9_io_uop_lrs2),
    .io_uop_lrs3(slots_9_io_uop_lrs3),
    .io_uop_ldst_val(slots_9_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_9_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_9_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_9_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_9_io_uop_frs3_en),
    .io_uop_fp_val(slots_9_io_uop_fp_val),
    .io_uop_fp_single(slots_9_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_9_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_9_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_9_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_9_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_9_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_9_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_9_io_uop_debug_tsrc),
    .io_debug_p1(slots_9_io_debug_p1),
    .io_debug_p2(slots_9_io_debug_p2),
    .io_debug_p3(slots_9_io_debug_p3),
    .io_debug_ppred(slots_9_io_debug_ppred),
    .io_debug_state(slots_9_io_debug_state)
  );
  IssueSlot slots_10 ( // @[issue-unit.scala 157:73]
    .clock(slots_10_clock),
    .reset(slots_10_reset),
    .io_valid(slots_10_io_valid),
    .io_will_be_valid(slots_10_io_will_be_valid),
    .io_request(slots_10_io_request),
    .io_request_hp(slots_10_io_request_hp),
    .io_grant(slots_10_io_grant),
    .io_brupdate_b1_resolve_mask(slots_10_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_10_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_10_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_10_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_10_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_10_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_10_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_10_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_10_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_10_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_10_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_10_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_10_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_10_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_10_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_10_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_10_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_10_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_10_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_10_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_10_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_10_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_10_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_10_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_10_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_10_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_10_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_10_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_10_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_10_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_10_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_10_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_10_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_10_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_10_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_10_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_10_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_10_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_10_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_10_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_10_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_10_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_10_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_10_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_10_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_10_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_10_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_10_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_10_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_10_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_10_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_10_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_10_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_10_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_10_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_10_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_10_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_10_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_10_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_10_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_10_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_10_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_10_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_10_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_10_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_10_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_10_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_10_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_10_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_10_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_10_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_10_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_10_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_10_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_10_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_10_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_10_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_10_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_10_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_10_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_10_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_10_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_10_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_10_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_10_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_10_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_10_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_10_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_10_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_10_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_10_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_10_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_10_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_10_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_10_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_10_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_10_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_10_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_10_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_10_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_10_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_10_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_10_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_10_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_10_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_10_io_brupdate_b2_target_offset),
    .io_kill(slots_10_io_kill),
    .io_clear(slots_10_io_clear),
    .io_ldspec_miss(slots_10_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_10_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_10_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_10_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_10_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_10_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_10_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_10_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_10_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_10_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_10_io_wakeup_ports_1_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_10_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_10_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_10_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_10_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_10_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_10_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_10_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_10_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_10_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_10_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_10_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_10_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_10_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_10_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_10_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_10_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_10_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_10_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_10_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_10_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_10_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_10_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_10_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_10_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_10_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_10_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_10_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_10_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_10_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_10_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_10_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_10_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_10_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_10_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_10_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_10_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_10_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_10_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_10_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_10_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_10_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_10_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_10_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_10_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_10_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_10_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_10_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_10_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_10_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_10_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_10_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_10_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_10_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_10_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_10_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_10_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_10_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_10_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_10_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_10_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_10_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_10_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_10_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_10_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_10_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_10_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_10_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_10_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_10_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_10_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_10_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_10_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_10_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_10_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_10_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_10_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_10_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_10_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_10_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_10_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_10_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_10_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_10_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_10_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_10_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_10_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_10_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_10_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_10_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_10_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_10_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_10_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_10_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_10_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_10_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_10_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_10_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_10_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_10_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_10_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_10_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_10_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_10_io_out_uop_switch),
    .io_out_uop_switch_off(slots_10_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_10_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_10_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_10_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_10_io_out_uop_rflag),
    .io_out_uop_wflag(slots_10_io_out_uop_wflag),
    .io_out_uop_prflag(slots_10_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_10_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_10_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_10_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_10_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_10_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_10_io_out_uop_split_num),
    .io_out_uop_self_index(slots_10_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_10_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_10_io_out_uop_address_num),
    .io_out_uop_uopc(slots_10_io_out_uop_uopc),
    .io_out_uop_inst(slots_10_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_10_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_10_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_10_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_10_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_10_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_10_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_10_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_10_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_10_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_10_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_10_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_10_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_10_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_10_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_10_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_10_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_10_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_10_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_10_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_10_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_10_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_10_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_10_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_10_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_10_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_10_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_10_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_10_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_10_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_10_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_10_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_10_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_10_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_10_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_10_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_10_io_out_uop_pdst),
    .io_out_uop_prs1(slots_10_io_out_uop_prs1),
    .io_out_uop_prs2(slots_10_io_out_uop_prs2),
    .io_out_uop_prs3(slots_10_io_out_uop_prs3),
    .io_out_uop_ppred(slots_10_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_10_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_10_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_10_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_10_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_10_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_10_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_10_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_10_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_10_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_10_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_10_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_10_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_10_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_10_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_10_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_10_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_10_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_10_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_10_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_10_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_10_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_10_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_10_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_10_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_10_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_10_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_10_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_10_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_10_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_10_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_10_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_10_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_10_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_10_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_10_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_10_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_10_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_10_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_10_io_uop_switch),
    .io_uop_switch_off(slots_10_io_uop_switch_off),
    .io_uop_is_unicore(slots_10_io_uop_is_unicore),
    .io_uop_shift(slots_10_io_uop_shift),
    .io_uop_lrs3_rtype(slots_10_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_10_io_uop_rflag),
    .io_uop_wflag(slots_10_io_uop_wflag),
    .io_uop_prflag(slots_10_io_uop_prflag),
    .io_uop_pwflag(slots_10_io_uop_pwflag),
    .io_uop_pflag_busy(slots_10_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_10_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_10_io_uop_op1_sel),
    .io_uop_op2_sel(slots_10_io_uop_op2_sel),
    .io_uop_split_num(slots_10_io_uop_split_num),
    .io_uop_self_index(slots_10_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_10_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_10_io_uop_address_num),
    .io_uop_uopc(slots_10_io_uop_uopc),
    .io_uop_inst(slots_10_io_uop_inst),
    .io_uop_debug_inst(slots_10_io_uop_debug_inst),
    .io_uop_is_rvc(slots_10_io_uop_is_rvc),
    .io_uop_debug_pc(slots_10_io_uop_debug_pc),
    .io_uop_iq_type(slots_10_io_uop_iq_type),
    .io_uop_fu_code(slots_10_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_10_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_10_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_10_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_10_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_10_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_10_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_10_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_10_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_10_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_10_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_10_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_10_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_10_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_10_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_10_io_uop_is_br),
    .io_uop_is_jalr(slots_10_io_uop_is_jalr),
    .io_uop_is_jal(slots_10_io_uop_is_jal),
    .io_uop_is_sfb(slots_10_io_uop_is_sfb),
    .io_uop_br_mask(slots_10_io_uop_br_mask),
    .io_uop_br_tag(slots_10_io_uop_br_tag),
    .io_uop_ftq_idx(slots_10_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_10_io_uop_edge_inst),
    .io_uop_pc_lob(slots_10_io_uop_pc_lob),
    .io_uop_taken(slots_10_io_uop_taken),
    .io_uop_imm_packed(slots_10_io_uop_imm_packed),
    .io_uop_csr_addr(slots_10_io_uop_csr_addr),
    .io_uop_rob_idx(slots_10_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_10_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_10_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_10_io_uop_rxq_idx),
    .io_uop_pdst(slots_10_io_uop_pdst),
    .io_uop_prs1(slots_10_io_uop_prs1),
    .io_uop_prs2(slots_10_io_uop_prs2),
    .io_uop_prs3(slots_10_io_uop_prs3),
    .io_uop_ppred(slots_10_io_uop_ppred),
    .io_uop_prs1_busy(slots_10_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_10_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_10_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_10_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_10_io_uop_stale_pdst),
    .io_uop_exception(slots_10_io_uop_exception),
    .io_uop_exc_cause(slots_10_io_uop_exc_cause),
    .io_uop_bypassable(slots_10_io_uop_bypassable),
    .io_uop_mem_cmd(slots_10_io_uop_mem_cmd),
    .io_uop_mem_size(slots_10_io_uop_mem_size),
    .io_uop_mem_signed(slots_10_io_uop_mem_signed),
    .io_uop_is_fence(slots_10_io_uop_is_fence),
    .io_uop_is_fencei(slots_10_io_uop_is_fencei),
    .io_uop_is_amo(slots_10_io_uop_is_amo),
    .io_uop_uses_ldq(slots_10_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_10_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_10_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_10_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_10_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_10_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_10_io_uop_ldst),
    .io_uop_lrs1(slots_10_io_uop_lrs1),
    .io_uop_lrs2(slots_10_io_uop_lrs2),
    .io_uop_lrs3(slots_10_io_uop_lrs3),
    .io_uop_ldst_val(slots_10_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_10_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_10_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_10_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_10_io_uop_frs3_en),
    .io_uop_fp_val(slots_10_io_uop_fp_val),
    .io_uop_fp_single(slots_10_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_10_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_10_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_10_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_10_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_10_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_10_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_10_io_uop_debug_tsrc),
    .io_debug_p1(slots_10_io_debug_p1),
    .io_debug_p2(slots_10_io_debug_p2),
    .io_debug_p3(slots_10_io_debug_p3),
    .io_debug_ppred(slots_10_io_debug_ppred),
    .io_debug_state(slots_10_io_debug_state)
  );
  IssueSlot slots_11 ( // @[issue-unit.scala 157:73]
    .clock(slots_11_clock),
    .reset(slots_11_reset),
    .io_valid(slots_11_io_valid),
    .io_will_be_valid(slots_11_io_will_be_valid),
    .io_request(slots_11_io_request),
    .io_request_hp(slots_11_io_request_hp),
    .io_grant(slots_11_io_grant),
    .io_brupdate_b1_resolve_mask(slots_11_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_11_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_11_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_11_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_11_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_11_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_11_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_11_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_11_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_11_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_11_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_11_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_11_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_11_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_11_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_11_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_11_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_11_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_11_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_11_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_11_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_11_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_11_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_11_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_11_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_11_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_11_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_11_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_11_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_11_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_11_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_11_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_11_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_11_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_11_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_11_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_11_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_11_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_11_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_11_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_11_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_11_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_11_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_11_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_11_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_11_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_11_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_11_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_11_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_11_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_11_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_11_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_11_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_11_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_11_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_11_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_11_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_11_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_11_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_11_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_11_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_11_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_11_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_11_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_11_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_11_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_11_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_11_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_11_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_11_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_11_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_11_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_11_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_11_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_11_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_11_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_11_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_11_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_11_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_11_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_11_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_11_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_11_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_11_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_11_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_11_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_11_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_11_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_11_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_11_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_11_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_11_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_11_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_11_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_11_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_11_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_11_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_11_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_11_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_11_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_11_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_11_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_11_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_11_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_11_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_11_io_brupdate_b2_target_offset),
    .io_kill(slots_11_io_kill),
    .io_clear(slots_11_io_clear),
    .io_ldspec_miss(slots_11_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_11_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_11_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_11_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_11_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_11_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_11_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_11_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_11_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_11_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_11_io_wakeup_ports_1_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_11_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_11_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_11_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_11_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_11_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_11_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_11_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_11_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_11_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_11_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_11_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_11_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_11_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_11_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_11_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_11_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_11_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_11_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_11_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_11_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_11_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_11_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_11_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_11_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_11_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_11_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_11_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_11_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_11_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_11_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_11_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_11_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_11_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_11_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_11_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_11_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_11_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_11_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_11_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_11_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_11_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_11_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_11_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_11_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_11_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_11_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_11_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_11_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_11_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_11_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_11_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_11_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_11_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_11_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_11_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_11_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_11_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_11_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_11_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_11_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_11_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_11_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_11_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_11_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_11_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_11_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_11_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_11_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_11_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_11_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_11_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_11_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_11_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_11_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_11_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_11_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_11_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_11_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_11_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_11_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_11_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_11_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_11_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_11_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_11_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_11_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_11_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_11_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_11_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_11_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_11_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_11_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_11_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_11_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_11_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_11_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_11_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_11_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_11_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_11_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_11_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_11_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_11_io_out_uop_switch),
    .io_out_uop_switch_off(slots_11_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_11_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_11_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_11_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_11_io_out_uop_rflag),
    .io_out_uop_wflag(slots_11_io_out_uop_wflag),
    .io_out_uop_prflag(slots_11_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_11_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_11_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_11_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_11_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_11_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_11_io_out_uop_split_num),
    .io_out_uop_self_index(slots_11_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_11_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_11_io_out_uop_address_num),
    .io_out_uop_uopc(slots_11_io_out_uop_uopc),
    .io_out_uop_inst(slots_11_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_11_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_11_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_11_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_11_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_11_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_11_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_11_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_11_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_11_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_11_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_11_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_11_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_11_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_11_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_11_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_11_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_11_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_11_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_11_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_11_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_11_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_11_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_11_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_11_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_11_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_11_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_11_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_11_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_11_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_11_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_11_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_11_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_11_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_11_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_11_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_11_io_out_uop_pdst),
    .io_out_uop_prs1(slots_11_io_out_uop_prs1),
    .io_out_uop_prs2(slots_11_io_out_uop_prs2),
    .io_out_uop_prs3(slots_11_io_out_uop_prs3),
    .io_out_uop_ppred(slots_11_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_11_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_11_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_11_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_11_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_11_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_11_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_11_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_11_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_11_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_11_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_11_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_11_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_11_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_11_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_11_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_11_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_11_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_11_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_11_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_11_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_11_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_11_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_11_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_11_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_11_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_11_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_11_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_11_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_11_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_11_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_11_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_11_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_11_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_11_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_11_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_11_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_11_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_11_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_11_io_uop_switch),
    .io_uop_switch_off(slots_11_io_uop_switch_off),
    .io_uop_is_unicore(slots_11_io_uop_is_unicore),
    .io_uop_shift(slots_11_io_uop_shift),
    .io_uop_lrs3_rtype(slots_11_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_11_io_uop_rflag),
    .io_uop_wflag(slots_11_io_uop_wflag),
    .io_uop_prflag(slots_11_io_uop_prflag),
    .io_uop_pwflag(slots_11_io_uop_pwflag),
    .io_uop_pflag_busy(slots_11_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_11_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_11_io_uop_op1_sel),
    .io_uop_op2_sel(slots_11_io_uop_op2_sel),
    .io_uop_split_num(slots_11_io_uop_split_num),
    .io_uop_self_index(slots_11_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_11_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_11_io_uop_address_num),
    .io_uop_uopc(slots_11_io_uop_uopc),
    .io_uop_inst(slots_11_io_uop_inst),
    .io_uop_debug_inst(slots_11_io_uop_debug_inst),
    .io_uop_is_rvc(slots_11_io_uop_is_rvc),
    .io_uop_debug_pc(slots_11_io_uop_debug_pc),
    .io_uop_iq_type(slots_11_io_uop_iq_type),
    .io_uop_fu_code(slots_11_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_11_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_11_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_11_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_11_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_11_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_11_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_11_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_11_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_11_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_11_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_11_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_11_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_11_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_11_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_11_io_uop_is_br),
    .io_uop_is_jalr(slots_11_io_uop_is_jalr),
    .io_uop_is_jal(slots_11_io_uop_is_jal),
    .io_uop_is_sfb(slots_11_io_uop_is_sfb),
    .io_uop_br_mask(slots_11_io_uop_br_mask),
    .io_uop_br_tag(slots_11_io_uop_br_tag),
    .io_uop_ftq_idx(slots_11_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_11_io_uop_edge_inst),
    .io_uop_pc_lob(slots_11_io_uop_pc_lob),
    .io_uop_taken(slots_11_io_uop_taken),
    .io_uop_imm_packed(slots_11_io_uop_imm_packed),
    .io_uop_csr_addr(slots_11_io_uop_csr_addr),
    .io_uop_rob_idx(slots_11_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_11_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_11_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_11_io_uop_rxq_idx),
    .io_uop_pdst(slots_11_io_uop_pdst),
    .io_uop_prs1(slots_11_io_uop_prs1),
    .io_uop_prs2(slots_11_io_uop_prs2),
    .io_uop_prs3(slots_11_io_uop_prs3),
    .io_uop_ppred(slots_11_io_uop_ppred),
    .io_uop_prs1_busy(slots_11_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_11_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_11_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_11_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_11_io_uop_stale_pdst),
    .io_uop_exception(slots_11_io_uop_exception),
    .io_uop_exc_cause(slots_11_io_uop_exc_cause),
    .io_uop_bypassable(slots_11_io_uop_bypassable),
    .io_uop_mem_cmd(slots_11_io_uop_mem_cmd),
    .io_uop_mem_size(slots_11_io_uop_mem_size),
    .io_uop_mem_signed(slots_11_io_uop_mem_signed),
    .io_uop_is_fence(slots_11_io_uop_is_fence),
    .io_uop_is_fencei(slots_11_io_uop_is_fencei),
    .io_uop_is_amo(slots_11_io_uop_is_amo),
    .io_uop_uses_ldq(slots_11_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_11_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_11_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_11_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_11_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_11_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_11_io_uop_ldst),
    .io_uop_lrs1(slots_11_io_uop_lrs1),
    .io_uop_lrs2(slots_11_io_uop_lrs2),
    .io_uop_lrs3(slots_11_io_uop_lrs3),
    .io_uop_ldst_val(slots_11_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_11_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_11_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_11_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_11_io_uop_frs3_en),
    .io_uop_fp_val(slots_11_io_uop_fp_val),
    .io_uop_fp_single(slots_11_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_11_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_11_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_11_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_11_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_11_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_11_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_11_io_uop_debug_tsrc),
    .io_debug_p1(slots_11_io_debug_p1),
    .io_debug_p2(slots_11_io_debug_p2),
    .io_debug_p3(slots_11_io_debug_p3),
    .io_debug_ppred(slots_11_io_debug_ppred),
    .io_debug_state(slots_11_io_debug_state)
  );
  IssueSlot slots_12 ( // @[issue-unit.scala 157:73]
    .clock(slots_12_clock),
    .reset(slots_12_reset),
    .io_valid(slots_12_io_valid),
    .io_will_be_valid(slots_12_io_will_be_valid),
    .io_request(slots_12_io_request),
    .io_request_hp(slots_12_io_request_hp),
    .io_grant(slots_12_io_grant),
    .io_brupdate_b1_resolve_mask(slots_12_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_12_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_12_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_12_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_12_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_12_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_12_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_12_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_12_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_12_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_12_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_12_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_12_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_12_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_12_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_12_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_12_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_12_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_12_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_12_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_12_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_12_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_12_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_12_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_12_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_12_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_12_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_12_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_12_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_12_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_12_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_12_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_12_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_12_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_12_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_12_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_12_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_12_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_12_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_12_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_12_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_12_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_12_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_12_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_12_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_12_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_12_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_12_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_12_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_12_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_12_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_12_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_12_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_12_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_12_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_12_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_12_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_12_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_12_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_12_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_12_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_12_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_12_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_12_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_12_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_12_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_12_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_12_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_12_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_12_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_12_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_12_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_12_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_12_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_12_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_12_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_12_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_12_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_12_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_12_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_12_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_12_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_12_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_12_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_12_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_12_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_12_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_12_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_12_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_12_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_12_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_12_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_12_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_12_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_12_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_12_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_12_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_12_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_12_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_12_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_12_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_12_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_12_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_12_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_12_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_12_io_brupdate_b2_target_offset),
    .io_kill(slots_12_io_kill),
    .io_clear(slots_12_io_clear),
    .io_ldspec_miss(slots_12_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_12_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_12_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_12_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_12_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_12_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_12_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_12_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_12_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_12_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_12_io_wakeup_ports_1_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_12_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_12_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_12_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_12_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_12_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_12_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_12_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_12_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_12_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_12_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_12_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_12_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_12_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_12_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_12_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_12_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_12_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_12_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_12_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_12_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_12_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_12_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_12_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_12_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_12_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_12_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_12_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_12_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_12_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_12_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_12_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_12_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_12_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_12_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_12_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_12_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_12_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_12_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_12_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_12_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_12_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_12_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_12_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_12_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_12_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_12_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_12_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_12_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_12_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_12_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_12_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_12_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_12_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_12_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_12_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_12_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_12_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_12_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_12_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_12_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_12_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_12_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_12_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_12_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_12_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_12_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_12_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_12_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_12_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_12_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_12_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_12_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_12_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_12_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_12_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_12_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_12_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_12_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_12_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_12_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_12_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_12_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_12_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_12_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_12_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_12_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_12_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_12_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_12_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_12_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_12_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_12_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_12_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_12_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_12_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_12_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_12_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_12_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_12_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_12_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_12_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_12_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_12_io_out_uop_switch),
    .io_out_uop_switch_off(slots_12_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_12_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_12_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_12_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_12_io_out_uop_rflag),
    .io_out_uop_wflag(slots_12_io_out_uop_wflag),
    .io_out_uop_prflag(slots_12_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_12_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_12_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_12_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_12_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_12_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_12_io_out_uop_split_num),
    .io_out_uop_self_index(slots_12_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_12_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_12_io_out_uop_address_num),
    .io_out_uop_uopc(slots_12_io_out_uop_uopc),
    .io_out_uop_inst(slots_12_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_12_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_12_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_12_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_12_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_12_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_12_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_12_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_12_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_12_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_12_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_12_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_12_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_12_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_12_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_12_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_12_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_12_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_12_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_12_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_12_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_12_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_12_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_12_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_12_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_12_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_12_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_12_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_12_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_12_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_12_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_12_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_12_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_12_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_12_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_12_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_12_io_out_uop_pdst),
    .io_out_uop_prs1(slots_12_io_out_uop_prs1),
    .io_out_uop_prs2(slots_12_io_out_uop_prs2),
    .io_out_uop_prs3(slots_12_io_out_uop_prs3),
    .io_out_uop_ppred(slots_12_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_12_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_12_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_12_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_12_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_12_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_12_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_12_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_12_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_12_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_12_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_12_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_12_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_12_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_12_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_12_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_12_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_12_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_12_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_12_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_12_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_12_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_12_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_12_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_12_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_12_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_12_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_12_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_12_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_12_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_12_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_12_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_12_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_12_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_12_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_12_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_12_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_12_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_12_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_12_io_uop_switch),
    .io_uop_switch_off(slots_12_io_uop_switch_off),
    .io_uop_is_unicore(slots_12_io_uop_is_unicore),
    .io_uop_shift(slots_12_io_uop_shift),
    .io_uop_lrs3_rtype(slots_12_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_12_io_uop_rflag),
    .io_uop_wflag(slots_12_io_uop_wflag),
    .io_uop_prflag(slots_12_io_uop_prflag),
    .io_uop_pwflag(slots_12_io_uop_pwflag),
    .io_uop_pflag_busy(slots_12_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_12_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_12_io_uop_op1_sel),
    .io_uop_op2_sel(slots_12_io_uop_op2_sel),
    .io_uop_split_num(slots_12_io_uop_split_num),
    .io_uop_self_index(slots_12_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_12_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_12_io_uop_address_num),
    .io_uop_uopc(slots_12_io_uop_uopc),
    .io_uop_inst(slots_12_io_uop_inst),
    .io_uop_debug_inst(slots_12_io_uop_debug_inst),
    .io_uop_is_rvc(slots_12_io_uop_is_rvc),
    .io_uop_debug_pc(slots_12_io_uop_debug_pc),
    .io_uop_iq_type(slots_12_io_uop_iq_type),
    .io_uop_fu_code(slots_12_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_12_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_12_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_12_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_12_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_12_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_12_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_12_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_12_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_12_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_12_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_12_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_12_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_12_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_12_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_12_io_uop_is_br),
    .io_uop_is_jalr(slots_12_io_uop_is_jalr),
    .io_uop_is_jal(slots_12_io_uop_is_jal),
    .io_uop_is_sfb(slots_12_io_uop_is_sfb),
    .io_uop_br_mask(slots_12_io_uop_br_mask),
    .io_uop_br_tag(slots_12_io_uop_br_tag),
    .io_uop_ftq_idx(slots_12_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_12_io_uop_edge_inst),
    .io_uop_pc_lob(slots_12_io_uop_pc_lob),
    .io_uop_taken(slots_12_io_uop_taken),
    .io_uop_imm_packed(slots_12_io_uop_imm_packed),
    .io_uop_csr_addr(slots_12_io_uop_csr_addr),
    .io_uop_rob_idx(slots_12_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_12_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_12_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_12_io_uop_rxq_idx),
    .io_uop_pdst(slots_12_io_uop_pdst),
    .io_uop_prs1(slots_12_io_uop_prs1),
    .io_uop_prs2(slots_12_io_uop_prs2),
    .io_uop_prs3(slots_12_io_uop_prs3),
    .io_uop_ppred(slots_12_io_uop_ppred),
    .io_uop_prs1_busy(slots_12_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_12_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_12_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_12_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_12_io_uop_stale_pdst),
    .io_uop_exception(slots_12_io_uop_exception),
    .io_uop_exc_cause(slots_12_io_uop_exc_cause),
    .io_uop_bypassable(slots_12_io_uop_bypassable),
    .io_uop_mem_cmd(slots_12_io_uop_mem_cmd),
    .io_uop_mem_size(slots_12_io_uop_mem_size),
    .io_uop_mem_signed(slots_12_io_uop_mem_signed),
    .io_uop_is_fence(slots_12_io_uop_is_fence),
    .io_uop_is_fencei(slots_12_io_uop_is_fencei),
    .io_uop_is_amo(slots_12_io_uop_is_amo),
    .io_uop_uses_ldq(slots_12_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_12_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_12_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_12_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_12_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_12_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_12_io_uop_ldst),
    .io_uop_lrs1(slots_12_io_uop_lrs1),
    .io_uop_lrs2(slots_12_io_uop_lrs2),
    .io_uop_lrs3(slots_12_io_uop_lrs3),
    .io_uop_ldst_val(slots_12_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_12_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_12_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_12_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_12_io_uop_frs3_en),
    .io_uop_fp_val(slots_12_io_uop_fp_val),
    .io_uop_fp_single(slots_12_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_12_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_12_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_12_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_12_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_12_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_12_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_12_io_uop_debug_tsrc),
    .io_debug_p1(slots_12_io_debug_p1),
    .io_debug_p2(slots_12_io_debug_p2),
    .io_debug_p3(slots_12_io_debug_p3),
    .io_debug_ppred(slots_12_io_debug_ppred),
    .io_debug_state(slots_12_io_debug_state)
  );
  IssueSlot slots_13 ( // @[issue-unit.scala 157:73]
    .clock(slots_13_clock),
    .reset(slots_13_reset),
    .io_valid(slots_13_io_valid),
    .io_will_be_valid(slots_13_io_will_be_valid),
    .io_request(slots_13_io_request),
    .io_request_hp(slots_13_io_request_hp),
    .io_grant(slots_13_io_grant),
    .io_brupdate_b1_resolve_mask(slots_13_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_13_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_13_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_13_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_13_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_13_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_13_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_13_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_13_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_13_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_13_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_13_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_13_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_13_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_13_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_13_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_13_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_13_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_13_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_13_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_13_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_13_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_13_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_13_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_13_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_13_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_13_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_13_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_13_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_13_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_13_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_13_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_13_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_13_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_13_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_13_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_13_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_13_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_13_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_13_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_13_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_13_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_13_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_13_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_13_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_13_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_13_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_13_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_13_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_13_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_13_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_13_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_13_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_13_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_13_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_13_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_13_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_13_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_13_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_13_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_13_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_13_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_13_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_13_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_13_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_13_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_13_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_13_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_13_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_13_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_13_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_13_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_13_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_13_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_13_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_13_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_13_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_13_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_13_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_13_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_13_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_13_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_13_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_13_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_13_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_13_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_13_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_13_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_13_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_13_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_13_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_13_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_13_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_13_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_13_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_13_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_13_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_13_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_13_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_13_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_13_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_13_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_13_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_13_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_13_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_13_io_brupdate_b2_target_offset),
    .io_kill(slots_13_io_kill),
    .io_clear(slots_13_io_clear),
    .io_ldspec_miss(slots_13_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_13_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_13_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_13_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_13_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_13_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_13_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_13_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_13_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_13_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_13_io_wakeup_ports_1_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_13_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_13_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_13_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_13_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_13_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_13_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_13_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_13_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_13_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_13_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_13_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_13_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_13_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_13_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_13_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_13_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_13_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_13_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_13_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_13_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_13_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_13_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_13_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_13_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_13_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_13_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_13_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_13_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_13_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_13_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_13_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_13_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_13_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_13_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_13_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_13_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_13_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_13_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_13_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_13_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_13_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_13_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_13_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_13_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_13_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_13_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_13_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_13_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_13_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_13_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_13_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_13_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_13_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_13_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_13_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_13_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_13_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_13_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_13_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_13_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_13_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_13_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_13_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_13_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_13_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_13_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_13_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_13_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_13_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_13_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_13_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_13_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_13_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_13_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_13_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_13_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_13_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_13_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_13_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_13_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_13_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_13_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_13_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_13_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_13_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_13_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_13_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_13_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_13_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_13_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_13_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_13_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_13_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_13_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_13_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_13_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_13_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_13_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_13_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_13_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_13_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_13_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_13_io_out_uop_switch),
    .io_out_uop_switch_off(slots_13_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_13_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_13_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_13_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_13_io_out_uop_rflag),
    .io_out_uop_wflag(slots_13_io_out_uop_wflag),
    .io_out_uop_prflag(slots_13_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_13_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_13_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_13_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_13_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_13_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_13_io_out_uop_split_num),
    .io_out_uop_self_index(slots_13_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_13_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_13_io_out_uop_address_num),
    .io_out_uop_uopc(slots_13_io_out_uop_uopc),
    .io_out_uop_inst(slots_13_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_13_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_13_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_13_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_13_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_13_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_13_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_13_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_13_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_13_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_13_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_13_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_13_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_13_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_13_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_13_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_13_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_13_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_13_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_13_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_13_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_13_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_13_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_13_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_13_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_13_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_13_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_13_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_13_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_13_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_13_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_13_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_13_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_13_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_13_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_13_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_13_io_out_uop_pdst),
    .io_out_uop_prs1(slots_13_io_out_uop_prs1),
    .io_out_uop_prs2(slots_13_io_out_uop_prs2),
    .io_out_uop_prs3(slots_13_io_out_uop_prs3),
    .io_out_uop_ppred(slots_13_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_13_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_13_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_13_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_13_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_13_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_13_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_13_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_13_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_13_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_13_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_13_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_13_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_13_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_13_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_13_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_13_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_13_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_13_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_13_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_13_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_13_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_13_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_13_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_13_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_13_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_13_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_13_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_13_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_13_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_13_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_13_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_13_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_13_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_13_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_13_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_13_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_13_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_13_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_13_io_uop_switch),
    .io_uop_switch_off(slots_13_io_uop_switch_off),
    .io_uop_is_unicore(slots_13_io_uop_is_unicore),
    .io_uop_shift(slots_13_io_uop_shift),
    .io_uop_lrs3_rtype(slots_13_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_13_io_uop_rflag),
    .io_uop_wflag(slots_13_io_uop_wflag),
    .io_uop_prflag(slots_13_io_uop_prflag),
    .io_uop_pwflag(slots_13_io_uop_pwflag),
    .io_uop_pflag_busy(slots_13_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_13_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_13_io_uop_op1_sel),
    .io_uop_op2_sel(slots_13_io_uop_op2_sel),
    .io_uop_split_num(slots_13_io_uop_split_num),
    .io_uop_self_index(slots_13_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_13_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_13_io_uop_address_num),
    .io_uop_uopc(slots_13_io_uop_uopc),
    .io_uop_inst(slots_13_io_uop_inst),
    .io_uop_debug_inst(slots_13_io_uop_debug_inst),
    .io_uop_is_rvc(slots_13_io_uop_is_rvc),
    .io_uop_debug_pc(slots_13_io_uop_debug_pc),
    .io_uop_iq_type(slots_13_io_uop_iq_type),
    .io_uop_fu_code(slots_13_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_13_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_13_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_13_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_13_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_13_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_13_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_13_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_13_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_13_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_13_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_13_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_13_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_13_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_13_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_13_io_uop_is_br),
    .io_uop_is_jalr(slots_13_io_uop_is_jalr),
    .io_uop_is_jal(slots_13_io_uop_is_jal),
    .io_uop_is_sfb(slots_13_io_uop_is_sfb),
    .io_uop_br_mask(slots_13_io_uop_br_mask),
    .io_uop_br_tag(slots_13_io_uop_br_tag),
    .io_uop_ftq_idx(slots_13_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_13_io_uop_edge_inst),
    .io_uop_pc_lob(slots_13_io_uop_pc_lob),
    .io_uop_taken(slots_13_io_uop_taken),
    .io_uop_imm_packed(slots_13_io_uop_imm_packed),
    .io_uop_csr_addr(slots_13_io_uop_csr_addr),
    .io_uop_rob_idx(slots_13_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_13_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_13_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_13_io_uop_rxq_idx),
    .io_uop_pdst(slots_13_io_uop_pdst),
    .io_uop_prs1(slots_13_io_uop_prs1),
    .io_uop_prs2(slots_13_io_uop_prs2),
    .io_uop_prs3(slots_13_io_uop_prs3),
    .io_uop_ppred(slots_13_io_uop_ppred),
    .io_uop_prs1_busy(slots_13_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_13_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_13_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_13_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_13_io_uop_stale_pdst),
    .io_uop_exception(slots_13_io_uop_exception),
    .io_uop_exc_cause(slots_13_io_uop_exc_cause),
    .io_uop_bypassable(slots_13_io_uop_bypassable),
    .io_uop_mem_cmd(slots_13_io_uop_mem_cmd),
    .io_uop_mem_size(slots_13_io_uop_mem_size),
    .io_uop_mem_signed(slots_13_io_uop_mem_signed),
    .io_uop_is_fence(slots_13_io_uop_is_fence),
    .io_uop_is_fencei(slots_13_io_uop_is_fencei),
    .io_uop_is_amo(slots_13_io_uop_is_amo),
    .io_uop_uses_ldq(slots_13_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_13_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_13_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_13_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_13_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_13_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_13_io_uop_ldst),
    .io_uop_lrs1(slots_13_io_uop_lrs1),
    .io_uop_lrs2(slots_13_io_uop_lrs2),
    .io_uop_lrs3(slots_13_io_uop_lrs3),
    .io_uop_ldst_val(slots_13_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_13_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_13_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_13_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_13_io_uop_frs3_en),
    .io_uop_fp_val(slots_13_io_uop_fp_val),
    .io_uop_fp_single(slots_13_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_13_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_13_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_13_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_13_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_13_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_13_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_13_io_uop_debug_tsrc),
    .io_debug_p1(slots_13_io_debug_p1),
    .io_debug_p2(slots_13_io_debug_p2),
    .io_debug_p3(slots_13_io_debug_p3),
    .io_debug_ppred(slots_13_io_debug_ppred),
    .io_debug_state(slots_13_io_debug_state)
  );
  IssueSlot slots_14 ( // @[issue-unit.scala 157:73]
    .clock(slots_14_clock),
    .reset(slots_14_reset),
    .io_valid(slots_14_io_valid),
    .io_will_be_valid(slots_14_io_will_be_valid),
    .io_request(slots_14_io_request),
    .io_request_hp(slots_14_io_request_hp),
    .io_grant(slots_14_io_grant),
    .io_brupdate_b1_resolve_mask(slots_14_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_14_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_14_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_14_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_14_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_14_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_14_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_14_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_14_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_14_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_14_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_14_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_14_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_14_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_14_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_14_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_14_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_14_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_14_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_14_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_14_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_14_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_14_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_14_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_14_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_14_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_14_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_14_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_14_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_14_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_14_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_14_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_14_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_14_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_14_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_14_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_14_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_14_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_14_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_14_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_14_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_14_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_14_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_14_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_14_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_14_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_14_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_14_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_14_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_14_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_14_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_14_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_14_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_14_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_14_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_14_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_14_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_14_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_14_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_14_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_14_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_14_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_14_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_14_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_14_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_14_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_14_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_14_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_14_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_14_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_14_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_14_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_14_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_14_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_14_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_14_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_14_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_14_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_14_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_14_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_14_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_14_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_14_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_14_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_14_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_14_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_14_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_14_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_14_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_14_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_14_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_14_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_14_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_14_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_14_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_14_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_14_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_14_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_14_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_14_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_14_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_14_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_14_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_14_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_14_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_14_io_brupdate_b2_target_offset),
    .io_kill(slots_14_io_kill),
    .io_clear(slots_14_io_clear),
    .io_ldspec_miss(slots_14_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_14_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_14_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_14_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_14_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_14_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_14_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_14_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_14_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_14_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_14_io_wakeup_ports_1_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_14_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_14_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_14_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_14_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_14_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_14_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_14_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_14_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_14_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_14_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_14_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_14_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_14_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_14_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_14_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_14_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_14_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_14_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_14_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_14_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_14_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_14_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_14_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_14_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_14_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_14_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_14_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_14_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_14_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_14_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_14_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_14_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_14_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_14_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_14_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_14_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_14_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_14_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_14_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_14_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_14_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_14_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_14_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_14_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_14_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_14_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_14_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_14_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_14_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_14_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_14_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_14_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_14_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_14_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_14_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_14_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_14_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_14_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_14_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_14_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_14_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_14_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_14_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_14_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_14_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_14_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_14_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_14_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_14_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_14_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_14_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_14_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_14_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_14_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_14_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_14_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_14_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_14_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_14_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_14_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_14_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_14_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_14_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_14_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_14_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_14_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_14_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_14_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_14_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_14_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_14_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_14_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_14_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_14_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_14_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_14_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_14_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_14_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_14_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_14_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_14_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_14_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_14_io_out_uop_switch),
    .io_out_uop_switch_off(slots_14_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_14_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_14_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_14_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_14_io_out_uop_rflag),
    .io_out_uop_wflag(slots_14_io_out_uop_wflag),
    .io_out_uop_prflag(slots_14_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_14_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_14_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_14_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_14_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_14_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_14_io_out_uop_split_num),
    .io_out_uop_self_index(slots_14_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_14_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_14_io_out_uop_address_num),
    .io_out_uop_uopc(slots_14_io_out_uop_uopc),
    .io_out_uop_inst(slots_14_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_14_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_14_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_14_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_14_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_14_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_14_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_14_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_14_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_14_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_14_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_14_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_14_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_14_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_14_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_14_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_14_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_14_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_14_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_14_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_14_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_14_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_14_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_14_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_14_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_14_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_14_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_14_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_14_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_14_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_14_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_14_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_14_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_14_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_14_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_14_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_14_io_out_uop_pdst),
    .io_out_uop_prs1(slots_14_io_out_uop_prs1),
    .io_out_uop_prs2(slots_14_io_out_uop_prs2),
    .io_out_uop_prs3(slots_14_io_out_uop_prs3),
    .io_out_uop_ppred(slots_14_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_14_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_14_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_14_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_14_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_14_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_14_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_14_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_14_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_14_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_14_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_14_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_14_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_14_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_14_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_14_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_14_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_14_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_14_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_14_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_14_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_14_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_14_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_14_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_14_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_14_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_14_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_14_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_14_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_14_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_14_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_14_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_14_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_14_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_14_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_14_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_14_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_14_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_14_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_14_io_uop_switch),
    .io_uop_switch_off(slots_14_io_uop_switch_off),
    .io_uop_is_unicore(slots_14_io_uop_is_unicore),
    .io_uop_shift(slots_14_io_uop_shift),
    .io_uop_lrs3_rtype(slots_14_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_14_io_uop_rflag),
    .io_uop_wflag(slots_14_io_uop_wflag),
    .io_uop_prflag(slots_14_io_uop_prflag),
    .io_uop_pwflag(slots_14_io_uop_pwflag),
    .io_uop_pflag_busy(slots_14_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_14_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_14_io_uop_op1_sel),
    .io_uop_op2_sel(slots_14_io_uop_op2_sel),
    .io_uop_split_num(slots_14_io_uop_split_num),
    .io_uop_self_index(slots_14_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_14_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_14_io_uop_address_num),
    .io_uop_uopc(slots_14_io_uop_uopc),
    .io_uop_inst(slots_14_io_uop_inst),
    .io_uop_debug_inst(slots_14_io_uop_debug_inst),
    .io_uop_is_rvc(slots_14_io_uop_is_rvc),
    .io_uop_debug_pc(slots_14_io_uop_debug_pc),
    .io_uop_iq_type(slots_14_io_uop_iq_type),
    .io_uop_fu_code(slots_14_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_14_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_14_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_14_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_14_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_14_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_14_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_14_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_14_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_14_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_14_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_14_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_14_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_14_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_14_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_14_io_uop_is_br),
    .io_uop_is_jalr(slots_14_io_uop_is_jalr),
    .io_uop_is_jal(slots_14_io_uop_is_jal),
    .io_uop_is_sfb(slots_14_io_uop_is_sfb),
    .io_uop_br_mask(slots_14_io_uop_br_mask),
    .io_uop_br_tag(slots_14_io_uop_br_tag),
    .io_uop_ftq_idx(slots_14_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_14_io_uop_edge_inst),
    .io_uop_pc_lob(slots_14_io_uop_pc_lob),
    .io_uop_taken(slots_14_io_uop_taken),
    .io_uop_imm_packed(slots_14_io_uop_imm_packed),
    .io_uop_csr_addr(slots_14_io_uop_csr_addr),
    .io_uop_rob_idx(slots_14_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_14_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_14_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_14_io_uop_rxq_idx),
    .io_uop_pdst(slots_14_io_uop_pdst),
    .io_uop_prs1(slots_14_io_uop_prs1),
    .io_uop_prs2(slots_14_io_uop_prs2),
    .io_uop_prs3(slots_14_io_uop_prs3),
    .io_uop_ppred(slots_14_io_uop_ppred),
    .io_uop_prs1_busy(slots_14_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_14_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_14_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_14_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_14_io_uop_stale_pdst),
    .io_uop_exception(slots_14_io_uop_exception),
    .io_uop_exc_cause(slots_14_io_uop_exc_cause),
    .io_uop_bypassable(slots_14_io_uop_bypassable),
    .io_uop_mem_cmd(slots_14_io_uop_mem_cmd),
    .io_uop_mem_size(slots_14_io_uop_mem_size),
    .io_uop_mem_signed(slots_14_io_uop_mem_signed),
    .io_uop_is_fence(slots_14_io_uop_is_fence),
    .io_uop_is_fencei(slots_14_io_uop_is_fencei),
    .io_uop_is_amo(slots_14_io_uop_is_amo),
    .io_uop_uses_ldq(slots_14_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_14_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_14_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_14_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_14_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_14_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_14_io_uop_ldst),
    .io_uop_lrs1(slots_14_io_uop_lrs1),
    .io_uop_lrs2(slots_14_io_uop_lrs2),
    .io_uop_lrs3(slots_14_io_uop_lrs3),
    .io_uop_ldst_val(slots_14_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_14_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_14_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_14_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_14_io_uop_frs3_en),
    .io_uop_fp_val(slots_14_io_uop_fp_val),
    .io_uop_fp_single(slots_14_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_14_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_14_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_14_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_14_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_14_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_14_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_14_io_uop_debug_tsrc),
    .io_debug_p1(slots_14_io_debug_p1),
    .io_debug_p2(slots_14_io_debug_p2),
    .io_debug_p3(slots_14_io_debug_p3),
    .io_debug_ppred(slots_14_io_debug_ppred),
    .io_debug_state(slots_14_io_debug_state)
  );
  IssueSlot slots_15 ( // @[issue-unit.scala 157:73]
    .clock(slots_15_clock),
    .reset(slots_15_reset),
    .io_valid(slots_15_io_valid),
    .io_will_be_valid(slots_15_io_will_be_valid),
    .io_request(slots_15_io_request),
    .io_request_hp(slots_15_io_request_hp),
    .io_grant(slots_15_io_grant),
    .io_brupdate_b1_resolve_mask(slots_15_io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask(slots_15_io_brupdate_b1_mispredict_mask),
    .io_brupdate_b2_uop_switch(slots_15_io_brupdate_b2_uop_switch),
    .io_brupdate_b2_uop_switch_off(slots_15_io_brupdate_b2_uop_switch_off),
    .io_brupdate_b2_uop_is_unicore(slots_15_io_brupdate_b2_uop_is_unicore),
    .io_brupdate_b2_uop_shift(slots_15_io_brupdate_b2_uop_shift),
    .io_brupdate_b2_uop_lrs3_rtype(slots_15_io_brupdate_b2_uop_lrs3_rtype),
    .io_brupdate_b2_uop_rflag(slots_15_io_brupdate_b2_uop_rflag),
    .io_brupdate_b2_uop_wflag(slots_15_io_brupdate_b2_uop_wflag),
    .io_brupdate_b2_uop_prflag(slots_15_io_brupdate_b2_uop_prflag),
    .io_brupdate_b2_uop_pwflag(slots_15_io_brupdate_b2_uop_pwflag),
    .io_brupdate_b2_uop_pflag_busy(slots_15_io_brupdate_b2_uop_pflag_busy),
    .io_brupdate_b2_uop_stale_pflag(slots_15_io_brupdate_b2_uop_stale_pflag),
    .io_brupdate_b2_uop_op1_sel(slots_15_io_brupdate_b2_uop_op1_sel),
    .io_brupdate_b2_uop_op2_sel(slots_15_io_brupdate_b2_uop_op2_sel),
    .io_brupdate_b2_uop_split_num(slots_15_io_brupdate_b2_uop_split_num),
    .io_brupdate_b2_uop_self_index(slots_15_io_brupdate_b2_uop_self_index),
    .io_brupdate_b2_uop_rob_inst_idx(slots_15_io_brupdate_b2_uop_rob_inst_idx),
    .io_brupdate_b2_uop_address_num(slots_15_io_brupdate_b2_uop_address_num),
    .io_brupdate_b2_uop_uopc(slots_15_io_brupdate_b2_uop_uopc),
    .io_brupdate_b2_uop_inst(slots_15_io_brupdate_b2_uop_inst),
    .io_brupdate_b2_uop_debug_inst(slots_15_io_brupdate_b2_uop_debug_inst),
    .io_brupdate_b2_uop_is_rvc(slots_15_io_brupdate_b2_uop_is_rvc),
    .io_brupdate_b2_uop_debug_pc(slots_15_io_brupdate_b2_uop_debug_pc),
    .io_brupdate_b2_uop_iq_type(slots_15_io_brupdate_b2_uop_iq_type),
    .io_brupdate_b2_uop_fu_code(slots_15_io_brupdate_b2_uop_fu_code),
    .io_brupdate_b2_uop_ctrl_br_type(slots_15_io_brupdate_b2_uop_ctrl_br_type),
    .io_brupdate_b2_uop_ctrl_op1_sel(slots_15_io_brupdate_b2_uop_ctrl_op1_sel),
    .io_brupdate_b2_uop_ctrl_op2_sel(slots_15_io_brupdate_b2_uop_ctrl_op2_sel),
    .io_brupdate_b2_uop_ctrl_imm_sel(slots_15_io_brupdate_b2_uop_ctrl_imm_sel),
    .io_brupdate_b2_uop_ctrl_op_fcn(slots_15_io_brupdate_b2_uop_ctrl_op_fcn),
    .io_brupdate_b2_uop_ctrl_fcn_dw(slots_15_io_brupdate_b2_uop_ctrl_fcn_dw),
    .io_brupdate_b2_uop_ctrl_csr_cmd(slots_15_io_brupdate_b2_uop_ctrl_csr_cmd),
    .io_brupdate_b2_uop_ctrl_is_load(slots_15_io_brupdate_b2_uop_ctrl_is_load),
    .io_brupdate_b2_uop_ctrl_is_sta(slots_15_io_brupdate_b2_uop_ctrl_is_sta),
    .io_brupdate_b2_uop_ctrl_is_std(slots_15_io_brupdate_b2_uop_ctrl_is_std),
    .io_brupdate_b2_uop_ctrl_op3_sel(slots_15_io_brupdate_b2_uop_ctrl_op3_sel),
    .io_brupdate_b2_uop_iw_state(slots_15_io_brupdate_b2_uop_iw_state),
    .io_brupdate_b2_uop_iw_p1_poisoned(slots_15_io_brupdate_b2_uop_iw_p1_poisoned),
    .io_brupdate_b2_uop_iw_p2_poisoned(slots_15_io_brupdate_b2_uop_iw_p2_poisoned),
    .io_brupdate_b2_uop_is_br(slots_15_io_brupdate_b2_uop_is_br),
    .io_brupdate_b2_uop_is_jalr(slots_15_io_brupdate_b2_uop_is_jalr),
    .io_brupdate_b2_uop_is_jal(slots_15_io_brupdate_b2_uop_is_jal),
    .io_brupdate_b2_uop_is_sfb(slots_15_io_brupdate_b2_uop_is_sfb),
    .io_brupdate_b2_uop_br_mask(slots_15_io_brupdate_b2_uop_br_mask),
    .io_brupdate_b2_uop_br_tag(slots_15_io_brupdate_b2_uop_br_tag),
    .io_brupdate_b2_uop_ftq_idx(slots_15_io_brupdate_b2_uop_ftq_idx),
    .io_brupdate_b2_uop_edge_inst(slots_15_io_brupdate_b2_uop_edge_inst),
    .io_brupdate_b2_uop_pc_lob(slots_15_io_brupdate_b2_uop_pc_lob),
    .io_brupdate_b2_uop_taken(slots_15_io_brupdate_b2_uop_taken),
    .io_brupdate_b2_uop_imm_packed(slots_15_io_brupdate_b2_uop_imm_packed),
    .io_brupdate_b2_uop_csr_addr(slots_15_io_brupdate_b2_uop_csr_addr),
    .io_brupdate_b2_uop_rob_idx(slots_15_io_brupdate_b2_uop_rob_idx),
    .io_brupdate_b2_uop_ldq_idx(slots_15_io_brupdate_b2_uop_ldq_idx),
    .io_brupdate_b2_uop_stq_idx(slots_15_io_brupdate_b2_uop_stq_idx),
    .io_brupdate_b2_uop_rxq_idx(slots_15_io_brupdate_b2_uop_rxq_idx),
    .io_brupdate_b2_uop_pdst(slots_15_io_brupdate_b2_uop_pdst),
    .io_brupdate_b2_uop_prs1(slots_15_io_brupdate_b2_uop_prs1),
    .io_brupdate_b2_uop_prs2(slots_15_io_brupdate_b2_uop_prs2),
    .io_brupdate_b2_uop_prs3(slots_15_io_brupdate_b2_uop_prs3),
    .io_brupdate_b2_uop_ppred(slots_15_io_brupdate_b2_uop_ppred),
    .io_brupdate_b2_uop_prs1_busy(slots_15_io_brupdate_b2_uop_prs1_busy),
    .io_brupdate_b2_uop_prs2_busy(slots_15_io_brupdate_b2_uop_prs2_busy),
    .io_brupdate_b2_uop_prs3_busy(slots_15_io_brupdate_b2_uop_prs3_busy),
    .io_brupdate_b2_uop_ppred_busy(slots_15_io_brupdate_b2_uop_ppred_busy),
    .io_brupdate_b2_uop_stale_pdst(slots_15_io_brupdate_b2_uop_stale_pdst),
    .io_brupdate_b2_uop_exception(slots_15_io_brupdate_b2_uop_exception),
    .io_brupdate_b2_uop_exc_cause(slots_15_io_brupdate_b2_uop_exc_cause),
    .io_brupdate_b2_uop_bypassable(slots_15_io_brupdate_b2_uop_bypassable),
    .io_brupdate_b2_uop_mem_cmd(slots_15_io_brupdate_b2_uop_mem_cmd),
    .io_brupdate_b2_uop_mem_size(slots_15_io_brupdate_b2_uop_mem_size),
    .io_brupdate_b2_uop_mem_signed(slots_15_io_brupdate_b2_uop_mem_signed),
    .io_brupdate_b2_uop_is_fence(slots_15_io_brupdate_b2_uop_is_fence),
    .io_brupdate_b2_uop_is_fencei(slots_15_io_brupdate_b2_uop_is_fencei),
    .io_brupdate_b2_uop_is_amo(slots_15_io_brupdate_b2_uop_is_amo),
    .io_brupdate_b2_uop_uses_ldq(slots_15_io_brupdate_b2_uop_uses_ldq),
    .io_brupdate_b2_uop_uses_stq(slots_15_io_brupdate_b2_uop_uses_stq),
    .io_brupdate_b2_uop_is_sys_pc2epc(slots_15_io_brupdate_b2_uop_is_sys_pc2epc),
    .io_brupdate_b2_uop_is_unique(slots_15_io_brupdate_b2_uop_is_unique),
    .io_brupdate_b2_uop_flush_on_commit(slots_15_io_brupdate_b2_uop_flush_on_commit),
    .io_brupdate_b2_uop_ldst_is_rs1(slots_15_io_brupdate_b2_uop_ldst_is_rs1),
    .io_brupdate_b2_uop_ldst(slots_15_io_brupdate_b2_uop_ldst),
    .io_brupdate_b2_uop_lrs1(slots_15_io_brupdate_b2_uop_lrs1),
    .io_brupdate_b2_uop_lrs2(slots_15_io_brupdate_b2_uop_lrs2),
    .io_brupdate_b2_uop_lrs3(slots_15_io_brupdate_b2_uop_lrs3),
    .io_brupdate_b2_uop_ldst_val(slots_15_io_brupdate_b2_uop_ldst_val),
    .io_brupdate_b2_uop_dst_rtype(slots_15_io_brupdate_b2_uop_dst_rtype),
    .io_brupdate_b2_uop_lrs1_rtype(slots_15_io_brupdate_b2_uop_lrs1_rtype),
    .io_brupdate_b2_uop_lrs2_rtype(slots_15_io_brupdate_b2_uop_lrs2_rtype),
    .io_brupdate_b2_uop_frs3_en(slots_15_io_brupdate_b2_uop_frs3_en),
    .io_brupdate_b2_uop_fp_val(slots_15_io_brupdate_b2_uop_fp_val),
    .io_brupdate_b2_uop_fp_single(slots_15_io_brupdate_b2_uop_fp_single),
    .io_brupdate_b2_uop_xcpt_pf_if(slots_15_io_brupdate_b2_uop_xcpt_pf_if),
    .io_brupdate_b2_uop_xcpt_ae_if(slots_15_io_brupdate_b2_uop_xcpt_ae_if),
    .io_brupdate_b2_uop_xcpt_ma_if(slots_15_io_brupdate_b2_uop_xcpt_ma_if),
    .io_brupdate_b2_uop_bp_debug_if(slots_15_io_brupdate_b2_uop_bp_debug_if),
    .io_brupdate_b2_uop_bp_xcpt_if(slots_15_io_brupdate_b2_uop_bp_xcpt_if),
    .io_brupdate_b2_uop_debug_fsrc(slots_15_io_brupdate_b2_uop_debug_fsrc),
    .io_brupdate_b2_uop_debug_tsrc(slots_15_io_brupdate_b2_uop_debug_tsrc),
    .io_brupdate_b2_valid(slots_15_io_brupdate_b2_valid),
    .io_brupdate_b2_mispredict(slots_15_io_brupdate_b2_mispredict),
    .io_brupdate_b2_taken(slots_15_io_brupdate_b2_taken),
    .io_brupdate_b2_cfi_type(slots_15_io_brupdate_b2_cfi_type),
    .io_brupdate_b2_pc_sel(slots_15_io_brupdate_b2_pc_sel),
    .io_brupdate_b2_jalr_target(slots_15_io_brupdate_b2_jalr_target),
    .io_brupdate_b2_target_offset(slots_15_io_brupdate_b2_target_offset),
    .io_kill(slots_15_io_kill),
    .io_clear(slots_15_io_clear),
    .io_ldspec_miss(slots_15_io_ldspec_miss),
    .io_wakeup_ports_0_valid(slots_15_io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst(slots_15_io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_0_bits_poisoned(slots_15_io_wakeup_ports_0_bits_poisoned),
    .io_wakeup_ports_0_bits_pwflag(slots_15_io_wakeup_ports_0_bits_pwflag),
    .io_wakeup_ports_0_bits_flag_valid(slots_15_io_wakeup_ports_0_bits_flag_valid),
    .io_wakeup_ports_1_valid(slots_15_io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst(slots_15_io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_1_bits_poisoned(slots_15_io_wakeup_ports_1_bits_poisoned),
    .io_wakeup_ports_1_bits_pwflag(slots_15_io_wakeup_ports_1_bits_pwflag),
    .io_wakeup_ports_1_bits_flag_valid(slots_15_io_wakeup_ports_1_bits_flag_valid),
    .io_pred_wakeup_port_valid(slots_15_io_pred_wakeup_port_valid),
    .io_pred_wakeup_port_bits(slots_15_io_pred_wakeup_port_bits),
    .io_spec_ld_wakeup_0_valid(slots_15_io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits(slots_15_io_spec_ld_wakeup_0_bits),
    .io_in_uop_valid(slots_15_io_in_uop_valid),
    .io_in_uop_bits_switch(slots_15_io_in_uop_bits_switch),
    .io_in_uop_bits_switch_off(slots_15_io_in_uop_bits_switch_off),
    .io_in_uop_bits_is_unicore(slots_15_io_in_uop_bits_is_unicore),
    .io_in_uop_bits_shift(slots_15_io_in_uop_bits_shift),
    .io_in_uop_bits_lrs3_rtype(slots_15_io_in_uop_bits_lrs3_rtype),
    .io_in_uop_bits_rflag(slots_15_io_in_uop_bits_rflag),
    .io_in_uop_bits_wflag(slots_15_io_in_uop_bits_wflag),
    .io_in_uop_bits_prflag(slots_15_io_in_uop_bits_prflag),
    .io_in_uop_bits_pwflag(slots_15_io_in_uop_bits_pwflag),
    .io_in_uop_bits_pflag_busy(slots_15_io_in_uop_bits_pflag_busy),
    .io_in_uop_bits_stale_pflag(slots_15_io_in_uop_bits_stale_pflag),
    .io_in_uop_bits_op1_sel(slots_15_io_in_uop_bits_op1_sel),
    .io_in_uop_bits_op2_sel(slots_15_io_in_uop_bits_op2_sel),
    .io_in_uop_bits_split_num(slots_15_io_in_uop_bits_split_num),
    .io_in_uop_bits_self_index(slots_15_io_in_uop_bits_self_index),
    .io_in_uop_bits_rob_inst_idx(slots_15_io_in_uop_bits_rob_inst_idx),
    .io_in_uop_bits_address_num(slots_15_io_in_uop_bits_address_num),
    .io_in_uop_bits_uopc(slots_15_io_in_uop_bits_uopc),
    .io_in_uop_bits_inst(slots_15_io_in_uop_bits_inst),
    .io_in_uop_bits_debug_inst(slots_15_io_in_uop_bits_debug_inst),
    .io_in_uop_bits_is_rvc(slots_15_io_in_uop_bits_is_rvc),
    .io_in_uop_bits_debug_pc(slots_15_io_in_uop_bits_debug_pc),
    .io_in_uop_bits_iq_type(slots_15_io_in_uop_bits_iq_type),
    .io_in_uop_bits_fu_code(slots_15_io_in_uop_bits_fu_code),
    .io_in_uop_bits_ctrl_br_type(slots_15_io_in_uop_bits_ctrl_br_type),
    .io_in_uop_bits_ctrl_op1_sel(slots_15_io_in_uop_bits_ctrl_op1_sel),
    .io_in_uop_bits_ctrl_op2_sel(slots_15_io_in_uop_bits_ctrl_op2_sel),
    .io_in_uop_bits_ctrl_imm_sel(slots_15_io_in_uop_bits_ctrl_imm_sel),
    .io_in_uop_bits_ctrl_op_fcn(slots_15_io_in_uop_bits_ctrl_op_fcn),
    .io_in_uop_bits_ctrl_fcn_dw(slots_15_io_in_uop_bits_ctrl_fcn_dw),
    .io_in_uop_bits_ctrl_csr_cmd(slots_15_io_in_uop_bits_ctrl_csr_cmd),
    .io_in_uop_bits_ctrl_is_load(slots_15_io_in_uop_bits_ctrl_is_load),
    .io_in_uop_bits_ctrl_is_sta(slots_15_io_in_uop_bits_ctrl_is_sta),
    .io_in_uop_bits_ctrl_is_std(slots_15_io_in_uop_bits_ctrl_is_std),
    .io_in_uop_bits_ctrl_op3_sel(slots_15_io_in_uop_bits_ctrl_op3_sel),
    .io_in_uop_bits_iw_state(slots_15_io_in_uop_bits_iw_state),
    .io_in_uop_bits_iw_p1_poisoned(slots_15_io_in_uop_bits_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned(slots_15_io_in_uop_bits_iw_p2_poisoned),
    .io_in_uop_bits_is_br(slots_15_io_in_uop_bits_is_br),
    .io_in_uop_bits_is_jalr(slots_15_io_in_uop_bits_is_jalr),
    .io_in_uop_bits_is_jal(slots_15_io_in_uop_bits_is_jal),
    .io_in_uop_bits_is_sfb(slots_15_io_in_uop_bits_is_sfb),
    .io_in_uop_bits_br_mask(slots_15_io_in_uop_bits_br_mask),
    .io_in_uop_bits_br_tag(slots_15_io_in_uop_bits_br_tag),
    .io_in_uop_bits_ftq_idx(slots_15_io_in_uop_bits_ftq_idx),
    .io_in_uop_bits_edge_inst(slots_15_io_in_uop_bits_edge_inst),
    .io_in_uop_bits_pc_lob(slots_15_io_in_uop_bits_pc_lob),
    .io_in_uop_bits_taken(slots_15_io_in_uop_bits_taken),
    .io_in_uop_bits_imm_packed(slots_15_io_in_uop_bits_imm_packed),
    .io_in_uop_bits_csr_addr(slots_15_io_in_uop_bits_csr_addr),
    .io_in_uop_bits_rob_idx(slots_15_io_in_uop_bits_rob_idx),
    .io_in_uop_bits_ldq_idx(slots_15_io_in_uop_bits_ldq_idx),
    .io_in_uop_bits_stq_idx(slots_15_io_in_uop_bits_stq_idx),
    .io_in_uop_bits_rxq_idx(slots_15_io_in_uop_bits_rxq_idx),
    .io_in_uop_bits_pdst(slots_15_io_in_uop_bits_pdst),
    .io_in_uop_bits_prs1(slots_15_io_in_uop_bits_prs1),
    .io_in_uop_bits_prs2(slots_15_io_in_uop_bits_prs2),
    .io_in_uop_bits_prs3(slots_15_io_in_uop_bits_prs3),
    .io_in_uop_bits_ppred(slots_15_io_in_uop_bits_ppred),
    .io_in_uop_bits_prs1_busy(slots_15_io_in_uop_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy(slots_15_io_in_uop_bits_prs2_busy),
    .io_in_uop_bits_prs3_busy(slots_15_io_in_uop_bits_prs3_busy),
    .io_in_uop_bits_ppred_busy(slots_15_io_in_uop_bits_ppred_busy),
    .io_in_uop_bits_stale_pdst(slots_15_io_in_uop_bits_stale_pdst),
    .io_in_uop_bits_exception(slots_15_io_in_uop_bits_exception),
    .io_in_uop_bits_exc_cause(slots_15_io_in_uop_bits_exc_cause),
    .io_in_uop_bits_bypassable(slots_15_io_in_uop_bits_bypassable),
    .io_in_uop_bits_mem_cmd(slots_15_io_in_uop_bits_mem_cmd),
    .io_in_uop_bits_mem_size(slots_15_io_in_uop_bits_mem_size),
    .io_in_uop_bits_mem_signed(slots_15_io_in_uop_bits_mem_signed),
    .io_in_uop_bits_is_fence(slots_15_io_in_uop_bits_is_fence),
    .io_in_uop_bits_is_fencei(slots_15_io_in_uop_bits_is_fencei),
    .io_in_uop_bits_is_amo(slots_15_io_in_uop_bits_is_amo),
    .io_in_uop_bits_uses_ldq(slots_15_io_in_uop_bits_uses_ldq),
    .io_in_uop_bits_uses_stq(slots_15_io_in_uop_bits_uses_stq),
    .io_in_uop_bits_is_sys_pc2epc(slots_15_io_in_uop_bits_is_sys_pc2epc),
    .io_in_uop_bits_is_unique(slots_15_io_in_uop_bits_is_unique),
    .io_in_uop_bits_flush_on_commit(slots_15_io_in_uop_bits_flush_on_commit),
    .io_in_uop_bits_ldst_is_rs1(slots_15_io_in_uop_bits_ldst_is_rs1),
    .io_in_uop_bits_ldst(slots_15_io_in_uop_bits_ldst),
    .io_in_uop_bits_lrs1(slots_15_io_in_uop_bits_lrs1),
    .io_in_uop_bits_lrs2(slots_15_io_in_uop_bits_lrs2),
    .io_in_uop_bits_lrs3(slots_15_io_in_uop_bits_lrs3),
    .io_in_uop_bits_ldst_val(slots_15_io_in_uop_bits_ldst_val),
    .io_in_uop_bits_dst_rtype(slots_15_io_in_uop_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype(slots_15_io_in_uop_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype(slots_15_io_in_uop_bits_lrs2_rtype),
    .io_in_uop_bits_frs3_en(slots_15_io_in_uop_bits_frs3_en),
    .io_in_uop_bits_fp_val(slots_15_io_in_uop_bits_fp_val),
    .io_in_uop_bits_fp_single(slots_15_io_in_uop_bits_fp_single),
    .io_in_uop_bits_xcpt_pf_if(slots_15_io_in_uop_bits_xcpt_pf_if),
    .io_in_uop_bits_xcpt_ae_if(slots_15_io_in_uop_bits_xcpt_ae_if),
    .io_in_uop_bits_xcpt_ma_if(slots_15_io_in_uop_bits_xcpt_ma_if),
    .io_in_uop_bits_bp_debug_if(slots_15_io_in_uop_bits_bp_debug_if),
    .io_in_uop_bits_bp_xcpt_if(slots_15_io_in_uop_bits_bp_xcpt_if),
    .io_in_uop_bits_debug_fsrc(slots_15_io_in_uop_bits_debug_fsrc),
    .io_in_uop_bits_debug_tsrc(slots_15_io_in_uop_bits_debug_tsrc),
    .io_out_uop_switch(slots_15_io_out_uop_switch),
    .io_out_uop_switch_off(slots_15_io_out_uop_switch_off),
    .io_out_uop_is_unicore(slots_15_io_out_uop_is_unicore),
    .io_out_uop_shift(slots_15_io_out_uop_shift),
    .io_out_uop_lrs3_rtype(slots_15_io_out_uop_lrs3_rtype),
    .io_out_uop_rflag(slots_15_io_out_uop_rflag),
    .io_out_uop_wflag(slots_15_io_out_uop_wflag),
    .io_out_uop_prflag(slots_15_io_out_uop_prflag),
    .io_out_uop_pwflag(slots_15_io_out_uop_pwflag),
    .io_out_uop_pflag_busy(slots_15_io_out_uop_pflag_busy),
    .io_out_uop_stale_pflag(slots_15_io_out_uop_stale_pflag),
    .io_out_uop_op1_sel(slots_15_io_out_uop_op1_sel),
    .io_out_uop_op2_sel(slots_15_io_out_uop_op2_sel),
    .io_out_uop_split_num(slots_15_io_out_uop_split_num),
    .io_out_uop_self_index(slots_15_io_out_uop_self_index),
    .io_out_uop_rob_inst_idx(slots_15_io_out_uop_rob_inst_idx),
    .io_out_uop_address_num(slots_15_io_out_uop_address_num),
    .io_out_uop_uopc(slots_15_io_out_uop_uopc),
    .io_out_uop_inst(slots_15_io_out_uop_inst),
    .io_out_uop_debug_inst(slots_15_io_out_uop_debug_inst),
    .io_out_uop_is_rvc(slots_15_io_out_uop_is_rvc),
    .io_out_uop_debug_pc(slots_15_io_out_uop_debug_pc),
    .io_out_uop_iq_type(slots_15_io_out_uop_iq_type),
    .io_out_uop_fu_code(slots_15_io_out_uop_fu_code),
    .io_out_uop_ctrl_br_type(slots_15_io_out_uop_ctrl_br_type),
    .io_out_uop_ctrl_op1_sel(slots_15_io_out_uop_ctrl_op1_sel),
    .io_out_uop_ctrl_op2_sel(slots_15_io_out_uop_ctrl_op2_sel),
    .io_out_uop_ctrl_imm_sel(slots_15_io_out_uop_ctrl_imm_sel),
    .io_out_uop_ctrl_op_fcn(slots_15_io_out_uop_ctrl_op_fcn),
    .io_out_uop_ctrl_fcn_dw(slots_15_io_out_uop_ctrl_fcn_dw),
    .io_out_uop_ctrl_csr_cmd(slots_15_io_out_uop_ctrl_csr_cmd),
    .io_out_uop_ctrl_is_load(slots_15_io_out_uop_ctrl_is_load),
    .io_out_uop_ctrl_is_sta(slots_15_io_out_uop_ctrl_is_sta),
    .io_out_uop_ctrl_is_std(slots_15_io_out_uop_ctrl_is_std),
    .io_out_uop_ctrl_op3_sel(slots_15_io_out_uop_ctrl_op3_sel),
    .io_out_uop_iw_state(slots_15_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned(slots_15_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned(slots_15_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br(slots_15_io_out_uop_is_br),
    .io_out_uop_is_jalr(slots_15_io_out_uop_is_jalr),
    .io_out_uop_is_jal(slots_15_io_out_uop_is_jal),
    .io_out_uop_is_sfb(slots_15_io_out_uop_is_sfb),
    .io_out_uop_br_mask(slots_15_io_out_uop_br_mask),
    .io_out_uop_br_tag(slots_15_io_out_uop_br_tag),
    .io_out_uop_ftq_idx(slots_15_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst(slots_15_io_out_uop_edge_inst),
    .io_out_uop_pc_lob(slots_15_io_out_uop_pc_lob),
    .io_out_uop_taken(slots_15_io_out_uop_taken),
    .io_out_uop_imm_packed(slots_15_io_out_uop_imm_packed),
    .io_out_uop_csr_addr(slots_15_io_out_uop_csr_addr),
    .io_out_uop_rob_idx(slots_15_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx(slots_15_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx(slots_15_io_out_uop_stq_idx),
    .io_out_uop_rxq_idx(slots_15_io_out_uop_rxq_idx),
    .io_out_uop_pdst(slots_15_io_out_uop_pdst),
    .io_out_uop_prs1(slots_15_io_out_uop_prs1),
    .io_out_uop_prs2(slots_15_io_out_uop_prs2),
    .io_out_uop_prs3(slots_15_io_out_uop_prs3),
    .io_out_uop_ppred(slots_15_io_out_uop_ppred),
    .io_out_uop_prs1_busy(slots_15_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy(slots_15_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy(slots_15_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy(slots_15_io_out_uop_ppred_busy),
    .io_out_uop_stale_pdst(slots_15_io_out_uop_stale_pdst),
    .io_out_uop_exception(slots_15_io_out_uop_exception),
    .io_out_uop_exc_cause(slots_15_io_out_uop_exc_cause),
    .io_out_uop_bypassable(slots_15_io_out_uop_bypassable),
    .io_out_uop_mem_cmd(slots_15_io_out_uop_mem_cmd),
    .io_out_uop_mem_size(slots_15_io_out_uop_mem_size),
    .io_out_uop_mem_signed(slots_15_io_out_uop_mem_signed),
    .io_out_uop_is_fence(slots_15_io_out_uop_is_fence),
    .io_out_uop_is_fencei(slots_15_io_out_uop_is_fencei),
    .io_out_uop_is_amo(slots_15_io_out_uop_is_amo),
    .io_out_uop_uses_ldq(slots_15_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq(slots_15_io_out_uop_uses_stq),
    .io_out_uop_is_sys_pc2epc(slots_15_io_out_uop_is_sys_pc2epc),
    .io_out_uop_is_unique(slots_15_io_out_uop_is_unique),
    .io_out_uop_flush_on_commit(slots_15_io_out_uop_flush_on_commit),
    .io_out_uop_ldst_is_rs1(slots_15_io_out_uop_ldst_is_rs1),
    .io_out_uop_ldst(slots_15_io_out_uop_ldst),
    .io_out_uop_lrs1(slots_15_io_out_uop_lrs1),
    .io_out_uop_lrs2(slots_15_io_out_uop_lrs2),
    .io_out_uop_lrs3(slots_15_io_out_uop_lrs3),
    .io_out_uop_ldst_val(slots_15_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype(slots_15_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype(slots_15_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype(slots_15_io_out_uop_lrs2_rtype),
    .io_out_uop_frs3_en(slots_15_io_out_uop_frs3_en),
    .io_out_uop_fp_val(slots_15_io_out_uop_fp_val),
    .io_out_uop_fp_single(slots_15_io_out_uop_fp_single),
    .io_out_uop_xcpt_pf_if(slots_15_io_out_uop_xcpt_pf_if),
    .io_out_uop_xcpt_ae_if(slots_15_io_out_uop_xcpt_ae_if),
    .io_out_uop_xcpt_ma_if(slots_15_io_out_uop_xcpt_ma_if),
    .io_out_uop_bp_debug_if(slots_15_io_out_uop_bp_debug_if),
    .io_out_uop_bp_xcpt_if(slots_15_io_out_uop_bp_xcpt_if),
    .io_out_uop_debug_fsrc(slots_15_io_out_uop_debug_fsrc),
    .io_out_uop_debug_tsrc(slots_15_io_out_uop_debug_tsrc),
    .io_uop_switch(slots_15_io_uop_switch),
    .io_uop_switch_off(slots_15_io_uop_switch_off),
    .io_uop_is_unicore(slots_15_io_uop_is_unicore),
    .io_uop_shift(slots_15_io_uop_shift),
    .io_uop_lrs3_rtype(slots_15_io_uop_lrs3_rtype),
    .io_uop_rflag(slots_15_io_uop_rflag),
    .io_uop_wflag(slots_15_io_uop_wflag),
    .io_uop_prflag(slots_15_io_uop_prflag),
    .io_uop_pwflag(slots_15_io_uop_pwflag),
    .io_uop_pflag_busy(slots_15_io_uop_pflag_busy),
    .io_uop_stale_pflag(slots_15_io_uop_stale_pflag),
    .io_uop_op1_sel(slots_15_io_uop_op1_sel),
    .io_uop_op2_sel(slots_15_io_uop_op2_sel),
    .io_uop_split_num(slots_15_io_uop_split_num),
    .io_uop_self_index(slots_15_io_uop_self_index),
    .io_uop_rob_inst_idx(slots_15_io_uop_rob_inst_idx),
    .io_uop_address_num(slots_15_io_uop_address_num),
    .io_uop_uopc(slots_15_io_uop_uopc),
    .io_uop_inst(slots_15_io_uop_inst),
    .io_uop_debug_inst(slots_15_io_uop_debug_inst),
    .io_uop_is_rvc(slots_15_io_uop_is_rvc),
    .io_uop_debug_pc(slots_15_io_uop_debug_pc),
    .io_uop_iq_type(slots_15_io_uop_iq_type),
    .io_uop_fu_code(slots_15_io_uop_fu_code),
    .io_uop_ctrl_br_type(slots_15_io_uop_ctrl_br_type),
    .io_uop_ctrl_op1_sel(slots_15_io_uop_ctrl_op1_sel),
    .io_uop_ctrl_op2_sel(slots_15_io_uop_ctrl_op2_sel),
    .io_uop_ctrl_imm_sel(slots_15_io_uop_ctrl_imm_sel),
    .io_uop_ctrl_op_fcn(slots_15_io_uop_ctrl_op_fcn),
    .io_uop_ctrl_fcn_dw(slots_15_io_uop_ctrl_fcn_dw),
    .io_uop_ctrl_csr_cmd(slots_15_io_uop_ctrl_csr_cmd),
    .io_uop_ctrl_is_load(slots_15_io_uop_ctrl_is_load),
    .io_uop_ctrl_is_sta(slots_15_io_uop_ctrl_is_sta),
    .io_uop_ctrl_is_std(slots_15_io_uop_ctrl_is_std),
    .io_uop_ctrl_op3_sel(slots_15_io_uop_ctrl_op3_sel),
    .io_uop_iw_state(slots_15_io_uop_iw_state),
    .io_uop_iw_p1_poisoned(slots_15_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned(slots_15_io_uop_iw_p2_poisoned),
    .io_uop_is_br(slots_15_io_uop_is_br),
    .io_uop_is_jalr(slots_15_io_uop_is_jalr),
    .io_uop_is_jal(slots_15_io_uop_is_jal),
    .io_uop_is_sfb(slots_15_io_uop_is_sfb),
    .io_uop_br_mask(slots_15_io_uop_br_mask),
    .io_uop_br_tag(slots_15_io_uop_br_tag),
    .io_uop_ftq_idx(slots_15_io_uop_ftq_idx),
    .io_uop_edge_inst(slots_15_io_uop_edge_inst),
    .io_uop_pc_lob(slots_15_io_uop_pc_lob),
    .io_uop_taken(slots_15_io_uop_taken),
    .io_uop_imm_packed(slots_15_io_uop_imm_packed),
    .io_uop_csr_addr(slots_15_io_uop_csr_addr),
    .io_uop_rob_idx(slots_15_io_uop_rob_idx),
    .io_uop_ldq_idx(slots_15_io_uop_ldq_idx),
    .io_uop_stq_idx(slots_15_io_uop_stq_idx),
    .io_uop_rxq_idx(slots_15_io_uop_rxq_idx),
    .io_uop_pdst(slots_15_io_uop_pdst),
    .io_uop_prs1(slots_15_io_uop_prs1),
    .io_uop_prs2(slots_15_io_uop_prs2),
    .io_uop_prs3(slots_15_io_uop_prs3),
    .io_uop_ppred(slots_15_io_uop_ppred),
    .io_uop_prs1_busy(slots_15_io_uop_prs1_busy),
    .io_uop_prs2_busy(slots_15_io_uop_prs2_busy),
    .io_uop_prs3_busy(slots_15_io_uop_prs3_busy),
    .io_uop_ppred_busy(slots_15_io_uop_ppred_busy),
    .io_uop_stale_pdst(slots_15_io_uop_stale_pdst),
    .io_uop_exception(slots_15_io_uop_exception),
    .io_uop_exc_cause(slots_15_io_uop_exc_cause),
    .io_uop_bypassable(slots_15_io_uop_bypassable),
    .io_uop_mem_cmd(slots_15_io_uop_mem_cmd),
    .io_uop_mem_size(slots_15_io_uop_mem_size),
    .io_uop_mem_signed(slots_15_io_uop_mem_signed),
    .io_uop_is_fence(slots_15_io_uop_is_fence),
    .io_uop_is_fencei(slots_15_io_uop_is_fencei),
    .io_uop_is_amo(slots_15_io_uop_is_amo),
    .io_uop_uses_ldq(slots_15_io_uop_uses_ldq),
    .io_uop_uses_stq(slots_15_io_uop_uses_stq),
    .io_uop_is_sys_pc2epc(slots_15_io_uop_is_sys_pc2epc),
    .io_uop_is_unique(slots_15_io_uop_is_unique),
    .io_uop_flush_on_commit(slots_15_io_uop_flush_on_commit),
    .io_uop_ldst_is_rs1(slots_15_io_uop_ldst_is_rs1),
    .io_uop_ldst(slots_15_io_uop_ldst),
    .io_uop_lrs1(slots_15_io_uop_lrs1),
    .io_uop_lrs2(slots_15_io_uop_lrs2),
    .io_uop_lrs3(slots_15_io_uop_lrs3),
    .io_uop_ldst_val(slots_15_io_uop_ldst_val),
    .io_uop_dst_rtype(slots_15_io_uop_dst_rtype),
    .io_uop_lrs1_rtype(slots_15_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype(slots_15_io_uop_lrs2_rtype),
    .io_uop_frs3_en(slots_15_io_uop_frs3_en),
    .io_uop_fp_val(slots_15_io_uop_fp_val),
    .io_uop_fp_single(slots_15_io_uop_fp_single),
    .io_uop_xcpt_pf_if(slots_15_io_uop_xcpt_pf_if),
    .io_uop_xcpt_ae_if(slots_15_io_uop_xcpt_ae_if),
    .io_uop_xcpt_ma_if(slots_15_io_uop_xcpt_ma_if),
    .io_uop_bp_debug_if(slots_15_io_uop_bp_debug_if),
    .io_uop_bp_xcpt_if(slots_15_io_uop_bp_xcpt_if),
    .io_uop_debug_fsrc(slots_15_io_uop_debug_fsrc),
    .io_uop_debug_tsrc(slots_15_io_uop_debug_tsrc),
    .io_debug_p1(slots_15_io_debug_p1),
    .io_debug_p2(slots_15_io_debug_p2),
    .io_debug_p3(slots_15_io_debug_p3),
    .io_debug_ppred(slots_15_io_debug_ppred),
    .io_debug_state(slots_15_io_debug_state)
  );
  assign io_dis_uops_0_ready = REG; // @[issue-unit-age-ordered.scala 87:26]
  assign io_dis_uops_1_ready = REG_1; // @[issue-unit-age-ordered.scala 87:26]
  assign io_iss_valids_0 = issue_slots_15_grant | (issue_slots_14_grant | (issue_slots_13_grant | (issue_slots_12_grant
     | (issue_slots_11_grant | (issue_slots_10_grant | (issue_slots_9_grant | (issue_slots_8_grant | (
    issue_slots_7_grant | (issue_slots_6_grant | (issue_slots_5_grant | (issue_slots_4_grant | (issue_slots_3_grant | (
    issue_slots_2_grant | (issue_slots_1_grant | issue_slots_0_grant)))))))))))))); // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 124:26]
  assign io_iss_uops_0_switch = issue_slots_15_grant ? issue_slots_15_uop_switch : _GEN_4657; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_switch_off = issue_slots_15_grant ? issue_slots_15_uop_switch_off : _GEN_4656; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_unicore = issue_slots_15_grant ? issue_slots_15_uop_is_unicore : _GEN_4655; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_shift = issue_slots_15_grant ? issue_slots_15_uop_shift : _GEN_4654; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_lrs3_rtype = issue_slots_15_grant ? issue_slots_15_uop_lrs3_rtype : _GEN_4653; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_rflag = issue_slots_15_grant ? issue_slots_15_uop_rflag : _GEN_4652; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_wflag = issue_slots_15_grant ? issue_slots_15_uop_wflag : _GEN_4651; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_prflag = issue_slots_15_grant ? issue_slots_15_uop_prflag : _GEN_4650; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_pwflag = issue_slots_15_grant ? issue_slots_15_uop_pwflag : _GEN_4649; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_pflag_busy = issue_slots_15_grant ? issue_slots_15_uop_pflag_busy : _GEN_4648; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_stale_pflag = issue_slots_15_grant ? issue_slots_15_uop_stale_pflag : _GEN_4647; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_op1_sel = issue_slots_15_grant ? issue_slots_15_uop_op1_sel : _GEN_4646; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_op2_sel = issue_slots_15_grant ? issue_slots_15_uop_op2_sel : _GEN_4645; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_split_num = issue_slots_15_grant ? issue_slots_15_uop_split_num : _GEN_4644; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_self_index = issue_slots_15_grant ? issue_slots_15_uop_self_index : _GEN_4643; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_rob_inst_idx = issue_slots_15_grant ? issue_slots_15_uop_rob_inst_idx : _GEN_4642; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_address_num = issue_slots_15_grant ? issue_slots_15_uop_address_num : _GEN_4641; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_uopc = issue_slots_15_grant ? issue_slots_15_uop_uopc : _GEN_4640; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_inst = issue_slots_15_grant ? issue_slots_15_uop_inst : _GEN_4639; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_debug_inst = issue_slots_15_grant ? issue_slots_15_uop_debug_inst : _GEN_4638; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_rvc = issue_slots_15_grant ? issue_slots_15_uop_is_rvc : _GEN_4637; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_debug_pc = issue_slots_15_grant ? issue_slots_15_uop_debug_pc : _GEN_4636; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_iq_type = issue_slots_15_grant ? issue_slots_15_uop_iq_type : _GEN_4635; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_fu_code = issue_slots_15_grant ? issue_slots_15_uop_fu_code : _GEN_4634; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_br_type = issue_slots_15_grant ? issue_slots_15_uop_ctrl_br_type : _GEN_4633; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_op1_sel = issue_slots_15_grant ? issue_slots_15_uop_ctrl_op1_sel : _GEN_4632; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_op2_sel = issue_slots_15_grant ? issue_slots_15_uop_ctrl_op2_sel : _GEN_4631; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_imm_sel = issue_slots_15_grant ? issue_slots_15_uop_ctrl_imm_sel : _GEN_4630; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_op_fcn = issue_slots_15_grant ? issue_slots_15_uop_ctrl_op_fcn : _GEN_4629; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_fcn_dw = issue_slots_15_grant ? issue_slots_15_uop_ctrl_fcn_dw : _GEN_4628; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_csr_cmd = issue_slots_15_grant ? issue_slots_15_uop_ctrl_csr_cmd : _GEN_4627; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_is_load = issue_slots_15_grant ? issue_slots_15_uop_ctrl_is_load : _GEN_4626; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_is_sta = issue_slots_15_grant ? issue_slots_15_uop_ctrl_is_sta : _GEN_4625; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_is_std = issue_slots_15_grant ? issue_slots_15_uop_ctrl_is_std : _GEN_4624; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ctrl_op3_sel = issue_slots_15_grant ? issue_slots_15_uop_ctrl_op3_sel : _GEN_4623; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_iw_state = issue_slots_15_grant ? issue_slots_15_uop_iw_state : _GEN_4622; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_iw_p1_poisoned = issue_slots_15_grant ? issue_slots_15_uop_iw_p1_poisoned : _GEN_4621; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_iw_p2_poisoned = issue_slots_15_grant ? issue_slots_15_uop_iw_p2_poisoned : _GEN_4620; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_br = issue_slots_15_grant ? issue_slots_15_uop_is_br : _GEN_4619; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_jalr = issue_slots_15_grant ? issue_slots_15_uop_is_jalr : _GEN_4618; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_jal = issue_slots_15_grant ? issue_slots_15_uop_is_jal : _GEN_4617; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_sfb = issue_slots_15_grant ? issue_slots_15_uop_is_sfb : _GEN_4616; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_br_mask = issue_slots_15_grant ? issue_slots_15_uop_br_mask : _GEN_4615; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_br_tag = issue_slots_15_grant ? issue_slots_15_uop_br_tag : _GEN_4614; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ftq_idx = issue_slots_15_grant ? issue_slots_15_uop_ftq_idx : _GEN_4613; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_edge_inst = issue_slots_15_grant ? issue_slots_15_uop_edge_inst : _GEN_4612; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_pc_lob = issue_slots_15_grant ? issue_slots_15_uop_pc_lob : _GEN_4611; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_taken = issue_slots_15_grant ? issue_slots_15_uop_taken : _GEN_4610; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_imm_packed = issue_slots_15_grant ? issue_slots_15_uop_imm_packed : _GEN_4609; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_csr_addr = issue_slots_15_grant ? issue_slots_15_uop_csr_addr : _GEN_4608; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_rob_idx = issue_slots_15_grant ? issue_slots_15_uop_rob_idx : _GEN_4607; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ldq_idx = issue_slots_15_grant ? issue_slots_15_uop_ldq_idx : _GEN_4606; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_stq_idx = issue_slots_15_grant ? issue_slots_15_uop_stq_idx : _GEN_4605; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_rxq_idx = issue_slots_15_grant ? issue_slots_15_uop_rxq_idx : _GEN_4604; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_pdst = issue_slots_15_grant ? issue_slots_15_uop_pdst : _GEN_4603; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_prs1 = issue_slots_15_grant ? issue_slots_15_uop_prs1 : _GEN_4602; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_prs2 = issue_slots_15_grant ? issue_slots_15_uop_prs2 : _GEN_4601; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_prs3 = issue_slots_15_grant ? issue_slots_15_uop_prs3 : _GEN_4600; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ppred = issue_slots_15_grant ? issue_slots_15_uop_ppred : _GEN_4599; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_prs1_busy = issue_slots_15_grant ? issue_slots_15_uop_prs1_busy : _GEN_4598; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_prs2_busy = issue_slots_15_grant ? issue_slots_15_uop_prs2_busy : _GEN_4597; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_prs3_busy = issue_slots_15_grant ? issue_slots_15_uop_prs3_busy : _GEN_4596; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ppred_busy = issue_slots_15_grant ? issue_slots_15_uop_ppred_busy : _GEN_4595; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_stale_pdst = issue_slots_15_grant ? issue_slots_15_uop_stale_pdst : _GEN_4594; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_exception = issue_slots_15_grant ? issue_slots_15_uop_exception : _GEN_4593; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_exc_cause = issue_slots_15_grant ? issue_slots_15_uop_exc_cause : _GEN_4592; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_bypassable = issue_slots_15_grant ? issue_slots_15_uop_bypassable : _GEN_4591; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_mem_cmd = issue_slots_15_grant ? issue_slots_15_uop_mem_cmd : _GEN_4590; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_mem_size = issue_slots_15_grant ? issue_slots_15_uop_mem_size : _GEN_4589; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_mem_signed = issue_slots_15_grant ? issue_slots_15_uop_mem_signed : _GEN_4588; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_fence = issue_slots_15_grant ? issue_slots_15_uop_is_fence : _GEN_4587; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_fencei = issue_slots_15_grant ? issue_slots_15_uop_is_fencei : _GEN_4586; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_amo = issue_slots_15_grant ? issue_slots_15_uop_is_amo : _GEN_4585; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_uses_ldq = issue_slots_15_grant ? issue_slots_15_uop_uses_ldq : _GEN_4584; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_uses_stq = issue_slots_15_grant ? issue_slots_15_uop_uses_stq : _GEN_4583; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_sys_pc2epc = issue_slots_15_grant ? issue_slots_15_uop_is_sys_pc2epc : _GEN_4582; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_is_unique = issue_slots_15_grant ? issue_slots_15_uop_is_unique : _GEN_4581; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_flush_on_commit = issue_slots_15_grant ? issue_slots_15_uop_flush_on_commit : _GEN_4580; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ldst_is_rs1 = issue_slots_15_grant ? issue_slots_15_uop_ldst_is_rs1 : _GEN_4579; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ldst = issue_slots_15_grant ? issue_slots_15_uop_ldst : _GEN_4578; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_lrs1 = issue_slots_15_grant ? issue_slots_15_uop_lrs1 : _GEN_4577; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_lrs2 = issue_slots_15_grant ? issue_slots_15_uop_lrs2 : _GEN_4576; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_lrs3 = issue_slots_15_grant ? issue_slots_15_uop_lrs3 : _GEN_4575; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_ldst_val = issue_slots_15_grant ? issue_slots_15_uop_ldst_val : _GEN_4574; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_dst_rtype = issue_slots_15_grant ? issue_slots_15_uop_dst_rtype : _GEN_4573; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_lrs1_rtype = issue_slots_15_grant ? issue_slots_15_uop_lrs1_rtype : _GEN_4572; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_lrs2_rtype = issue_slots_15_grant ? issue_slots_15_uop_lrs2_rtype : _GEN_4571; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_frs3_en = issue_slots_15_grant ? issue_slots_15_uop_frs3_en : _GEN_4570; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_fp_val = issue_slots_15_grant ? issue_slots_15_uop_fp_val : _GEN_4569; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_fp_single = issue_slots_15_grant ? issue_slots_15_uop_fp_single : _GEN_4568; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_xcpt_pf_if = issue_slots_15_grant ? issue_slots_15_uop_xcpt_pf_if : _GEN_4567; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_xcpt_ae_if = issue_slots_15_grant ? issue_slots_15_uop_xcpt_ae_if : _GEN_4566; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_xcpt_ma_if = issue_slots_15_grant ? issue_slots_15_uop_xcpt_ma_if : _GEN_4565; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_bp_debug_if = issue_slots_15_grant ? issue_slots_15_uop_bp_debug_if : _GEN_4564; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_bp_xcpt_if = issue_slots_15_grant ? issue_slots_15_uop_bp_xcpt_if : _GEN_4563; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_debug_fsrc = issue_slots_15_grant ? issue_slots_15_uop_debug_fsrc : _GEN_4562; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_iss_uops_0_debug_tsrc = issue_slots_15_grant ? issue_slots_15_uop_debug_tsrc : _GEN_4561; // @[issue-unit-age-ordered.scala 122:76 issue-unit-age-ordered.scala 125:24]
  assign io_event_empty = ~(issue_slots_0_valid | issue_slots_1_valid | issue_slots_2_valid | issue_slots_3_valid |
    issue_slots_4_valid | issue_slots_5_valid | issue_slots_6_valid | issue_slots_7_valid | issue_slots_8_valid |
    issue_slots_9_valid | issue_slots_10_valid | issue_slots_11_valid | issue_slots_12_valid | issue_slots_13_valid |
    issue_slots_14_valid | issue_slots_15_valid); // @[issue-unit.scala 169:21]
  assign slots_0_clock = clock;
  assign slots_0_reset = reset;
  assign slots_0_io_grant = issue_slots_0_request & _T_333; // @[issue-unit-age-ordered.scala 122:40]
  assign slots_0_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_0_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_0_io_clear = 1'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_0_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_0_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_0_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_0_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_0_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_0_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_0_io_in_uop_valid = _GEN_7[1:0] == 2'h2 ? issue_slots_2_will_be_valid : _GEN_38; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_0_io_in_uop_bits_switch = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_switch :
    issue_slots_1_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_switch_off = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_switch_off :
    issue_slots_1_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_unicore = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_is_unicore :
    issue_slots_1_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_shift = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_shift : issue_slots_1_out_uop_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_lrs3_rtype = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_lrs3_rtype :
    issue_slots_1_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_rflag = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_rflag : issue_slots_1_out_uop_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_wflag = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_wflag : issue_slots_1_out_uop_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_prflag = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_prflag :
    issue_slots_1_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_pwflag = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_pwflag :
    issue_slots_1_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_pflag_busy = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_pflag_busy :
    issue_slots_1_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_stale_pflag = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_stale_pflag :
    issue_slots_1_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_op1_sel = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_op1_sel :
    issue_slots_1_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_op2_sel = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_op2_sel :
    issue_slots_1_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_split_num = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_split_num :
    issue_slots_1_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_self_index = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_self_index :
    issue_slots_1_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_rob_inst_idx = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_rob_inst_idx :
    issue_slots_1_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_address_num = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_address_num :
    issue_slots_1_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_uopc = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_uopc : issue_slots_1_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_inst = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_inst : issue_slots_1_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_debug_inst = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_debug_inst :
    issue_slots_1_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_rvc = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_is_rvc :
    issue_slots_1_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_debug_pc = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_debug_pc :
    issue_slots_1_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_iq_type = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_iq_type :
    issue_slots_1_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_fu_code = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_fu_code :
    issue_slots_1_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_br_type = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_br_type :
    issue_slots_1_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_op1_sel = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_op1_sel :
    issue_slots_1_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_op2_sel = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_op2_sel :
    issue_slots_1_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_imm_sel = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_imm_sel :
    issue_slots_1_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_op_fcn = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_op_fcn :
    issue_slots_1_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_fcn_dw = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_fcn_dw :
    issue_slots_1_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_csr_cmd = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_csr_cmd :
    issue_slots_1_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_is_load = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_is_load :
    issue_slots_1_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_is_sta = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_is_sta :
    issue_slots_1_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_is_std = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_is_std :
    issue_slots_1_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ctrl_op3_sel = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_ctrl_op3_sel :
    issue_slots_1_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_iw_state = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_iw_state :
    issue_slots_1_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_iw_p1_poisoned = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_iw_p1_poisoned :
    issue_slots_1_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_iw_p2_poisoned = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_iw_p2_poisoned :
    issue_slots_1_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_br = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_is_br : issue_slots_1_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_jalr = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_is_jalr :
    issue_slots_1_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_jal = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_is_jal :
    issue_slots_1_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_sfb = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_is_sfb :
    issue_slots_1_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_br_mask = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_br_mask :
    issue_slots_1_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_br_tag = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_br_tag :
    issue_slots_1_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ftq_idx = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_ftq_idx :
    issue_slots_1_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_edge_inst = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_edge_inst :
    issue_slots_1_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_pc_lob = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_pc_lob :
    issue_slots_1_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_taken = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_taken : issue_slots_1_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_imm_packed = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_imm_packed :
    issue_slots_1_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_csr_addr = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_csr_addr :
    issue_slots_1_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_rob_idx = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_rob_idx :
    issue_slots_1_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ldq_idx = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_ldq_idx :
    issue_slots_1_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_stq_idx = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_stq_idx :
    issue_slots_1_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_rxq_idx = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_rxq_idx :
    issue_slots_1_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_pdst = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_pdst : issue_slots_1_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_prs1 = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_prs1 : issue_slots_1_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_prs2 = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_prs2 : issue_slots_1_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_prs3 = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_prs3 : issue_slots_1_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ppred = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_ppred : issue_slots_1_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_prs1_busy = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_prs1_busy :
    issue_slots_1_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_prs2_busy = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_prs2_busy :
    issue_slots_1_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_prs3_busy = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_prs3_busy :
    issue_slots_1_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ppred_busy = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_ppred_busy :
    issue_slots_1_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_stale_pdst = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_stale_pdst :
    issue_slots_1_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_exception = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_exception :
    issue_slots_1_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_exc_cause = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_exc_cause :
    issue_slots_1_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_bypassable = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_bypassable :
    issue_slots_1_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_mem_cmd = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_mem_cmd :
    issue_slots_1_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_mem_size = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_mem_size :
    issue_slots_1_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_mem_signed = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_mem_signed :
    issue_slots_1_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_fence = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_is_fence :
    issue_slots_1_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_fencei = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_is_fencei :
    issue_slots_1_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_amo = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_is_amo :
    issue_slots_1_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_uses_ldq = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_uses_ldq :
    issue_slots_1_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_uses_stq = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_uses_stq :
    issue_slots_1_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_sys_pc2epc = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_is_sys_pc2epc :
    issue_slots_1_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_is_unique = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_is_unique :
    issue_slots_1_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_flush_on_commit = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_flush_on_commit :
    issue_slots_1_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ldst_is_rs1 = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_ldst_is_rs1 :
    issue_slots_1_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ldst = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_ldst : issue_slots_1_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_lrs1 = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_lrs1 : issue_slots_1_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_lrs2 = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_lrs2 : issue_slots_1_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_lrs3 = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_lrs3 : issue_slots_1_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_ldst_val = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_ldst_val :
    issue_slots_1_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_dst_rtype = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_dst_rtype :
    issue_slots_1_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_lrs1_rtype = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_lrs1_rtype :
    issue_slots_1_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_lrs2_rtype = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_lrs2_rtype :
    issue_slots_1_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_frs3_en = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_frs3_en :
    issue_slots_1_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_fp_val = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_fp_val :
    issue_slots_1_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_fp_single = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_fp_single :
    issue_slots_1_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_xcpt_pf_if = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_xcpt_pf_if :
    issue_slots_1_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_xcpt_ae_if = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_xcpt_ae_if :
    issue_slots_1_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_xcpt_ma_if = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_xcpt_ma_if :
    issue_slots_1_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_bp_debug_if = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_bp_debug_if :
    issue_slots_1_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_bp_xcpt_if = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_bp_xcpt_if :
    issue_slots_1_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_debug_fsrc = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_debug_fsrc :
    issue_slots_1_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_0_io_in_uop_bits_debug_tsrc = _GEN_7[1:0] == 2'h2 ? issue_slots_2_out_uop_debug_tsrc :
    issue_slots_1_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_clock = clock;
  assign slots_1_reset = reset;
  assign slots_1_io_grant = issue_slots_1_request & _T_348 & ~issue_slots_0_grant; // @[issue-unit-age-ordered.scala 122:56]
  assign slots_1_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_1_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_1_io_clear = _GEN_5[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_1_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_1_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_1_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_1_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_1_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_1_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_1_io_in_uop_valid = _GEN_9[1:0] == 2'h2 ? issue_slots_3_will_be_valid : _GEN_234; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_1_io_in_uop_bits_switch = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_switch :
    issue_slots_2_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_switch_off = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_switch_off :
    issue_slots_2_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_unicore = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_is_unicore :
    issue_slots_2_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_shift = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_shift : issue_slots_2_out_uop_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_lrs3_rtype = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_lrs3_rtype :
    issue_slots_2_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_rflag = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_rflag : issue_slots_2_out_uop_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_wflag = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_wflag : issue_slots_2_out_uop_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_prflag = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_prflag :
    issue_slots_2_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_pwflag = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_pwflag :
    issue_slots_2_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_pflag_busy = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_pflag_busy :
    issue_slots_2_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_stale_pflag = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_stale_pflag :
    issue_slots_2_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_op1_sel = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_op1_sel :
    issue_slots_2_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_op2_sel = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_op2_sel :
    issue_slots_2_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_split_num = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_split_num :
    issue_slots_2_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_self_index = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_self_index :
    issue_slots_2_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_rob_inst_idx = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_rob_inst_idx :
    issue_slots_2_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_address_num = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_address_num :
    issue_slots_2_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_uopc = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_uopc : issue_slots_2_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_inst = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_inst : issue_slots_2_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_debug_inst = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_debug_inst :
    issue_slots_2_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_rvc = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_is_rvc :
    issue_slots_2_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_debug_pc = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_debug_pc :
    issue_slots_2_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_iq_type = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_iq_type :
    issue_slots_2_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_fu_code = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_fu_code :
    issue_slots_2_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_br_type = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_br_type :
    issue_slots_2_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_op1_sel = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_op1_sel :
    issue_slots_2_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_op2_sel = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_op2_sel :
    issue_slots_2_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_imm_sel = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_imm_sel :
    issue_slots_2_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_op_fcn = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_op_fcn :
    issue_slots_2_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_fcn_dw = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_fcn_dw :
    issue_slots_2_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_csr_cmd = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_csr_cmd :
    issue_slots_2_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_is_load = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_is_load :
    issue_slots_2_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_is_sta = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_is_sta :
    issue_slots_2_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_is_std = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_is_std :
    issue_slots_2_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ctrl_op3_sel = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_ctrl_op3_sel :
    issue_slots_2_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_iw_state = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_iw_state :
    issue_slots_2_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_iw_p1_poisoned = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_iw_p1_poisoned :
    issue_slots_2_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_iw_p2_poisoned = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_iw_p2_poisoned :
    issue_slots_2_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_br = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_is_br : issue_slots_2_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_jalr = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_is_jalr :
    issue_slots_2_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_jal = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_is_jal :
    issue_slots_2_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_sfb = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_is_sfb :
    issue_slots_2_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_br_mask = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_br_mask :
    issue_slots_2_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_br_tag = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_br_tag :
    issue_slots_2_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ftq_idx = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_ftq_idx :
    issue_slots_2_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_edge_inst = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_edge_inst :
    issue_slots_2_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_pc_lob = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_pc_lob :
    issue_slots_2_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_taken = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_taken : issue_slots_2_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_imm_packed = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_imm_packed :
    issue_slots_2_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_csr_addr = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_csr_addr :
    issue_slots_2_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_rob_idx = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_rob_idx :
    issue_slots_2_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ldq_idx = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_ldq_idx :
    issue_slots_2_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_stq_idx = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_stq_idx :
    issue_slots_2_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_rxq_idx = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_rxq_idx :
    issue_slots_2_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_pdst = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_pdst : issue_slots_2_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_prs1 = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_prs1 : issue_slots_2_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_prs2 = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_prs2 : issue_slots_2_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_prs3 = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_prs3 : issue_slots_2_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ppred = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_ppred : issue_slots_2_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_prs1_busy = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_prs1_busy :
    issue_slots_2_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_prs2_busy = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_prs2_busy :
    issue_slots_2_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_prs3_busy = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_prs3_busy :
    issue_slots_2_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ppred_busy = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_ppred_busy :
    issue_slots_2_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_stale_pdst = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_stale_pdst :
    issue_slots_2_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_exception = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_exception :
    issue_slots_2_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_exc_cause = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_exc_cause :
    issue_slots_2_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_bypassable = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_bypassable :
    issue_slots_2_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_mem_cmd = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_mem_cmd :
    issue_slots_2_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_mem_size = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_mem_size :
    issue_slots_2_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_mem_signed = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_mem_signed :
    issue_slots_2_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_fence = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_is_fence :
    issue_slots_2_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_fencei = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_is_fencei :
    issue_slots_2_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_amo = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_is_amo :
    issue_slots_2_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_uses_ldq = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_uses_ldq :
    issue_slots_2_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_uses_stq = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_uses_stq :
    issue_slots_2_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_sys_pc2epc = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_is_sys_pc2epc :
    issue_slots_2_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_is_unique = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_is_unique :
    issue_slots_2_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_flush_on_commit = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_flush_on_commit :
    issue_slots_2_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ldst_is_rs1 = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_ldst_is_rs1 :
    issue_slots_2_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ldst = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_ldst : issue_slots_2_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_lrs1 = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_lrs1 : issue_slots_2_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_lrs2 = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_lrs2 : issue_slots_2_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_lrs3 = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_lrs3 : issue_slots_2_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_ldst_val = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_ldst_val :
    issue_slots_2_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_dst_rtype = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_dst_rtype :
    issue_slots_2_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_lrs1_rtype = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_lrs1_rtype :
    issue_slots_2_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_lrs2_rtype = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_lrs2_rtype :
    issue_slots_2_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_frs3_en = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_frs3_en :
    issue_slots_2_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_fp_val = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_fp_val :
    issue_slots_2_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_fp_single = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_fp_single :
    issue_slots_2_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_xcpt_pf_if = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_xcpt_pf_if :
    issue_slots_2_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_xcpt_ae_if = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_xcpt_ae_if :
    issue_slots_2_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_xcpt_ma_if = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_xcpt_ma_if :
    issue_slots_2_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_bp_debug_if = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_bp_debug_if :
    issue_slots_2_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_bp_xcpt_if = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_bp_xcpt_if :
    issue_slots_2_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_debug_fsrc = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_debug_fsrc :
    issue_slots_2_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_1_io_in_uop_bits_debug_tsrc = _GEN_9[1:0] == 2'h2 ? issue_slots_3_out_uop_debug_tsrc :
    issue_slots_2_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_clock = clock;
  assign slots_2_reset = reset;
  assign slots_2_io_grant = issue_slots_2_request & _T_363 & ~_T_357; // @[issue-unit-age-ordered.scala 122:56]
  assign slots_2_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_2_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_2_io_clear = _GEN_7[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_2_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_2_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_2_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_2_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_2_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_2_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_2_io_in_uop_valid = _GEN_11[1:0] == 2'h2 ? issue_slots_4_will_be_valid : _GEN_430; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_2_io_in_uop_bits_switch = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_switch :
    issue_slots_3_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_switch_off = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_switch_off :
    issue_slots_3_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_unicore = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_is_unicore :
    issue_slots_3_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_shift = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_shift : issue_slots_3_out_uop_shift
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_lrs3_rtype = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_lrs3_rtype :
    issue_slots_3_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_rflag = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_rflag : issue_slots_3_out_uop_rflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_wflag = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_wflag : issue_slots_3_out_uop_wflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_prflag = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_prflag :
    issue_slots_3_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_pwflag = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_pwflag :
    issue_slots_3_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_pflag_busy = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_pflag_busy :
    issue_slots_3_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_stale_pflag = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_stale_pflag :
    issue_slots_3_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_op1_sel = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_op1_sel :
    issue_slots_3_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_op2_sel = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_op2_sel :
    issue_slots_3_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_split_num = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_split_num :
    issue_slots_3_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_self_index = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_self_index :
    issue_slots_3_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_rob_inst_idx = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_rob_inst_idx :
    issue_slots_3_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_address_num = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_address_num :
    issue_slots_3_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_uopc = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_uopc : issue_slots_3_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_inst = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_inst : issue_slots_3_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_debug_inst = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_debug_inst :
    issue_slots_3_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_rvc = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_is_rvc :
    issue_slots_3_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_debug_pc = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_debug_pc :
    issue_slots_3_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_iq_type = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_iq_type :
    issue_slots_3_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_fu_code = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_fu_code :
    issue_slots_3_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_br_type = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_br_type :
    issue_slots_3_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_op1_sel = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_op1_sel :
    issue_slots_3_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_op2_sel = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_op2_sel :
    issue_slots_3_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_imm_sel = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_imm_sel :
    issue_slots_3_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_op_fcn = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_op_fcn :
    issue_slots_3_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_fcn_dw = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_fcn_dw :
    issue_slots_3_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_csr_cmd = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_csr_cmd :
    issue_slots_3_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_is_load = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_is_load :
    issue_slots_3_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_is_sta = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_is_sta :
    issue_slots_3_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_is_std = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_is_std :
    issue_slots_3_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ctrl_op3_sel = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_ctrl_op3_sel :
    issue_slots_3_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_iw_state = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_iw_state :
    issue_slots_3_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_iw_p1_poisoned = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_iw_p1_poisoned :
    issue_slots_3_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_iw_p2_poisoned = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_iw_p2_poisoned :
    issue_slots_3_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_br = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_is_br : issue_slots_3_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_jalr = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_is_jalr :
    issue_slots_3_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_jal = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_is_jal :
    issue_slots_3_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_sfb = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_is_sfb :
    issue_slots_3_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_br_mask = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_br_mask :
    issue_slots_3_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_br_tag = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_br_tag :
    issue_slots_3_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ftq_idx = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_ftq_idx :
    issue_slots_3_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_edge_inst = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_edge_inst :
    issue_slots_3_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_pc_lob = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_pc_lob :
    issue_slots_3_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_taken = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_taken : issue_slots_3_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_imm_packed = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_imm_packed :
    issue_slots_3_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_csr_addr = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_csr_addr :
    issue_slots_3_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_rob_idx = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_rob_idx :
    issue_slots_3_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ldq_idx = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_ldq_idx :
    issue_slots_3_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_stq_idx = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_stq_idx :
    issue_slots_3_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_rxq_idx = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_rxq_idx :
    issue_slots_3_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_pdst = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_pdst : issue_slots_3_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_prs1 = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_prs1 : issue_slots_3_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_prs2 = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_prs2 : issue_slots_3_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_prs3 = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_prs3 : issue_slots_3_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ppred = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_ppred : issue_slots_3_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_prs1_busy = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_prs1_busy :
    issue_slots_3_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_prs2_busy = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_prs2_busy :
    issue_slots_3_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_prs3_busy = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_prs3_busy :
    issue_slots_3_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ppred_busy = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_ppred_busy :
    issue_slots_3_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_stale_pdst = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_stale_pdst :
    issue_slots_3_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_exception = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_exception :
    issue_slots_3_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_exc_cause = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_exc_cause :
    issue_slots_3_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_bypassable = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_bypassable :
    issue_slots_3_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_mem_cmd = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_mem_cmd :
    issue_slots_3_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_mem_size = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_mem_size :
    issue_slots_3_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_mem_signed = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_mem_signed :
    issue_slots_3_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_fence = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_is_fence :
    issue_slots_3_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_fencei = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_is_fencei :
    issue_slots_3_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_amo = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_is_amo :
    issue_slots_3_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_uses_ldq = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_uses_ldq :
    issue_slots_3_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_uses_stq = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_uses_stq :
    issue_slots_3_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_sys_pc2epc = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_is_sys_pc2epc :
    issue_slots_3_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_is_unique = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_is_unique :
    issue_slots_3_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_flush_on_commit = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_flush_on_commit :
    issue_slots_3_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ldst_is_rs1 = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_ldst_is_rs1 :
    issue_slots_3_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ldst = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_ldst : issue_slots_3_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_lrs1 = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_lrs1 : issue_slots_3_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_lrs2 = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_lrs2 : issue_slots_3_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_lrs3 = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_lrs3 : issue_slots_3_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_ldst_val = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_ldst_val :
    issue_slots_3_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_dst_rtype = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_dst_rtype :
    issue_slots_3_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_lrs1_rtype = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_lrs1_rtype :
    issue_slots_3_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_lrs2_rtype = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_lrs2_rtype :
    issue_slots_3_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_frs3_en = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_frs3_en :
    issue_slots_3_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_fp_val = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_fp_val :
    issue_slots_3_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_fp_single = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_fp_single :
    issue_slots_3_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_xcpt_pf_if = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_xcpt_pf_if :
    issue_slots_3_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_xcpt_ae_if = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_xcpt_ae_if :
    issue_slots_3_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_xcpt_ma_if = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_xcpt_ma_if :
    issue_slots_3_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_bp_debug_if = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_bp_debug_if :
    issue_slots_3_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_bp_xcpt_if = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_bp_xcpt_if :
    issue_slots_3_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_debug_fsrc = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_debug_fsrc :
    issue_slots_3_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_2_io_in_uop_bits_debug_tsrc = _GEN_11[1:0] == 2'h2 ? issue_slots_4_out_uop_debug_tsrc :
    issue_slots_3_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_clock = clock;
  assign slots_3_reset = reset;
  assign slots_3_io_grant = issue_slots_3_request & _T_378 & ~_T_372; // @[issue-unit-age-ordered.scala 122:56]
  assign slots_3_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_3_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_3_io_clear = _GEN_9[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_3_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_3_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_3_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_3_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_3_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_3_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_3_io_in_uop_valid = _GEN_13[1:0] == 2'h2 ? issue_slots_5_will_be_valid : _GEN_626; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_3_io_in_uop_bits_switch = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_switch :
    issue_slots_4_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_switch_off = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_switch_off :
    issue_slots_4_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_unicore = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_is_unicore :
    issue_slots_4_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_shift = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_shift : issue_slots_4_out_uop_shift
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_lrs3_rtype = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_lrs3_rtype :
    issue_slots_4_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_rflag = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_rflag : issue_slots_4_out_uop_rflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_wflag = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_wflag : issue_slots_4_out_uop_wflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_prflag = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_prflag :
    issue_slots_4_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_pwflag = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_pwflag :
    issue_slots_4_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_pflag_busy = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_pflag_busy :
    issue_slots_4_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_stale_pflag = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_stale_pflag :
    issue_slots_4_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_op1_sel = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_op1_sel :
    issue_slots_4_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_op2_sel = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_op2_sel :
    issue_slots_4_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_split_num = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_split_num :
    issue_slots_4_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_self_index = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_self_index :
    issue_slots_4_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_rob_inst_idx = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_rob_inst_idx :
    issue_slots_4_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_address_num = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_address_num :
    issue_slots_4_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_uopc = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_uopc : issue_slots_4_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_inst = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_inst : issue_slots_4_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_debug_inst = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_debug_inst :
    issue_slots_4_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_rvc = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_is_rvc :
    issue_slots_4_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_debug_pc = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_debug_pc :
    issue_slots_4_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_iq_type = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_iq_type :
    issue_slots_4_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_fu_code = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_fu_code :
    issue_slots_4_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_br_type = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_br_type :
    issue_slots_4_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_op1_sel = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_op1_sel :
    issue_slots_4_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_op2_sel = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_op2_sel :
    issue_slots_4_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_imm_sel = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_imm_sel :
    issue_slots_4_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_op_fcn = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_op_fcn :
    issue_slots_4_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_fcn_dw = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_fcn_dw :
    issue_slots_4_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_csr_cmd = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_csr_cmd :
    issue_slots_4_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_is_load = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_is_load :
    issue_slots_4_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_is_sta = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_is_sta :
    issue_slots_4_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_is_std = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_is_std :
    issue_slots_4_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ctrl_op3_sel = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_ctrl_op3_sel :
    issue_slots_4_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_iw_state = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_iw_state :
    issue_slots_4_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_iw_p1_poisoned = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_iw_p1_poisoned :
    issue_slots_4_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_iw_p2_poisoned = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_iw_p2_poisoned :
    issue_slots_4_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_br = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_is_br : issue_slots_4_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_jalr = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_is_jalr :
    issue_slots_4_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_jal = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_is_jal :
    issue_slots_4_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_sfb = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_is_sfb :
    issue_slots_4_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_br_mask = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_br_mask :
    issue_slots_4_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_br_tag = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_br_tag :
    issue_slots_4_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ftq_idx = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_ftq_idx :
    issue_slots_4_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_edge_inst = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_edge_inst :
    issue_slots_4_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_pc_lob = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_pc_lob :
    issue_slots_4_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_taken = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_taken : issue_slots_4_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_imm_packed = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_imm_packed :
    issue_slots_4_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_csr_addr = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_csr_addr :
    issue_slots_4_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_rob_idx = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_rob_idx :
    issue_slots_4_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ldq_idx = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_ldq_idx :
    issue_slots_4_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_stq_idx = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_stq_idx :
    issue_slots_4_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_rxq_idx = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_rxq_idx :
    issue_slots_4_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_pdst = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_pdst : issue_slots_4_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_prs1 = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_prs1 : issue_slots_4_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_prs2 = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_prs2 : issue_slots_4_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_prs3 = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_prs3 : issue_slots_4_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ppred = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_ppred : issue_slots_4_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_prs1_busy = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_prs1_busy :
    issue_slots_4_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_prs2_busy = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_prs2_busy :
    issue_slots_4_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_prs3_busy = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_prs3_busy :
    issue_slots_4_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ppred_busy = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_ppred_busy :
    issue_slots_4_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_stale_pdst = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_stale_pdst :
    issue_slots_4_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_exception = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_exception :
    issue_slots_4_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_exc_cause = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_exc_cause :
    issue_slots_4_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_bypassable = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_bypassable :
    issue_slots_4_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_mem_cmd = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_mem_cmd :
    issue_slots_4_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_mem_size = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_mem_size :
    issue_slots_4_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_mem_signed = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_mem_signed :
    issue_slots_4_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_fence = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_is_fence :
    issue_slots_4_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_fencei = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_is_fencei :
    issue_slots_4_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_amo = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_is_amo :
    issue_slots_4_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_uses_ldq = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_uses_ldq :
    issue_slots_4_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_uses_stq = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_uses_stq :
    issue_slots_4_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_sys_pc2epc = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_is_sys_pc2epc :
    issue_slots_4_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_is_unique = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_is_unique :
    issue_slots_4_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_flush_on_commit = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_flush_on_commit :
    issue_slots_4_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ldst_is_rs1 = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_ldst_is_rs1 :
    issue_slots_4_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ldst = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_ldst : issue_slots_4_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_lrs1 = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_lrs1 : issue_slots_4_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_lrs2 = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_lrs2 : issue_slots_4_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_lrs3 = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_lrs3 : issue_slots_4_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_ldst_val = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_ldst_val :
    issue_slots_4_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_dst_rtype = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_dst_rtype :
    issue_slots_4_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_lrs1_rtype = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_lrs1_rtype :
    issue_slots_4_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_lrs2_rtype = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_lrs2_rtype :
    issue_slots_4_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_frs3_en = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_frs3_en :
    issue_slots_4_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_fp_val = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_fp_val :
    issue_slots_4_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_fp_single = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_fp_single :
    issue_slots_4_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_xcpt_pf_if = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_xcpt_pf_if :
    issue_slots_4_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_xcpt_ae_if = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_xcpt_ae_if :
    issue_slots_4_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_xcpt_ma_if = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_xcpt_ma_if :
    issue_slots_4_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_bp_debug_if = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_bp_debug_if :
    issue_slots_4_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_bp_xcpt_if = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_bp_xcpt_if :
    issue_slots_4_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_debug_fsrc = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_debug_fsrc :
    issue_slots_4_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_3_io_in_uop_bits_debug_tsrc = _GEN_13[1:0] == 2'h2 ? issue_slots_5_out_uop_debug_tsrc :
    issue_slots_4_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_clock = clock;
  assign slots_4_reset = reset;
  assign slots_4_io_grant = issue_slots_4_request & _T_393 & ~_T_387; // @[issue-unit-age-ordered.scala 122:56]
  assign slots_4_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_4_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_4_io_clear = _GEN_11[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_4_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_4_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_4_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_4_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_4_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_4_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_4_io_in_uop_valid = _GEN_15[1:0] == 2'h2 ? issue_slots_6_will_be_valid : _GEN_822; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_4_io_in_uop_bits_switch = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_switch :
    issue_slots_5_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_switch_off = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_switch_off :
    issue_slots_5_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_unicore = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_is_unicore :
    issue_slots_5_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_shift = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_shift : issue_slots_5_out_uop_shift
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_lrs3_rtype = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_lrs3_rtype :
    issue_slots_5_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_rflag = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_rflag : issue_slots_5_out_uop_rflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_wflag = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_wflag : issue_slots_5_out_uop_wflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_prflag = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_prflag :
    issue_slots_5_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_pwflag = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_pwflag :
    issue_slots_5_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_pflag_busy = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_pflag_busy :
    issue_slots_5_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_stale_pflag = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_stale_pflag :
    issue_slots_5_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_op1_sel = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_op1_sel :
    issue_slots_5_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_op2_sel = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_op2_sel :
    issue_slots_5_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_split_num = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_split_num :
    issue_slots_5_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_self_index = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_self_index :
    issue_slots_5_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_rob_inst_idx = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_rob_inst_idx :
    issue_slots_5_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_address_num = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_address_num :
    issue_slots_5_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_uopc = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_uopc : issue_slots_5_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_inst = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_inst : issue_slots_5_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_debug_inst = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_debug_inst :
    issue_slots_5_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_rvc = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_is_rvc :
    issue_slots_5_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_debug_pc = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_debug_pc :
    issue_slots_5_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_iq_type = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_iq_type :
    issue_slots_5_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_fu_code = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_fu_code :
    issue_slots_5_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_br_type = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_br_type :
    issue_slots_5_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_op1_sel = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_op1_sel :
    issue_slots_5_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_op2_sel = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_op2_sel :
    issue_slots_5_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_imm_sel = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_imm_sel :
    issue_slots_5_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_op_fcn = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_op_fcn :
    issue_slots_5_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_fcn_dw = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_fcn_dw :
    issue_slots_5_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_csr_cmd = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_csr_cmd :
    issue_slots_5_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_is_load = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_is_load :
    issue_slots_5_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_is_sta = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_is_sta :
    issue_slots_5_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_is_std = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_is_std :
    issue_slots_5_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ctrl_op3_sel = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_ctrl_op3_sel :
    issue_slots_5_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_iw_state = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_iw_state :
    issue_slots_5_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_iw_p1_poisoned = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_iw_p1_poisoned :
    issue_slots_5_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_iw_p2_poisoned = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_iw_p2_poisoned :
    issue_slots_5_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_br = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_is_br : issue_slots_5_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_jalr = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_is_jalr :
    issue_slots_5_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_jal = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_is_jal :
    issue_slots_5_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_sfb = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_is_sfb :
    issue_slots_5_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_br_mask = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_br_mask :
    issue_slots_5_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_br_tag = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_br_tag :
    issue_slots_5_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ftq_idx = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_ftq_idx :
    issue_slots_5_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_edge_inst = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_edge_inst :
    issue_slots_5_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_pc_lob = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_pc_lob :
    issue_slots_5_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_taken = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_taken : issue_slots_5_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_imm_packed = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_imm_packed :
    issue_slots_5_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_csr_addr = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_csr_addr :
    issue_slots_5_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_rob_idx = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_rob_idx :
    issue_slots_5_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ldq_idx = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_ldq_idx :
    issue_slots_5_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_stq_idx = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_stq_idx :
    issue_slots_5_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_rxq_idx = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_rxq_idx :
    issue_slots_5_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_pdst = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_pdst : issue_slots_5_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_prs1 = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_prs1 : issue_slots_5_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_prs2 = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_prs2 : issue_slots_5_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_prs3 = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_prs3 : issue_slots_5_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ppred = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_ppred : issue_slots_5_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_prs1_busy = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_prs1_busy :
    issue_slots_5_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_prs2_busy = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_prs2_busy :
    issue_slots_5_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_prs3_busy = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_prs3_busy :
    issue_slots_5_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ppred_busy = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_ppred_busy :
    issue_slots_5_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_stale_pdst = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_stale_pdst :
    issue_slots_5_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_exception = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_exception :
    issue_slots_5_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_exc_cause = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_exc_cause :
    issue_slots_5_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_bypassable = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_bypassable :
    issue_slots_5_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_mem_cmd = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_mem_cmd :
    issue_slots_5_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_mem_size = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_mem_size :
    issue_slots_5_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_mem_signed = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_mem_signed :
    issue_slots_5_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_fence = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_is_fence :
    issue_slots_5_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_fencei = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_is_fencei :
    issue_slots_5_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_amo = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_is_amo :
    issue_slots_5_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_uses_ldq = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_uses_ldq :
    issue_slots_5_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_uses_stq = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_uses_stq :
    issue_slots_5_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_sys_pc2epc = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_is_sys_pc2epc :
    issue_slots_5_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_is_unique = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_is_unique :
    issue_slots_5_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_flush_on_commit = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_flush_on_commit :
    issue_slots_5_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ldst_is_rs1 = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_ldst_is_rs1 :
    issue_slots_5_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ldst = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_ldst : issue_slots_5_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_lrs1 = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_lrs1 : issue_slots_5_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_lrs2 = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_lrs2 : issue_slots_5_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_lrs3 = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_lrs3 : issue_slots_5_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_ldst_val = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_ldst_val :
    issue_slots_5_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_dst_rtype = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_dst_rtype :
    issue_slots_5_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_lrs1_rtype = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_lrs1_rtype :
    issue_slots_5_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_lrs2_rtype = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_lrs2_rtype :
    issue_slots_5_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_frs3_en = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_frs3_en :
    issue_slots_5_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_fp_val = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_fp_val :
    issue_slots_5_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_fp_single = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_fp_single :
    issue_slots_5_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_xcpt_pf_if = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_xcpt_pf_if :
    issue_slots_5_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_xcpt_ae_if = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_xcpt_ae_if :
    issue_slots_5_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_xcpt_ma_if = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_xcpt_ma_if :
    issue_slots_5_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_bp_debug_if = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_bp_debug_if :
    issue_slots_5_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_bp_xcpt_if = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_bp_xcpt_if :
    issue_slots_5_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_debug_fsrc = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_debug_fsrc :
    issue_slots_5_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_4_io_in_uop_bits_debug_tsrc = _GEN_15[1:0] == 2'h2 ? issue_slots_6_out_uop_debug_tsrc :
    issue_slots_5_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_clock = clock;
  assign slots_5_reset = reset;
  assign slots_5_io_grant = issue_slots_5_request & _T_408 & ~_T_402; // @[issue-unit-age-ordered.scala 122:56]
  assign slots_5_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_5_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_5_io_clear = _GEN_13[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_5_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_5_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_5_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_5_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_5_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_5_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_5_io_in_uop_valid = _GEN_17[1:0] == 2'h2 ? issue_slots_7_will_be_valid : _GEN_1018; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_5_io_in_uop_bits_switch = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_switch :
    issue_slots_6_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_switch_off = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_switch_off :
    issue_slots_6_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_unicore = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_is_unicore :
    issue_slots_6_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_shift = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_shift : issue_slots_6_out_uop_shift
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_lrs3_rtype = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_lrs3_rtype :
    issue_slots_6_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_rflag = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_rflag : issue_slots_6_out_uop_rflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_wflag = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_wflag : issue_slots_6_out_uop_wflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_prflag = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_prflag :
    issue_slots_6_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_pwflag = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_pwflag :
    issue_slots_6_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_pflag_busy = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_pflag_busy :
    issue_slots_6_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_stale_pflag = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_stale_pflag :
    issue_slots_6_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_op1_sel = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_op1_sel :
    issue_slots_6_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_op2_sel = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_op2_sel :
    issue_slots_6_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_split_num = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_split_num :
    issue_slots_6_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_self_index = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_self_index :
    issue_slots_6_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_rob_inst_idx = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_rob_inst_idx :
    issue_slots_6_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_address_num = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_address_num :
    issue_slots_6_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_uopc = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_uopc : issue_slots_6_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_inst = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_inst : issue_slots_6_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_debug_inst = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_debug_inst :
    issue_slots_6_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_rvc = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_is_rvc :
    issue_slots_6_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_debug_pc = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_debug_pc :
    issue_slots_6_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_iq_type = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_iq_type :
    issue_slots_6_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_fu_code = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_fu_code :
    issue_slots_6_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_br_type = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_br_type :
    issue_slots_6_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_op1_sel = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_op1_sel :
    issue_slots_6_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_op2_sel = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_op2_sel :
    issue_slots_6_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_imm_sel = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_imm_sel :
    issue_slots_6_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_op_fcn = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_op_fcn :
    issue_slots_6_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_fcn_dw = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_fcn_dw :
    issue_slots_6_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_csr_cmd = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_csr_cmd :
    issue_slots_6_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_is_load = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_is_load :
    issue_slots_6_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_is_sta = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_is_sta :
    issue_slots_6_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_is_std = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_is_std :
    issue_slots_6_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ctrl_op3_sel = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_ctrl_op3_sel :
    issue_slots_6_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_iw_state = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_iw_state :
    issue_slots_6_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_iw_p1_poisoned = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_iw_p1_poisoned :
    issue_slots_6_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_iw_p2_poisoned = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_iw_p2_poisoned :
    issue_slots_6_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_br = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_is_br : issue_slots_6_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_jalr = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_is_jalr :
    issue_slots_6_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_jal = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_is_jal :
    issue_slots_6_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_sfb = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_is_sfb :
    issue_slots_6_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_br_mask = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_br_mask :
    issue_slots_6_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_br_tag = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_br_tag :
    issue_slots_6_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ftq_idx = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_ftq_idx :
    issue_slots_6_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_edge_inst = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_edge_inst :
    issue_slots_6_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_pc_lob = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_pc_lob :
    issue_slots_6_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_taken = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_taken : issue_slots_6_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_imm_packed = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_imm_packed :
    issue_slots_6_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_csr_addr = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_csr_addr :
    issue_slots_6_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_rob_idx = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_rob_idx :
    issue_slots_6_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ldq_idx = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_ldq_idx :
    issue_slots_6_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_stq_idx = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_stq_idx :
    issue_slots_6_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_rxq_idx = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_rxq_idx :
    issue_slots_6_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_pdst = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_pdst : issue_slots_6_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_prs1 = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_prs1 : issue_slots_6_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_prs2 = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_prs2 : issue_slots_6_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_prs3 = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_prs3 : issue_slots_6_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ppred = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_ppred : issue_slots_6_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_prs1_busy = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_prs1_busy :
    issue_slots_6_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_prs2_busy = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_prs2_busy :
    issue_slots_6_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_prs3_busy = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_prs3_busy :
    issue_slots_6_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ppred_busy = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_ppred_busy :
    issue_slots_6_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_stale_pdst = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_stale_pdst :
    issue_slots_6_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_exception = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_exception :
    issue_slots_6_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_exc_cause = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_exc_cause :
    issue_slots_6_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_bypassable = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_bypassable :
    issue_slots_6_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_mem_cmd = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_mem_cmd :
    issue_slots_6_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_mem_size = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_mem_size :
    issue_slots_6_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_mem_signed = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_mem_signed :
    issue_slots_6_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_fence = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_is_fence :
    issue_slots_6_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_fencei = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_is_fencei :
    issue_slots_6_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_amo = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_is_amo :
    issue_slots_6_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_uses_ldq = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_uses_ldq :
    issue_slots_6_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_uses_stq = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_uses_stq :
    issue_slots_6_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_sys_pc2epc = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_is_sys_pc2epc :
    issue_slots_6_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_is_unique = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_is_unique :
    issue_slots_6_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_flush_on_commit = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_flush_on_commit :
    issue_slots_6_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ldst_is_rs1 = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_ldst_is_rs1 :
    issue_slots_6_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ldst = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_ldst : issue_slots_6_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_lrs1 = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_lrs1 : issue_slots_6_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_lrs2 = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_lrs2 : issue_slots_6_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_lrs3 = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_lrs3 : issue_slots_6_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_ldst_val = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_ldst_val :
    issue_slots_6_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_dst_rtype = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_dst_rtype :
    issue_slots_6_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_lrs1_rtype = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_lrs1_rtype :
    issue_slots_6_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_lrs2_rtype = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_lrs2_rtype :
    issue_slots_6_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_frs3_en = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_frs3_en :
    issue_slots_6_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_fp_val = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_fp_val :
    issue_slots_6_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_fp_single = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_fp_single :
    issue_slots_6_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_xcpt_pf_if = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_xcpt_pf_if :
    issue_slots_6_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_xcpt_ae_if = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_xcpt_ae_if :
    issue_slots_6_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_xcpt_ma_if = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_xcpt_ma_if :
    issue_slots_6_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_bp_debug_if = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_bp_debug_if :
    issue_slots_6_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_bp_xcpt_if = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_bp_xcpt_if :
    issue_slots_6_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_debug_fsrc = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_debug_fsrc :
    issue_slots_6_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_5_io_in_uop_bits_debug_tsrc = _GEN_17[1:0] == 2'h2 ? issue_slots_7_out_uop_debug_tsrc :
    issue_slots_6_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_clock = clock;
  assign slots_6_reset = reset;
  assign slots_6_io_grant = issue_slots_6_request & _T_423 & ~_T_417; // @[issue-unit-age-ordered.scala 122:56]
  assign slots_6_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_6_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_6_io_clear = _GEN_15[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_6_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_6_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_6_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_6_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_6_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_6_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_6_io_in_uop_valid = _GEN_19[1:0] == 2'h2 ? issue_slots_8_will_be_valid : _GEN_1214; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_6_io_in_uop_bits_switch = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_switch :
    issue_slots_7_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_switch_off = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_switch_off :
    issue_slots_7_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_unicore = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_is_unicore :
    issue_slots_7_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_shift = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_shift : issue_slots_7_out_uop_shift
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_lrs3_rtype = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_lrs3_rtype :
    issue_slots_7_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_rflag = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_rflag : issue_slots_7_out_uop_rflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_wflag = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_wflag : issue_slots_7_out_uop_wflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_prflag = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_prflag :
    issue_slots_7_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_pwflag = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_pwflag :
    issue_slots_7_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_pflag_busy = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_pflag_busy :
    issue_slots_7_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_stale_pflag = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_stale_pflag :
    issue_slots_7_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_op1_sel = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_op1_sel :
    issue_slots_7_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_op2_sel = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_op2_sel :
    issue_slots_7_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_split_num = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_split_num :
    issue_slots_7_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_self_index = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_self_index :
    issue_slots_7_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_rob_inst_idx = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_rob_inst_idx :
    issue_slots_7_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_address_num = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_address_num :
    issue_slots_7_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_uopc = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_uopc : issue_slots_7_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_inst = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_inst : issue_slots_7_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_debug_inst = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_debug_inst :
    issue_slots_7_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_rvc = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_is_rvc :
    issue_slots_7_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_debug_pc = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_debug_pc :
    issue_slots_7_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_iq_type = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_iq_type :
    issue_slots_7_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_fu_code = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_fu_code :
    issue_slots_7_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_br_type = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_br_type :
    issue_slots_7_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_op1_sel = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_op1_sel :
    issue_slots_7_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_op2_sel = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_op2_sel :
    issue_slots_7_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_imm_sel = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_imm_sel :
    issue_slots_7_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_op_fcn = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_op_fcn :
    issue_slots_7_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_fcn_dw = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_fcn_dw :
    issue_slots_7_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_csr_cmd = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_csr_cmd :
    issue_slots_7_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_is_load = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_is_load :
    issue_slots_7_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_is_sta = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_is_sta :
    issue_slots_7_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_is_std = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_is_std :
    issue_slots_7_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ctrl_op3_sel = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_ctrl_op3_sel :
    issue_slots_7_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_iw_state = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_iw_state :
    issue_slots_7_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_iw_p1_poisoned = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_iw_p1_poisoned :
    issue_slots_7_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_iw_p2_poisoned = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_iw_p2_poisoned :
    issue_slots_7_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_br = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_is_br : issue_slots_7_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_jalr = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_is_jalr :
    issue_slots_7_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_jal = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_is_jal :
    issue_slots_7_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_sfb = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_is_sfb :
    issue_slots_7_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_br_mask = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_br_mask :
    issue_slots_7_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_br_tag = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_br_tag :
    issue_slots_7_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ftq_idx = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_ftq_idx :
    issue_slots_7_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_edge_inst = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_edge_inst :
    issue_slots_7_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_pc_lob = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_pc_lob :
    issue_slots_7_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_taken = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_taken : issue_slots_7_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_imm_packed = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_imm_packed :
    issue_slots_7_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_csr_addr = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_csr_addr :
    issue_slots_7_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_rob_idx = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_rob_idx :
    issue_slots_7_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ldq_idx = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_ldq_idx :
    issue_slots_7_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_stq_idx = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_stq_idx :
    issue_slots_7_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_rxq_idx = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_rxq_idx :
    issue_slots_7_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_pdst = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_pdst : issue_slots_7_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_prs1 = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_prs1 : issue_slots_7_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_prs2 = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_prs2 : issue_slots_7_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_prs3 = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_prs3 : issue_slots_7_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ppred = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_ppred : issue_slots_7_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_prs1_busy = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_prs1_busy :
    issue_slots_7_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_prs2_busy = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_prs2_busy :
    issue_slots_7_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_prs3_busy = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_prs3_busy :
    issue_slots_7_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ppred_busy = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_ppred_busy :
    issue_slots_7_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_stale_pdst = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_stale_pdst :
    issue_slots_7_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_exception = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_exception :
    issue_slots_7_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_exc_cause = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_exc_cause :
    issue_slots_7_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_bypassable = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_bypassable :
    issue_slots_7_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_mem_cmd = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_mem_cmd :
    issue_slots_7_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_mem_size = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_mem_size :
    issue_slots_7_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_mem_signed = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_mem_signed :
    issue_slots_7_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_fence = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_is_fence :
    issue_slots_7_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_fencei = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_is_fencei :
    issue_slots_7_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_amo = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_is_amo :
    issue_slots_7_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_uses_ldq = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_uses_ldq :
    issue_slots_7_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_uses_stq = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_uses_stq :
    issue_slots_7_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_sys_pc2epc = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_is_sys_pc2epc :
    issue_slots_7_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_is_unique = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_is_unique :
    issue_slots_7_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_flush_on_commit = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_flush_on_commit :
    issue_slots_7_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ldst_is_rs1 = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_ldst_is_rs1 :
    issue_slots_7_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ldst = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_ldst : issue_slots_7_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_lrs1 = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_lrs1 : issue_slots_7_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_lrs2 = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_lrs2 : issue_slots_7_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_lrs3 = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_lrs3 : issue_slots_7_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_ldst_val = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_ldst_val :
    issue_slots_7_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_dst_rtype = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_dst_rtype :
    issue_slots_7_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_lrs1_rtype = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_lrs1_rtype :
    issue_slots_7_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_lrs2_rtype = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_lrs2_rtype :
    issue_slots_7_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_frs3_en = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_frs3_en :
    issue_slots_7_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_fp_val = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_fp_val :
    issue_slots_7_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_fp_single = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_fp_single :
    issue_slots_7_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_xcpt_pf_if = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_xcpt_pf_if :
    issue_slots_7_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_xcpt_ae_if = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_xcpt_ae_if :
    issue_slots_7_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_xcpt_ma_if = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_xcpt_ma_if :
    issue_slots_7_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_bp_debug_if = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_bp_debug_if :
    issue_slots_7_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_bp_xcpt_if = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_bp_xcpt_if :
    issue_slots_7_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_debug_fsrc = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_debug_fsrc :
    issue_slots_7_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_6_io_in_uop_bits_debug_tsrc = _GEN_19[1:0] == 2'h2 ? issue_slots_8_out_uop_debug_tsrc :
    issue_slots_7_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_clock = clock;
  assign slots_7_reset = reset;
  assign slots_7_io_grant = issue_slots_7_request & _T_438 & ~_T_432; // @[issue-unit-age-ordered.scala 122:56]
  assign slots_7_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_7_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_7_io_clear = _GEN_17[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_7_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_7_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_7_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_7_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_7_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_7_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_7_io_in_uop_valid = _GEN_21[1:0] == 2'h2 ? issue_slots_9_will_be_valid : _GEN_1410; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_7_io_in_uop_bits_switch = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_switch :
    issue_slots_8_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_switch_off = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_switch_off :
    issue_slots_8_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_unicore = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_is_unicore :
    issue_slots_8_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_shift = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_shift : issue_slots_8_out_uop_shift
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_lrs3_rtype = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_lrs3_rtype :
    issue_slots_8_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_rflag = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_rflag : issue_slots_8_out_uop_rflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_wflag = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_wflag : issue_slots_8_out_uop_wflag
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_prflag = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_prflag :
    issue_slots_8_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_pwflag = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_pwflag :
    issue_slots_8_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_pflag_busy = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_pflag_busy :
    issue_slots_8_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_stale_pflag = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_stale_pflag :
    issue_slots_8_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_op1_sel = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_op1_sel :
    issue_slots_8_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_op2_sel = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_op2_sel :
    issue_slots_8_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_split_num = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_split_num :
    issue_slots_8_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_self_index = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_self_index :
    issue_slots_8_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_rob_inst_idx = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_rob_inst_idx :
    issue_slots_8_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_address_num = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_address_num :
    issue_slots_8_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_uopc = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_uopc : issue_slots_8_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_inst = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_inst : issue_slots_8_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_debug_inst = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_debug_inst :
    issue_slots_8_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_rvc = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_is_rvc :
    issue_slots_8_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_debug_pc = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_debug_pc :
    issue_slots_8_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_iq_type = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_iq_type :
    issue_slots_8_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_fu_code = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_fu_code :
    issue_slots_8_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_br_type = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_br_type :
    issue_slots_8_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_op1_sel = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_op1_sel :
    issue_slots_8_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_op2_sel = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_op2_sel :
    issue_slots_8_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_imm_sel = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_imm_sel :
    issue_slots_8_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_op_fcn = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_op_fcn :
    issue_slots_8_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_fcn_dw = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_fcn_dw :
    issue_slots_8_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_csr_cmd = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_csr_cmd :
    issue_slots_8_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_is_load = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_is_load :
    issue_slots_8_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_is_sta = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_is_sta :
    issue_slots_8_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_is_std = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_is_std :
    issue_slots_8_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ctrl_op3_sel = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_ctrl_op3_sel :
    issue_slots_8_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_iw_state = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_iw_state :
    issue_slots_8_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_iw_p1_poisoned = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_iw_p1_poisoned :
    issue_slots_8_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_iw_p2_poisoned = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_iw_p2_poisoned :
    issue_slots_8_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_br = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_is_br : issue_slots_8_out_uop_is_br
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_jalr = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_is_jalr :
    issue_slots_8_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_jal = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_is_jal :
    issue_slots_8_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_sfb = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_is_sfb :
    issue_slots_8_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_br_mask = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_br_mask :
    issue_slots_8_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_br_tag = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_br_tag :
    issue_slots_8_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ftq_idx = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_ftq_idx :
    issue_slots_8_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_edge_inst = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_edge_inst :
    issue_slots_8_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_pc_lob = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_pc_lob :
    issue_slots_8_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_taken = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_taken : issue_slots_8_out_uop_taken
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_imm_packed = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_imm_packed :
    issue_slots_8_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_csr_addr = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_csr_addr :
    issue_slots_8_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_rob_idx = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_rob_idx :
    issue_slots_8_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ldq_idx = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_ldq_idx :
    issue_slots_8_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_stq_idx = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_stq_idx :
    issue_slots_8_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_rxq_idx = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_rxq_idx :
    issue_slots_8_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_pdst = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_pdst : issue_slots_8_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_prs1 = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_prs1 : issue_slots_8_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_prs2 = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_prs2 : issue_slots_8_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_prs3 = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_prs3 : issue_slots_8_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ppred = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_ppred : issue_slots_8_out_uop_ppred
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_prs1_busy = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_prs1_busy :
    issue_slots_8_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_prs2_busy = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_prs2_busy :
    issue_slots_8_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_prs3_busy = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_prs3_busy :
    issue_slots_8_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ppred_busy = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_ppred_busy :
    issue_slots_8_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_stale_pdst = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_stale_pdst :
    issue_slots_8_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_exception = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_exception :
    issue_slots_8_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_exc_cause = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_exc_cause :
    issue_slots_8_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_bypassable = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_bypassable :
    issue_slots_8_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_mem_cmd = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_mem_cmd :
    issue_slots_8_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_mem_size = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_mem_size :
    issue_slots_8_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_mem_signed = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_mem_signed :
    issue_slots_8_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_fence = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_is_fence :
    issue_slots_8_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_fencei = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_is_fencei :
    issue_slots_8_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_amo = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_is_amo :
    issue_slots_8_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_uses_ldq = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_uses_ldq :
    issue_slots_8_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_uses_stq = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_uses_stq :
    issue_slots_8_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_sys_pc2epc = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_is_sys_pc2epc :
    issue_slots_8_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_is_unique = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_is_unique :
    issue_slots_8_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_flush_on_commit = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_flush_on_commit :
    issue_slots_8_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ldst_is_rs1 = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_ldst_is_rs1 :
    issue_slots_8_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ldst = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_ldst : issue_slots_8_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_lrs1 = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_lrs1 : issue_slots_8_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_lrs2 = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_lrs2 : issue_slots_8_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_lrs3 = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_lrs3 : issue_slots_8_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_ldst_val = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_ldst_val :
    issue_slots_8_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_dst_rtype = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_dst_rtype :
    issue_slots_8_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_lrs1_rtype = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_lrs1_rtype :
    issue_slots_8_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_lrs2_rtype = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_lrs2_rtype :
    issue_slots_8_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_frs3_en = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_frs3_en :
    issue_slots_8_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_fp_val = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_fp_val :
    issue_slots_8_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_fp_single = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_fp_single :
    issue_slots_8_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_xcpt_pf_if = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_xcpt_pf_if :
    issue_slots_8_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_xcpt_ae_if = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_xcpt_ae_if :
    issue_slots_8_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_xcpt_ma_if = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_xcpt_ma_if :
    issue_slots_8_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_bp_debug_if = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_bp_debug_if :
    issue_slots_8_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_bp_xcpt_if = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_bp_xcpt_if :
    issue_slots_8_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_debug_fsrc = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_debug_fsrc :
    issue_slots_8_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_7_io_in_uop_bits_debug_tsrc = _GEN_21[1:0] == 2'h2 ? issue_slots_9_out_uop_debug_tsrc :
    issue_slots_8_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_clock = clock;
  assign slots_8_reset = reset;
  assign slots_8_io_grant = issue_slots_8_request & _T_453 & ~_T_447; // @[issue-unit-age-ordered.scala 122:56]
  assign slots_8_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_8_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_8_io_clear = _GEN_19[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_8_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_8_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_8_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_8_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_8_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_8_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_8_io_in_uop_valid = _GEN_23[1:0] == 2'h2 ? issue_slots_10_will_be_valid : _GEN_1606; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_8_io_in_uop_bits_switch = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_switch :
    issue_slots_9_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_switch_off = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_switch_off :
    issue_slots_9_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_unicore = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_is_unicore :
    issue_slots_9_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_shift = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_shift :
    issue_slots_9_out_uop_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_lrs3_rtype = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_lrs3_rtype :
    issue_slots_9_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_rflag = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_rflag :
    issue_slots_9_out_uop_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_wflag = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_wflag :
    issue_slots_9_out_uop_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_prflag = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_prflag :
    issue_slots_9_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_pwflag = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_pwflag :
    issue_slots_9_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_pflag_busy = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_pflag_busy :
    issue_slots_9_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_stale_pflag = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_stale_pflag :
    issue_slots_9_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_op1_sel = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_op1_sel :
    issue_slots_9_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_op2_sel = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_op2_sel :
    issue_slots_9_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_split_num = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_split_num :
    issue_slots_9_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_self_index = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_self_index :
    issue_slots_9_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_rob_inst_idx = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_rob_inst_idx :
    issue_slots_9_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_address_num = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_address_num :
    issue_slots_9_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_uopc = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_uopc : issue_slots_9_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_inst = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_inst : issue_slots_9_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_debug_inst = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_debug_inst :
    issue_slots_9_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_rvc = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_is_rvc :
    issue_slots_9_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_debug_pc = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_debug_pc :
    issue_slots_9_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_iq_type = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_iq_type :
    issue_slots_9_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_fu_code = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_fu_code :
    issue_slots_9_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_br_type = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_br_type :
    issue_slots_9_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_op1_sel = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_op1_sel :
    issue_slots_9_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_op2_sel = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_op2_sel :
    issue_slots_9_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_imm_sel = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_imm_sel :
    issue_slots_9_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_op_fcn = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_op_fcn :
    issue_slots_9_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_fcn_dw = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_fcn_dw :
    issue_slots_9_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_csr_cmd = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_csr_cmd :
    issue_slots_9_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_is_load = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_is_load :
    issue_slots_9_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_is_sta = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_is_sta :
    issue_slots_9_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_is_std = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_is_std :
    issue_slots_9_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ctrl_op3_sel = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_ctrl_op3_sel :
    issue_slots_9_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_iw_state = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_iw_state :
    issue_slots_9_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_iw_p1_poisoned = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_iw_p1_poisoned :
    issue_slots_9_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_iw_p2_poisoned = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_iw_p2_poisoned :
    issue_slots_9_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_br = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_is_br :
    issue_slots_9_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_jalr = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_is_jalr :
    issue_slots_9_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_jal = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_is_jal :
    issue_slots_9_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_sfb = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_is_sfb :
    issue_slots_9_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_br_mask = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_br_mask :
    issue_slots_9_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_br_tag = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_br_tag :
    issue_slots_9_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ftq_idx = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_ftq_idx :
    issue_slots_9_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_edge_inst = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_edge_inst :
    issue_slots_9_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_pc_lob = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_pc_lob :
    issue_slots_9_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_taken = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_taken :
    issue_slots_9_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_imm_packed = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_imm_packed :
    issue_slots_9_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_csr_addr = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_csr_addr :
    issue_slots_9_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_rob_idx = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_rob_idx :
    issue_slots_9_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ldq_idx = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_ldq_idx :
    issue_slots_9_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_stq_idx = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_stq_idx :
    issue_slots_9_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_rxq_idx = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_rxq_idx :
    issue_slots_9_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_pdst = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_pdst : issue_slots_9_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_prs1 = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_prs1 : issue_slots_9_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_prs2 = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_prs2 : issue_slots_9_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_prs3 = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_prs3 : issue_slots_9_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ppred = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_ppred :
    issue_slots_9_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_prs1_busy = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_prs1_busy :
    issue_slots_9_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_prs2_busy = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_prs2_busy :
    issue_slots_9_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_prs3_busy = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_prs3_busy :
    issue_slots_9_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ppred_busy = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_ppred_busy :
    issue_slots_9_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_stale_pdst = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_stale_pdst :
    issue_slots_9_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_exception = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_exception :
    issue_slots_9_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_exc_cause = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_exc_cause :
    issue_slots_9_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_bypassable = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_bypassable :
    issue_slots_9_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_mem_cmd = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_mem_cmd :
    issue_slots_9_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_mem_size = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_mem_size :
    issue_slots_9_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_mem_signed = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_mem_signed :
    issue_slots_9_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_fence = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_is_fence :
    issue_slots_9_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_fencei = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_is_fencei :
    issue_slots_9_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_amo = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_is_amo :
    issue_slots_9_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_uses_ldq = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_uses_ldq :
    issue_slots_9_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_uses_stq = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_uses_stq :
    issue_slots_9_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_sys_pc2epc = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_is_sys_pc2epc :
    issue_slots_9_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_is_unique = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_is_unique :
    issue_slots_9_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_flush_on_commit = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_flush_on_commit :
    issue_slots_9_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ldst_is_rs1 = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_ldst_is_rs1 :
    issue_slots_9_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ldst = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_ldst : issue_slots_9_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_lrs1 = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_lrs1 : issue_slots_9_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_lrs2 = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_lrs2 : issue_slots_9_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_lrs3 = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_lrs3 : issue_slots_9_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_ldst_val = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_ldst_val :
    issue_slots_9_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_dst_rtype = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_dst_rtype :
    issue_slots_9_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_lrs1_rtype = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_lrs1_rtype :
    issue_slots_9_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_lrs2_rtype = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_lrs2_rtype :
    issue_slots_9_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_frs3_en = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_frs3_en :
    issue_slots_9_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_fp_val = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_fp_val :
    issue_slots_9_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_fp_single = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_fp_single :
    issue_slots_9_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_xcpt_pf_if = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_xcpt_pf_if :
    issue_slots_9_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_xcpt_ae_if = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_xcpt_ae_if :
    issue_slots_9_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_xcpt_ma_if = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_xcpt_ma_if :
    issue_slots_9_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_bp_debug_if = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_bp_debug_if :
    issue_slots_9_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_bp_xcpt_if = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_bp_xcpt_if :
    issue_slots_9_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_debug_fsrc = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_debug_fsrc :
    issue_slots_9_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_8_io_in_uop_bits_debug_tsrc = _GEN_23[1:0] == 2'h2 ? issue_slots_10_out_uop_debug_tsrc :
    issue_slots_9_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_clock = clock;
  assign slots_9_reset = reset;
  assign slots_9_io_grant = issue_slots_9_request & _T_468 & ~_T_462; // @[issue-unit-age-ordered.scala 122:56]
  assign slots_9_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_9_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_9_io_clear = _GEN_21[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_9_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_9_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_9_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_9_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_9_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_9_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_9_io_in_uop_valid = _GEN_25[1:0] == 2'h2 ? issue_slots_11_will_be_valid : _GEN_1802; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_9_io_in_uop_bits_switch = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_switch :
    issue_slots_10_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_switch_off = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_switch_off :
    issue_slots_10_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_unicore = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_is_unicore :
    issue_slots_10_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_shift = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_shift :
    issue_slots_10_out_uop_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_lrs3_rtype = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_lrs3_rtype :
    issue_slots_10_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_rflag = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_rflag :
    issue_slots_10_out_uop_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_wflag = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_wflag :
    issue_slots_10_out_uop_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_prflag = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_prflag :
    issue_slots_10_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_pwflag = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_pwflag :
    issue_slots_10_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_pflag_busy = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_pflag_busy :
    issue_slots_10_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_stale_pflag = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_stale_pflag :
    issue_slots_10_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_op1_sel = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_op1_sel :
    issue_slots_10_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_op2_sel = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_op2_sel :
    issue_slots_10_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_split_num = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_split_num :
    issue_slots_10_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_self_index = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_self_index :
    issue_slots_10_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_rob_inst_idx = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_rob_inst_idx :
    issue_slots_10_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_address_num = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_address_num :
    issue_slots_10_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_uopc = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_uopc : issue_slots_10_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_inst = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_inst : issue_slots_10_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_debug_inst = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_debug_inst :
    issue_slots_10_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_rvc = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_is_rvc :
    issue_slots_10_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_debug_pc = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_debug_pc :
    issue_slots_10_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_iq_type = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_iq_type :
    issue_slots_10_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_fu_code = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_fu_code :
    issue_slots_10_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_br_type = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_br_type :
    issue_slots_10_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_op1_sel = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_op1_sel :
    issue_slots_10_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_op2_sel = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_op2_sel :
    issue_slots_10_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_imm_sel = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_imm_sel :
    issue_slots_10_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_op_fcn = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_op_fcn :
    issue_slots_10_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_fcn_dw = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_fcn_dw :
    issue_slots_10_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_csr_cmd = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_csr_cmd :
    issue_slots_10_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_is_load = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_is_load :
    issue_slots_10_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_is_sta = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_is_sta :
    issue_slots_10_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_is_std = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_is_std :
    issue_slots_10_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ctrl_op3_sel = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_ctrl_op3_sel :
    issue_slots_10_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_iw_state = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_iw_state :
    issue_slots_10_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_iw_p1_poisoned = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_iw_p1_poisoned :
    issue_slots_10_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_iw_p2_poisoned = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_iw_p2_poisoned :
    issue_slots_10_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_br = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_is_br :
    issue_slots_10_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_jalr = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_is_jalr :
    issue_slots_10_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_jal = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_is_jal :
    issue_slots_10_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_sfb = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_is_sfb :
    issue_slots_10_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_br_mask = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_br_mask :
    issue_slots_10_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_br_tag = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_br_tag :
    issue_slots_10_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ftq_idx = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_ftq_idx :
    issue_slots_10_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_edge_inst = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_edge_inst :
    issue_slots_10_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_pc_lob = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_pc_lob :
    issue_slots_10_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_taken = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_taken :
    issue_slots_10_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_imm_packed = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_imm_packed :
    issue_slots_10_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_csr_addr = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_csr_addr :
    issue_slots_10_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_rob_idx = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_rob_idx :
    issue_slots_10_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ldq_idx = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_ldq_idx :
    issue_slots_10_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_stq_idx = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_stq_idx :
    issue_slots_10_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_rxq_idx = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_rxq_idx :
    issue_slots_10_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_pdst = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_pdst : issue_slots_10_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_prs1 = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_prs1 : issue_slots_10_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_prs2 = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_prs2 : issue_slots_10_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_prs3 = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_prs3 : issue_slots_10_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ppred = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_ppred :
    issue_slots_10_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_prs1_busy = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_prs1_busy :
    issue_slots_10_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_prs2_busy = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_prs2_busy :
    issue_slots_10_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_prs3_busy = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_prs3_busy :
    issue_slots_10_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ppred_busy = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_ppred_busy :
    issue_slots_10_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_stale_pdst = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_stale_pdst :
    issue_slots_10_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_exception = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_exception :
    issue_slots_10_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_exc_cause = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_exc_cause :
    issue_slots_10_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_bypassable = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_bypassable :
    issue_slots_10_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_mem_cmd = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_mem_cmd :
    issue_slots_10_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_mem_size = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_mem_size :
    issue_slots_10_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_mem_signed = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_mem_signed :
    issue_slots_10_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_fence = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_is_fence :
    issue_slots_10_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_fencei = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_is_fencei :
    issue_slots_10_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_amo = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_is_amo :
    issue_slots_10_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_uses_ldq = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_uses_ldq :
    issue_slots_10_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_uses_stq = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_uses_stq :
    issue_slots_10_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_sys_pc2epc = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_is_sys_pc2epc :
    issue_slots_10_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_is_unique = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_is_unique :
    issue_slots_10_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_flush_on_commit = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_flush_on_commit :
    issue_slots_10_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ldst_is_rs1 = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_ldst_is_rs1 :
    issue_slots_10_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ldst = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_ldst : issue_slots_10_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_lrs1 = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_lrs1 : issue_slots_10_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_lrs2 = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_lrs2 : issue_slots_10_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_lrs3 = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_lrs3 : issue_slots_10_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_ldst_val = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_ldst_val :
    issue_slots_10_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_dst_rtype = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_dst_rtype :
    issue_slots_10_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_lrs1_rtype = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_lrs1_rtype :
    issue_slots_10_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_lrs2_rtype = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_lrs2_rtype :
    issue_slots_10_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_frs3_en = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_frs3_en :
    issue_slots_10_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_fp_val = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_fp_val :
    issue_slots_10_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_fp_single = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_fp_single :
    issue_slots_10_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_xcpt_pf_if = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_xcpt_pf_if :
    issue_slots_10_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_xcpt_ae_if = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_xcpt_ae_if :
    issue_slots_10_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_xcpt_ma_if = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_xcpt_ma_if :
    issue_slots_10_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_bp_debug_if = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_bp_debug_if :
    issue_slots_10_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_bp_xcpt_if = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_bp_xcpt_if :
    issue_slots_10_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_debug_fsrc = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_debug_fsrc :
    issue_slots_10_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_9_io_in_uop_bits_debug_tsrc = _GEN_25[1:0] == 2'h2 ? issue_slots_11_out_uop_debug_tsrc :
    issue_slots_10_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_clock = clock;
  assign slots_10_reset = reset;
  assign slots_10_io_grant = issue_slots_10_request & _T_483 & ~_T_477; // @[issue-unit-age-ordered.scala 122:56]
  assign slots_10_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_10_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_10_io_clear = _GEN_23[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_10_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_10_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_10_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_10_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_10_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_10_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_10_io_in_uop_valid = _GEN_27[1:0] == 2'h2 ? issue_slots_12_will_be_valid : _GEN_1998; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_10_io_in_uop_bits_switch = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_switch :
    issue_slots_11_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_switch_off = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_switch_off :
    issue_slots_11_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_unicore = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_is_unicore :
    issue_slots_11_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_shift = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_shift :
    issue_slots_11_out_uop_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_lrs3_rtype = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_lrs3_rtype :
    issue_slots_11_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_rflag = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_rflag :
    issue_slots_11_out_uop_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_wflag = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_wflag :
    issue_slots_11_out_uop_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_prflag = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_prflag :
    issue_slots_11_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_pwflag = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_pwflag :
    issue_slots_11_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_pflag_busy = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_pflag_busy :
    issue_slots_11_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_stale_pflag = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_stale_pflag :
    issue_slots_11_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_op1_sel = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_op1_sel :
    issue_slots_11_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_op2_sel = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_op2_sel :
    issue_slots_11_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_split_num = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_split_num :
    issue_slots_11_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_self_index = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_self_index :
    issue_slots_11_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_rob_inst_idx = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_rob_inst_idx :
    issue_slots_11_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_address_num = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_address_num :
    issue_slots_11_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_uopc = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_uopc : issue_slots_11_out_uop_uopc
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_inst = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_inst : issue_slots_11_out_uop_inst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_debug_inst = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_debug_inst :
    issue_slots_11_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_rvc = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_is_rvc :
    issue_slots_11_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_debug_pc = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_debug_pc :
    issue_slots_11_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_iq_type = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_iq_type :
    issue_slots_11_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_fu_code = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_fu_code :
    issue_slots_11_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_br_type = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_br_type :
    issue_slots_11_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_op1_sel = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_op1_sel :
    issue_slots_11_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_op2_sel = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_op2_sel :
    issue_slots_11_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_imm_sel = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_imm_sel :
    issue_slots_11_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_op_fcn = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_op_fcn :
    issue_slots_11_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_fcn_dw = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_fcn_dw :
    issue_slots_11_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_csr_cmd = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_csr_cmd :
    issue_slots_11_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_is_load = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_is_load :
    issue_slots_11_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_is_sta = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_is_sta :
    issue_slots_11_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_is_std = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_is_std :
    issue_slots_11_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ctrl_op3_sel = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_ctrl_op3_sel :
    issue_slots_11_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_iw_state = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_iw_state :
    issue_slots_11_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_iw_p1_poisoned = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_iw_p1_poisoned :
    issue_slots_11_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_iw_p2_poisoned = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_iw_p2_poisoned :
    issue_slots_11_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_br = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_is_br :
    issue_slots_11_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_jalr = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_is_jalr :
    issue_slots_11_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_jal = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_is_jal :
    issue_slots_11_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_sfb = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_is_sfb :
    issue_slots_11_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_br_mask = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_br_mask :
    issue_slots_11_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_br_tag = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_br_tag :
    issue_slots_11_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ftq_idx = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_ftq_idx :
    issue_slots_11_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_edge_inst = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_edge_inst :
    issue_slots_11_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_pc_lob = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_pc_lob :
    issue_slots_11_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_taken = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_taken :
    issue_slots_11_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_imm_packed = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_imm_packed :
    issue_slots_11_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_csr_addr = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_csr_addr :
    issue_slots_11_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_rob_idx = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_rob_idx :
    issue_slots_11_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ldq_idx = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_ldq_idx :
    issue_slots_11_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_stq_idx = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_stq_idx :
    issue_slots_11_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_rxq_idx = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_rxq_idx :
    issue_slots_11_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_pdst = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_pdst : issue_slots_11_out_uop_pdst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_prs1 = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_prs1 : issue_slots_11_out_uop_prs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_prs2 = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_prs2 : issue_slots_11_out_uop_prs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_prs3 = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_prs3 : issue_slots_11_out_uop_prs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ppred = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_ppred :
    issue_slots_11_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_prs1_busy = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_prs1_busy :
    issue_slots_11_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_prs2_busy = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_prs2_busy :
    issue_slots_11_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_prs3_busy = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_prs3_busy :
    issue_slots_11_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ppred_busy = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_ppred_busy :
    issue_slots_11_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_stale_pdst = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_stale_pdst :
    issue_slots_11_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_exception = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_exception :
    issue_slots_11_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_exc_cause = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_exc_cause :
    issue_slots_11_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_bypassable = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_bypassable :
    issue_slots_11_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_mem_cmd = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_mem_cmd :
    issue_slots_11_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_mem_size = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_mem_size :
    issue_slots_11_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_mem_signed = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_mem_signed :
    issue_slots_11_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_fence = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_is_fence :
    issue_slots_11_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_fencei = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_is_fencei :
    issue_slots_11_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_amo = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_is_amo :
    issue_slots_11_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_uses_ldq = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_uses_ldq :
    issue_slots_11_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_uses_stq = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_uses_stq :
    issue_slots_11_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_sys_pc2epc = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_is_sys_pc2epc :
    issue_slots_11_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_is_unique = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_is_unique :
    issue_slots_11_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_flush_on_commit = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_flush_on_commit :
    issue_slots_11_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ldst_is_rs1 = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_ldst_is_rs1 :
    issue_slots_11_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ldst = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_ldst : issue_slots_11_out_uop_ldst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_lrs1 = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_lrs1 : issue_slots_11_out_uop_lrs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_lrs2 = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_lrs2 : issue_slots_11_out_uop_lrs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_lrs3 = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_lrs3 : issue_slots_11_out_uop_lrs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_ldst_val = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_ldst_val :
    issue_slots_11_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_dst_rtype = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_dst_rtype :
    issue_slots_11_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_lrs1_rtype = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_lrs1_rtype :
    issue_slots_11_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_lrs2_rtype = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_lrs2_rtype :
    issue_slots_11_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_frs3_en = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_frs3_en :
    issue_slots_11_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_fp_val = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_fp_val :
    issue_slots_11_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_fp_single = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_fp_single :
    issue_slots_11_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_xcpt_pf_if = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_xcpt_pf_if :
    issue_slots_11_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_xcpt_ae_if = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_xcpt_ae_if :
    issue_slots_11_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_xcpt_ma_if = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_xcpt_ma_if :
    issue_slots_11_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_bp_debug_if = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_bp_debug_if :
    issue_slots_11_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_bp_xcpt_if = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_bp_xcpt_if :
    issue_slots_11_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_debug_fsrc = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_debug_fsrc :
    issue_slots_11_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_10_io_in_uop_bits_debug_tsrc = _GEN_27[1:0] == 2'h2 ? issue_slots_12_out_uop_debug_tsrc :
    issue_slots_11_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_clock = clock;
  assign slots_11_reset = reset;
  assign slots_11_io_grant = issue_slots_11_request & _T_498 & ~_T_492; // @[issue-unit-age-ordered.scala 122:56]
  assign slots_11_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_11_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_11_io_clear = _GEN_25[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_11_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_11_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_11_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_11_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_11_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_11_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_11_io_in_uop_valid = _GEN_29[1:0] == 2'h2 ? issue_slots_13_will_be_valid : _GEN_2194; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_11_io_in_uop_bits_switch = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_switch :
    issue_slots_12_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_switch_off = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_switch_off :
    issue_slots_12_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_unicore = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_is_unicore :
    issue_slots_12_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_shift = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_shift :
    issue_slots_12_out_uop_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_lrs3_rtype = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_lrs3_rtype :
    issue_slots_12_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_rflag = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_rflag :
    issue_slots_12_out_uop_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_wflag = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_wflag :
    issue_slots_12_out_uop_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_prflag = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_prflag :
    issue_slots_12_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_pwflag = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_pwflag :
    issue_slots_12_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_pflag_busy = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_pflag_busy :
    issue_slots_12_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_stale_pflag = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_stale_pflag :
    issue_slots_12_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_op1_sel = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_op1_sel :
    issue_slots_12_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_op2_sel = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_op2_sel :
    issue_slots_12_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_split_num = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_split_num :
    issue_slots_12_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_self_index = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_self_index :
    issue_slots_12_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_rob_inst_idx = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_rob_inst_idx :
    issue_slots_12_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_address_num = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_address_num :
    issue_slots_12_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_uopc = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_uopc : issue_slots_12_out_uop_uopc
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_inst = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_inst : issue_slots_12_out_uop_inst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_debug_inst = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_debug_inst :
    issue_slots_12_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_rvc = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_is_rvc :
    issue_slots_12_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_debug_pc = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_debug_pc :
    issue_slots_12_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_iq_type = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_iq_type :
    issue_slots_12_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_fu_code = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_fu_code :
    issue_slots_12_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_br_type = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_br_type :
    issue_slots_12_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_op1_sel = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_op1_sel :
    issue_slots_12_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_op2_sel = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_op2_sel :
    issue_slots_12_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_imm_sel = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_imm_sel :
    issue_slots_12_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_op_fcn = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_op_fcn :
    issue_slots_12_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_fcn_dw = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_fcn_dw :
    issue_slots_12_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_csr_cmd = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_csr_cmd :
    issue_slots_12_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_is_load = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_is_load :
    issue_slots_12_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_is_sta = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_is_sta :
    issue_slots_12_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_is_std = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_is_std :
    issue_slots_12_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ctrl_op3_sel = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_ctrl_op3_sel :
    issue_slots_12_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_iw_state = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_iw_state :
    issue_slots_12_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_iw_p1_poisoned = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_iw_p1_poisoned :
    issue_slots_12_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_iw_p2_poisoned = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_iw_p2_poisoned :
    issue_slots_12_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_br = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_is_br :
    issue_slots_12_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_jalr = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_is_jalr :
    issue_slots_12_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_jal = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_is_jal :
    issue_slots_12_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_sfb = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_is_sfb :
    issue_slots_12_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_br_mask = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_br_mask :
    issue_slots_12_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_br_tag = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_br_tag :
    issue_slots_12_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ftq_idx = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_ftq_idx :
    issue_slots_12_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_edge_inst = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_edge_inst :
    issue_slots_12_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_pc_lob = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_pc_lob :
    issue_slots_12_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_taken = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_taken :
    issue_slots_12_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_imm_packed = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_imm_packed :
    issue_slots_12_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_csr_addr = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_csr_addr :
    issue_slots_12_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_rob_idx = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_rob_idx :
    issue_slots_12_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ldq_idx = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_ldq_idx :
    issue_slots_12_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_stq_idx = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_stq_idx :
    issue_slots_12_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_rxq_idx = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_rxq_idx :
    issue_slots_12_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_pdst = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_pdst : issue_slots_12_out_uop_pdst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_prs1 = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_prs1 : issue_slots_12_out_uop_prs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_prs2 = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_prs2 : issue_slots_12_out_uop_prs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_prs3 = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_prs3 : issue_slots_12_out_uop_prs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ppred = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_ppred :
    issue_slots_12_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_prs1_busy = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_prs1_busy :
    issue_slots_12_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_prs2_busy = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_prs2_busy :
    issue_slots_12_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_prs3_busy = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_prs3_busy :
    issue_slots_12_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ppred_busy = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_ppred_busy :
    issue_slots_12_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_stale_pdst = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_stale_pdst :
    issue_slots_12_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_exception = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_exception :
    issue_slots_12_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_exc_cause = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_exc_cause :
    issue_slots_12_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_bypassable = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_bypassable :
    issue_slots_12_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_mem_cmd = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_mem_cmd :
    issue_slots_12_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_mem_size = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_mem_size :
    issue_slots_12_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_mem_signed = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_mem_signed :
    issue_slots_12_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_fence = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_is_fence :
    issue_slots_12_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_fencei = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_is_fencei :
    issue_slots_12_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_amo = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_is_amo :
    issue_slots_12_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_uses_ldq = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_uses_ldq :
    issue_slots_12_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_uses_stq = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_uses_stq :
    issue_slots_12_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_sys_pc2epc = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_is_sys_pc2epc :
    issue_slots_12_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_is_unique = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_is_unique :
    issue_slots_12_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_flush_on_commit = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_flush_on_commit :
    issue_slots_12_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ldst_is_rs1 = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_ldst_is_rs1 :
    issue_slots_12_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ldst = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_ldst : issue_slots_12_out_uop_ldst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_lrs1 = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_lrs1 : issue_slots_12_out_uop_lrs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_lrs2 = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_lrs2 : issue_slots_12_out_uop_lrs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_lrs3 = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_lrs3 : issue_slots_12_out_uop_lrs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_ldst_val = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_ldst_val :
    issue_slots_12_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_dst_rtype = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_dst_rtype :
    issue_slots_12_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_lrs1_rtype = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_lrs1_rtype :
    issue_slots_12_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_lrs2_rtype = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_lrs2_rtype :
    issue_slots_12_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_frs3_en = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_frs3_en :
    issue_slots_12_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_fp_val = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_fp_val :
    issue_slots_12_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_fp_single = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_fp_single :
    issue_slots_12_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_xcpt_pf_if = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_xcpt_pf_if :
    issue_slots_12_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_xcpt_ae_if = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_xcpt_ae_if :
    issue_slots_12_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_xcpt_ma_if = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_xcpt_ma_if :
    issue_slots_12_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_bp_debug_if = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_bp_debug_if :
    issue_slots_12_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_bp_xcpt_if = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_bp_xcpt_if :
    issue_slots_12_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_debug_fsrc = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_debug_fsrc :
    issue_slots_12_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_11_io_in_uop_bits_debug_tsrc = _GEN_29[1:0] == 2'h2 ? issue_slots_13_out_uop_debug_tsrc :
    issue_slots_12_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_clock = clock;
  assign slots_12_reset = reset;
  assign slots_12_io_grant = issue_slots_12_request & _T_513 & ~_T_507; // @[issue-unit-age-ordered.scala 122:56]
  assign slots_12_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_12_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_12_io_clear = _GEN_27[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_12_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_12_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_12_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_12_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_12_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_12_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_12_io_in_uop_valid = _GEN_31[1:0] == 2'h2 ? issue_slots_14_will_be_valid : _GEN_2390; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_12_io_in_uop_bits_switch = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_switch :
    issue_slots_13_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_switch_off = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_switch_off :
    issue_slots_13_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_unicore = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_is_unicore :
    issue_slots_13_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_shift = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_shift :
    issue_slots_13_out_uop_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_lrs3_rtype = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_lrs3_rtype :
    issue_slots_13_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_rflag = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_rflag :
    issue_slots_13_out_uop_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_wflag = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_wflag :
    issue_slots_13_out_uop_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_prflag = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_prflag :
    issue_slots_13_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_pwflag = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_pwflag :
    issue_slots_13_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_pflag_busy = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_pflag_busy :
    issue_slots_13_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_stale_pflag = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_stale_pflag :
    issue_slots_13_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_op1_sel = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_op1_sel :
    issue_slots_13_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_op2_sel = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_op2_sel :
    issue_slots_13_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_split_num = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_split_num :
    issue_slots_13_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_self_index = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_self_index :
    issue_slots_13_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_rob_inst_idx = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_rob_inst_idx :
    issue_slots_13_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_address_num = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_address_num :
    issue_slots_13_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_uopc = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_uopc : issue_slots_13_out_uop_uopc
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_inst = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_inst : issue_slots_13_out_uop_inst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_debug_inst = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_debug_inst :
    issue_slots_13_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_rvc = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_is_rvc :
    issue_slots_13_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_debug_pc = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_debug_pc :
    issue_slots_13_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_iq_type = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_iq_type :
    issue_slots_13_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_fu_code = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_fu_code :
    issue_slots_13_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_br_type = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_br_type :
    issue_slots_13_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_op1_sel = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_op1_sel :
    issue_slots_13_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_op2_sel = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_op2_sel :
    issue_slots_13_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_imm_sel = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_imm_sel :
    issue_slots_13_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_op_fcn = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_op_fcn :
    issue_slots_13_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_fcn_dw = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_fcn_dw :
    issue_slots_13_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_csr_cmd = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_csr_cmd :
    issue_slots_13_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_is_load = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_is_load :
    issue_slots_13_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_is_sta = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_is_sta :
    issue_slots_13_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_is_std = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_is_std :
    issue_slots_13_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ctrl_op3_sel = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_ctrl_op3_sel :
    issue_slots_13_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_iw_state = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_iw_state :
    issue_slots_13_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_iw_p1_poisoned = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_iw_p1_poisoned :
    issue_slots_13_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_iw_p2_poisoned = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_iw_p2_poisoned :
    issue_slots_13_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_br = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_is_br :
    issue_slots_13_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_jalr = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_is_jalr :
    issue_slots_13_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_jal = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_is_jal :
    issue_slots_13_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_sfb = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_is_sfb :
    issue_slots_13_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_br_mask = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_br_mask :
    issue_slots_13_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_br_tag = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_br_tag :
    issue_slots_13_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ftq_idx = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_ftq_idx :
    issue_slots_13_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_edge_inst = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_edge_inst :
    issue_slots_13_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_pc_lob = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_pc_lob :
    issue_slots_13_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_taken = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_taken :
    issue_slots_13_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_imm_packed = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_imm_packed :
    issue_slots_13_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_csr_addr = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_csr_addr :
    issue_slots_13_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_rob_idx = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_rob_idx :
    issue_slots_13_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ldq_idx = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_ldq_idx :
    issue_slots_13_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_stq_idx = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_stq_idx :
    issue_slots_13_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_rxq_idx = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_rxq_idx :
    issue_slots_13_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_pdst = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_pdst : issue_slots_13_out_uop_pdst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_prs1 = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_prs1 : issue_slots_13_out_uop_prs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_prs2 = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_prs2 : issue_slots_13_out_uop_prs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_prs3 = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_prs3 : issue_slots_13_out_uop_prs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ppred = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_ppred :
    issue_slots_13_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_prs1_busy = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_prs1_busy :
    issue_slots_13_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_prs2_busy = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_prs2_busy :
    issue_slots_13_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_prs3_busy = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_prs3_busy :
    issue_slots_13_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ppred_busy = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_ppred_busy :
    issue_slots_13_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_stale_pdst = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_stale_pdst :
    issue_slots_13_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_exception = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_exception :
    issue_slots_13_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_exc_cause = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_exc_cause :
    issue_slots_13_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_bypassable = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_bypassable :
    issue_slots_13_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_mem_cmd = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_mem_cmd :
    issue_slots_13_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_mem_size = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_mem_size :
    issue_slots_13_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_mem_signed = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_mem_signed :
    issue_slots_13_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_fence = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_is_fence :
    issue_slots_13_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_fencei = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_is_fencei :
    issue_slots_13_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_amo = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_is_amo :
    issue_slots_13_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_uses_ldq = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_uses_ldq :
    issue_slots_13_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_uses_stq = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_uses_stq :
    issue_slots_13_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_sys_pc2epc = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_is_sys_pc2epc :
    issue_slots_13_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_is_unique = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_is_unique :
    issue_slots_13_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_flush_on_commit = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_flush_on_commit :
    issue_slots_13_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ldst_is_rs1 = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_ldst_is_rs1 :
    issue_slots_13_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ldst = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_ldst : issue_slots_13_out_uop_ldst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_lrs1 = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_lrs1 : issue_slots_13_out_uop_lrs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_lrs2 = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_lrs2 : issue_slots_13_out_uop_lrs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_lrs3 = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_lrs3 : issue_slots_13_out_uop_lrs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_ldst_val = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_ldst_val :
    issue_slots_13_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_dst_rtype = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_dst_rtype :
    issue_slots_13_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_lrs1_rtype = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_lrs1_rtype :
    issue_slots_13_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_lrs2_rtype = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_lrs2_rtype :
    issue_slots_13_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_frs3_en = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_frs3_en :
    issue_slots_13_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_fp_val = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_fp_val :
    issue_slots_13_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_fp_single = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_fp_single :
    issue_slots_13_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_xcpt_pf_if = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_xcpt_pf_if :
    issue_slots_13_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_xcpt_ae_if = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_xcpt_ae_if :
    issue_slots_13_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_xcpt_ma_if = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_xcpt_ma_if :
    issue_slots_13_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_bp_debug_if = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_bp_debug_if :
    issue_slots_13_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_bp_xcpt_if = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_bp_xcpt_if :
    issue_slots_13_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_debug_fsrc = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_debug_fsrc :
    issue_slots_13_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_12_io_in_uop_bits_debug_tsrc = _GEN_31[1:0] == 2'h2 ? issue_slots_14_out_uop_debug_tsrc :
    issue_slots_13_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_clock = clock;
  assign slots_13_reset = reset;
  assign slots_13_io_grant = issue_slots_13_request & _T_528 & ~_T_522; // @[issue-unit-age-ordered.scala 122:56]
  assign slots_13_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_13_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_13_io_clear = _GEN_29[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_13_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_13_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_13_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_13_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_13_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_13_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_13_io_in_uop_valid = _GEN_33[1:0] == 2'h2 ? issue_slots_15_will_be_valid : _GEN_2586; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_13_io_in_uop_bits_switch = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_switch :
    issue_slots_14_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_switch_off = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_switch_off :
    issue_slots_14_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_unicore = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_is_unicore :
    issue_slots_14_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_shift = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_shift :
    issue_slots_14_out_uop_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_lrs3_rtype = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_lrs3_rtype :
    issue_slots_14_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_rflag = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_rflag :
    issue_slots_14_out_uop_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_wflag = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_wflag :
    issue_slots_14_out_uop_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_prflag = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_prflag :
    issue_slots_14_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_pwflag = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_pwflag :
    issue_slots_14_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_pflag_busy = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_pflag_busy :
    issue_slots_14_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_stale_pflag = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_stale_pflag :
    issue_slots_14_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_op1_sel = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_op1_sel :
    issue_slots_14_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_op2_sel = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_op2_sel :
    issue_slots_14_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_split_num = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_split_num :
    issue_slots_14_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_self_index = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_self_index :
    issue_slots_14_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_rob_inst_idx = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_rob_inst_idx :
    issue_slots_14_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_address_num = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_address_num :
    issue_slots_14_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_uopc = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_uopc : issue_slots_14_out_uop_uopc
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_inst = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_inst : issue_slots_14_out_uop_inst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_debug_inst = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_debug_inst :
    issue_slots_14_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_rvc = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_is_rvc :
    issue_slots_14_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_debug_pc = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_debug_pc :
    issue_slots_14_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_iq_type = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_iq_type :
    issue_slots_14_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_fu_code = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_fu_code :
    issue_slots_14_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_br_type = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_br_type :
    issue_slots_14_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_op1_sel = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_op1_sel :
    issue_slots_14_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_op2_sel = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_op2_sel :
    issue_slots_14_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_imm_sel = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_imm_sel :
    issue_slots_14_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_op_fcn = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_op_fcn :
    issue_slots_14_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_fcn_dw = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_fcn_dw :
    issue_slots_14_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_csr_cmd = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_csr_cmd :
    issue_slots_14_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_is_load = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_is_load :
    issue_slots_14_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_is_sta = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_is_sta :
    issue_slots_14_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_is_std = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_is_std :
    issue_slots_14_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ctrl_op3_sel = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_ctrl_op3_sel :
    issue_slots_14_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_iw_state = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_iw_state :
    issue_slots_14_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_iw_p1_poisoned = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_iw_p1_poisoned :
    issue_slots_14_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_iw_p2_poisoned = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_iw_p2_poisoned :
    issue_slots_14_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_br = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_is_br :
    issue_slots_14_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_jalr = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_is_jalr :
    issue_slots_14_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_jal = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_is_jal :
    issue_slots_14_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_sfb = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_is_sfb :
    issue_slots_14_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_br_mask = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_br_mask :
    issue_slots_14_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_br_tag = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_br_tag :
    issue_slots_14_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ftq_idx = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_ftq_idx :
    issue_slots_14_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_edge_inst = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_edge_inst :
    issue_slots_14_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_pc_lob = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_pc_lob :
    issue_slots_14_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_taken = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_taken :
    issue_slots_14_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_imm_packed = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_imm_packed :
    issue_slots_14_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_csr_addr = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_csr_addr :
    issue_slots_14_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_rob_idx = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_rob_idx :
    issue_slots_14_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ldq_idx = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_ldq_idx :
    issue_slots_14_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_stq_idx = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_stq_idx :
    issue_slots_14_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_rxq_idx = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_rxq_idx :
    issue_slots_14_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_pdst = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_pdst : issue_slots_14_out_uop_pdst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_prs1 = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_prs1 : issue_slots_14_out_uop_prs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_prs2 = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_prs2 : issue_slots_14_out_uop_prs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_prs3 = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_prs3 : issue_slots_14_out_uop_prs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ppred = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_ppred :
    issue_slots_14_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_prs1_busy = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_prs1_busy :
    issue_slots_14_out_uop_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_prs2_busy = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_prs2_busy :
    issue_slots_14_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_prs3_busy = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_prs3_busy :
    issue_slots_14_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ppred_busy = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_ppred_busy :
    issue_slots_14_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_stale_pdst = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_stale_pdst :
    issue_slots_14_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_exception = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_exception :
    issue_slots_14_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_exc_cause = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_exc_cause :
    issue_slots_14_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_bypassable = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_bypassable :
    issue_slots_14_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_mem_cmd = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_mem_cmd :
    issue_slots_14_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_mem_size = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_mem_size :
    issue_slots_14_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_mem_signed = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_mem_signed :
    issue_slots_14_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_fence = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_is_fence :
    issue_slots_14_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_fencei = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_is_fencei :
    issue_slots_14_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_amo = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_is_amo :
    issue_slots_14_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_uses_ldq = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_uses_ldq :
    issue_slots_14_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_uses_stq = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_uses_stq :
    issue_slots_14_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_sys_pc2epc = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_is_sys_pc2epc :
    issue_slots_14_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_is_unique = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_is_unique :
    issue_slots_14_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_flush_on_commit = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_flush_on_commit :
    issue_slots_14_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ldst_is_rs1 = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_ldst_is_rs1 :
    issue_slots_14_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ldst = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_ldst : issue_slots_14_out_uop_ldst
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_lrs1 = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_lrs1 : issue_slots_14_out_uop_lrs1
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_lrs2 = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_lrs2 : issue_slots_14_out_uop_lrs2
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_lrs3 = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_lrs3 : issue_slots_14_out_uop_lrs3
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_ldst_val = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_ldst_val :
    issue_slots_14_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_dst_rtype = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_dst_rtype :
    issue_slots_14_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_lrs1_rtype = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_lrs1_rtype :
    issue_slots_14_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_lrs2_rtype = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_lrs2_rtype :
    issue_slots_14_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_frs3_en = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_frs3_en :
    issue_slots_14_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_fp_val = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_fp_val :
    issue_slots_14_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_fp_single = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_fp_single :
    issue_slots_14_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_xcpt_pf_if = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_xcpt_pf_if :
    issue_slots_14_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_xcpt_ae_if = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_xcpt_ae_if :
    issue_slots_14_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_xcpt_ma_if = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_xcpt_ma_if :
    issue_slots_14_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_bp_debug_if = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_bp_debug_if :
    issue_slots_14_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_bp_xcpt_if = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_bp_xcpt_if :
    issue_slots_14_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_debug_fsrc = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_debug_fsrc :
    issue_slots_14_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_13_io_in_uop_bits_debug_tsrc = _GEN_33[1:0] == 2'h2 ? issue_slots_15_out_uop_debug_tsrc :
    issue_slots_14_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_clock = clock;
  assign slots_14_reset = reset;
  assign slots_14_io_grant = issue_slots_14_request & _T_543 & ~_T_537; // @[issue-unit-age-ordered.scala 122:56]
  assign slots_14_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_14_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_14_io_clear = _GEN_31[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_14_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_14_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_14_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_14_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_14_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_14_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_14_io_in_uop_valid = _GEN_35[1:0] == 2'h2 ? will_be_valid_16 : _GEN_2782; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_14_io_in_uop_bits_switch = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_switch :
    issue_slots_15_out_uop_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_switch_off = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_switch_off :
    issue_slots_15_out_uop_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_unicore = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_is_unicore :
    issue_slots_15_out_uop_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_shift = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_shift : issue_slots_15_out_uop_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_lrs3_rtype = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_lrs3_rtype :
    issue_slots_15_out_uop_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_rflag = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_rflag : issue_slots_15_out_uop_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_wflag = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_wflag : issue_slots_15_out_uop_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_prflag = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_prflag :
    issue_slots_15_out_uop_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_pwflag = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_pwflag :
    issue_slots_15_out_uop_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_pflag_busy = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_pflag_busy :
    issue_slots_15_out_uop_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_stale_pflag = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_stale_pflag :
    issue_slots_15_out_uop_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_op1_sel = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_op1_sel :
    issue_slots_15_out_uop_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_op2_sel = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_op2_sel :
    issue_slots_15_out_uop_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_split_num = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_split_num :
    issue_slots_15_out_uop_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_self_index = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_self_index :
    issue_slots_15_out_uop_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_rob_inst_idx = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_rob_inst_idx :
    issue_slots_15_out_uop_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_address_num = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_address_num :
    issue_slots_15_out_uop_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_uopc = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_uopc : issue_slots_15_out_uop_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_inst = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_inst : issue_slots_15_out_uop_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_debug_inst = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_debug_inst :
    issue_slots_15_out_uop_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_rvc = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_is_rvc :
    issue_slots_15_out_uop_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_debug_pc = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_debug_pc :
    issue_slots_15_out_uop_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_iq_type = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_iq_type :
    issue_slots_15_out_uop_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_fu_code = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_fu_code :
    issue_slots_15_out_uop_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_br_type = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_br_type :
    issue_slots_15_out_uop_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_op1_sel = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_op1_sel :
    issue_slots_15_out_uop_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_op2_sel = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_op2_sel :
    issue_slots_15_out_uop_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_imm_sel = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_imm_sel :
    issue_slots_15_out_uop_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_op_fcn = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_op_fcn :
    issue_slots_15_out_uop_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_fcn_dw = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_fcn_dw :
    issue_slots_15_out_uop_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_csr_cmd = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_csr_cmd :
    issue_slots_15_out_uop_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_is_load = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_is_load :
    issue_slots_15_out_uop_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_is_sta = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_is_sta :
    issue_slots_15_out_uop_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_is_std = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_is_std :
    issue_slots_15_out_uop_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ctrl_op3_sel = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_ctrl_op3_sel :
    issue_slots_15_out_uop_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_iw_state = _GEN_35[1:0] == 2'h2 ? 2'h1 : issue_slots_15_out_uop_iw_state; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_iw_p1_poisoned = _GEN_35[1:0] == 2'h2 ? 1'h0 : issue_slots_15_out_uop_iw_p1_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_iw_p2_poisoned = _GEN_35[1:0] == 2'h2 ? 1'h0 : issue_slots_15_out_uop_iw_p2_poisoned; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_br = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_is_br : issue_slots_15_out_uop_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_jalr = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_is_jalr :
    issue_slots_15_out_uop_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_jal = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_is_jal :
    issue_slots_15_out_uop_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_sfb = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_is_sfb :
    issue_slots_15_out_uop_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_br_mask = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_br_mask :
    issue_slots_15_out_uop_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_br_tag = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_br_tag :
    issue_slots_15_out_uop_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ftq_idx = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_ftq_idx :
    issue_slots_15_out_uop_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_edge_inst = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_edge_inst :
    issue_slots_15_out_uop_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_pc_lob = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_pc_lob :
    issue_slots_15_out_uop_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_taken = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_taken : issue_slots_15_out_uop_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_imm_packed = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_imm_packed :
    issue_slots_15_out_uop_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_csr_addr = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_csr_addr :
    issue_slots_15_out_uop_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_rob_idx = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_rob_idx :
    issue_slots_15_out_uop_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ldq_idx = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_ldq_idx :
    issue_slots_15_out_uop_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_stq_idx = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_stq_idx :
    issue_slots_15_out_uop_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_rxq_idx = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_rxq_idx :
    issue_slots_15_out_uop_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_pdst = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_pdst : issue_slots_15_out_uop_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_prs1 = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_prs1 : issue_slots_15_out_uop_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_prs2 = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_prs2 : issue_slots_15_out_uop_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_prs3 = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_prs3 : issue_slots_15_out_uop_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ppred = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_ppred : issue_slots_15_out_uop_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_prs1_busy = _GEN_35[1:0] == 2'h2 ? uops_16_prs1_busy : issue_slots_15_out_uop_prs1_busy
    ; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_prs2_busy = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_prs2_busy :
    issue_slots_15_out_uop_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_prs3_busy = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_prs3_busy :
    issue_slots_15_out_uop_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ppred_busy = _GEN_35[1:0] == 2'h2 ? 1'h0 : issue_slots_15_out_uop_ppred_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_stale_pdst = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_stale_pdst :
    issue_slots_15_out_uop_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_exception = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_exception :
    issue_slots_15_out_uop_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_exc_cause = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_exc_cause :
    issue_slots_15_out_uop_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_bypassable = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_bypassable :
    issue_slots_15_out_uop_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_mem_cmd = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_mem_cmd :
    issue_slots_15_out_uop_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_mem_size = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_mem_size :
    issue_slots_15_out_uop_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_mem_signed = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_mem_signed :
    issue_slots_15_out_uop_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_fence = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_is_fence :
    issue_slots_15_out_uop_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_fencei = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_is_fencei :
    issue_slots_15_out_uop_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_amo = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_is_amo :
    issue_slots_15_out_uop_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_uses_ldq = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_uses_ldq :
    issue_slots_15_out_uop_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_uses_stq = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_uses_stq :
    issue_slots_15_out_uop_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_sys_pc2epc = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_is_sys_pc2epc :
    issue_slots_15_out_uop_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_is_unique = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_is_unique :
    issue_slots_15_out_uop_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_flush_on_commit = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_flush_on_commit :
    issue_slots_15_out_uop_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ldst_is_rs1 = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_ldst_is_rs1 :
    issue_slots_15_out_uop_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ldst = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_ldst : issue_slots_15_out_uop_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_lrs1 = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_lrs1 : issue_slots_15_out_uop_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_lrs2 = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_lrs2 : issue_slots_15_out_uop_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_lrs3 = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_lrs3 : issue_slots_15_out_uop_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_ldst_val = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_ldst_val :
    issue_slots_15_out_uop_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_dst_rtype = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_dst_rtype :
    issue_slots_15_out_uop_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_lrs1_rtype = _GEN_35[1:0] == 2'h2 ? uops_16_lrs1_rtype :
    issue_slots_15_out_uop_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_lrs2_rtype = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_lrs2_rtype :
    issue_slots_15_out_uop_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_frs3_en = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_frs3_en :
    issue_slots_15_out_uop_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_fp_val = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_fp_val :
    issue_slots_15_out_uop_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_fp_single = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_fp_single :
    issue_slots_15_out_uop_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_xcpt_pf_if = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_xcpt_pf_if :
    issue_slots_15_out_uop_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_xcpt_ae_if = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_xcpt_ae_if :
    issue_slots_15_out_uop_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_xcpt_ma_if = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_xcpt_ma_if :
    issue_slots_15_out_uop_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_bp_debug_if = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_bp_debug_if :
    issue_slots_15_out_uop_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_bp_xcpt_if = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_bp_xcpt_if :
    issue_slots_15_out_uop_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_debug_fsrc = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_debug_fsrc :
    issue_slots_15_out_uop_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_14_io_in_uop_bits_debug_tsrc = _GEN_35[1:0] == 2'h2 ? io_dis_uops_0_bits_debug_tsrc :
    issue_slots_15_out_uop_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_clock = clock;
  assign slots_15_reset = reset;
  assign slots_15_io_grant = issue_slots_15_request & _T_558 & ~_T_552; // @[issue-unit-age-ordered.scala 122:56]
  assign slots_15_io_brupdate_b1_resolve_mask = io_brupdate_b1_resolve_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b1_mispredict_mask = io_brupdate_b1_mispredict_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_switch = io_brupdate_b2_uop_switch; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_switch_off = io_brupdate_b2_uop_switch_off; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_unicore = io_brupdate_b2_uop_is_unicore; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_shift = io_brupdate_b2_uop_shift; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_lrs3_rtype = io_brupdate_b2_uop_lrs3_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_rflag = io_brupdate_b2_uop_rflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_wflag = io_brupdate_b2_uop_wflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_prflag = io_brupdate_b2_uop_prflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_pwflag = io_brupdate_b2_uop_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_pflag_busy = io_brupdate_b2_uop_pflag_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_stale_pflag = io_brupdate_b2_uop_stale_pflag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_op1_sel = io_brupdate_b2_uop_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_op2_sel = io_brupdate_b2_uop_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_split_num = io_brupdate_b2_uop_split_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_self_index = io_brupdate_b2_uop_self_index; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_rob_inst_idx = io_brupdate_b2_uop_rob_inst_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_address_num = io_brupdate_b2_uop_address_num; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_uopc = io_brupdate_b2_uop_uopc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_inst = io_brupdate_b2_uop_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_debug_inst = io_brupdate_b2_uop_debug_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_rvc = io_brupdate_b2_uop_is_rvc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_debug_pc = io_brupdate_b2_uop_debug_pc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_iq_type = io_brupdate_b2_uop_iq_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_fu_code = io_brupdate_b2_uop_fu_code; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_br_type = io_brupdate_b2_uop_ctrl_br_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_op1_sel = io_brupdate_b2_uop_ctrl_op1_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_op2_sel = io_brupdate_b2_uop_ctrl_op2_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_imm_sel = io_brupdate_b2_uop_ctrl_imm_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_op_fcn = io_brupdate_b2_uop_ctrl_op_fcn; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_fcn_dw = io_brupdate_b2_uop_ctrl_fcn_dw; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_csr_cmd = io_brupdate_b2_uop_ctrl_csr_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_is_load = io_brupdate_b2_uop_ctrl_is_load; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_is_sta = io_brupdate_b2_uop_ctrl_is_sta; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_is_std = io_brupdate_b2_uop_ctrl_is_std; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ctrl_op3_sel = io_brupdate_b2_uop_ctrl_op3_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_iw_state = io_brupdate_b2_uop_iw_state; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_iw_p1_poisoned = io_brupdate_b2_uop_iw_p1_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_iw_p2_poisoned = io_brupdate_b2_uop_iw_p2_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_br = io_brupdate_b2_uop_is_br; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_jalr = io_brupdate_b2_uop_is_jalr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_jal = io_brupdate_b2_uop_is_jal; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_sfb = io_brupdate_b2_uop_is_sfb; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_br_mask = io_brupdate_b2_uop_br_mask; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_br_tag = io_brupdate_b2_uop_br_tag; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ftq_idx = io_brupdate_b2_uop_ftq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_edge_inst = io_brupdate_b2_uop_edge_inst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_pc_lob = io_brupdate_b2_uop_pc_lob; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_taken = io_brupdate_b2_uop_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_imm_packed = io_brupdate_b2_uop_imm_packed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_csr_addr = io_brupdate_b2_uop_csr_addr; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_rob_idx = io_brupdate_b2_uop_rob_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ldq_idx = io_brupdate_b2_uop_ldq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_stq_idx = io_brupdate_b2_uop_stq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_rxq_idx = io_brupdate_b2_uop_rxq_idx; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_pdst = io_brupdate_b2_uop_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_prs1 = io_brupdate_b2_uop_prs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_prs2 = io_brupdate_b2_uop_prs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_prs3 = io_brupdate_b2_uop_prs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ppred = io_brupdate_b2_uop_ppred; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_prs1_busy = io_brupdate_b2_uop_prs1_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_prs2_busy = io_brupdate_b2_uop_prs2_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_prs3_busy = io_brupdate_b2_uop_prs3_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ppred_busy = io_brupdate_b2_uop_ppred_busy; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_stale_pdst = io_brupdate_b2_uop_stale_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_exception = io_brupdate_b2_uop_exception; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_exc_cause = io_brupdate_b2_uop_exc_cause; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_bypassable = io_brupdate_b2_uop_bypassable; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_mem_cmd = io_brupdate_b2_uop_mem_cmd; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_mem_size = io_brupdate_b2_uop_mem_size; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_mem_signed = io_brupdate_b2_uop_mem_signed; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_fence = io_brupdate_b2_uop_is_fence; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_fencei = io_brupdate_b2_uop_is_fencei; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_amo = io_brupdate_b2_uop_is_amo; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_uses_ldq = io_brupdate_b2_uop_uses_ldq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_uses_stq = io_brupdate_b2_uop_uses_stq; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_sys_pc2epc = io_brupdate_b2_uop_is_sys_pc2epc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_is_unique = io_brupdate_b2_uop_is_unique; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_flush_on_commit = io_brupdate_b2_uop_flush_on_commit; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ldst_is_rs1 = io_brupdate_b2_uop_ldst_is_rs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ldst = io_brupdate_b2_uop_ldst; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_lrs1 = io_brupdate_b2_uop_lrs1; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_lrs2 = io_brupdate_b2_uop_lrs2; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_lrs3 = io_brupdate_b2_uop_lrs3; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_ldst_val = io_brupdate_b2_uop_ldst_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_dst_rtype = io_brupdate_b2_uop_dst_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_lrs1_rtype = io_brupdate_b2_uop_lrs1_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_lrs2_rtype = io_brupdate_b2_uop_lrs2_rtype; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_frs3_en = io_brupdate_b2_uop_frs3_en; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_fp_val = io_brupdate_b2_uop_fp_val; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_fp_single = io_brupdate_b2_uop_fp_single; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_xcpt_pf_if = io_brupdate_b2_uop_xcpt_pf_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_xcpt_ae_if = io_brupdate_b2_uop_xcpt_ae_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_xcpt_ma_if = io_brupdate_b2_uop_xcpt_ma_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_bp_debug_if = io_brupdate_b2_uop_bp_debug_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_bp_xcpt_if = io_brupdate_b2_uop_bp_xcpt_if; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_debug_fsrc = io_brupdate_b2_uop_debug_fsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_uop_debug_tsrc = io_brupdate_b2_uop_debug_tsrc; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_valid = io_brupdate_b2_valid; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_mispredict = io_brupdate_b2_mispredict; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_taken = io_brupdate_b2_taken; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_cfi_type = io_brupdate_b2_cfi_type; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_pc_sel = io_brupdate_b2_pc_sel; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_jalr_target = io_brupdate_b2_jalr_target; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_brupdate_b2_target_offset = io_brupdate_b2_target_offset; // @[issue-unit.scala 158:28 issue-unit.scala 165:37]
  assign slots_15_io_kill = io_flush_pipeline; // @[issue-unit.scala 158:28 issue-unit.scala 166:37]
  assign slots_15_io_clear = _GEN_33[1:0] != 2'h0; // @[issue-unit-age-ordered.scala 76:49]
  assign slots_15_io_ldspec_miss = io_ld_miss; // @[issue-unit.scala 158:28 issue-unit.scala 164:37]
  assign slots_15_io_wakeup_ports_0_valid = io_wakeup_ports_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_0_bits_pdst = io_wakeup_ports_0_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_0_bits_poisoned = io_wakeup_ports_0_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_0_bits_pwflag = io_wakeup_ports_0_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_0_bits_flag_valid = io_wakeup_ports_0_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_1_valid = io_wakeup_ports_1_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_1_bits_pdst = io_wakeup_ports_1_bits_pdst; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_1_bits_poisoned = io_wakeup_ports_1_bits_poisoned; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_1_bits_pwflag = io_wakeup_ports_1_bits_pwflag; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_wakeup_ports_1_bits_flag_valid = io_wakeup_ports_1_bits_flag_valid; // @[issue-unit.scala 158:28 issue-unit.scala 161:37]
  assign slots_15_io_pred_wakeup_port_valid = io_pred_wakeup_port_valid; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_15_io_pred_wakeup_port_bits = io_pred_wakeup_port_bits; // @[issue-unit.scala 158:28 issue-unit.scala 162:37]
  assign slots_15_io_spec_ld_wakeup_0_valid = io_spec_ld_wakeup_0_valid; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_15_io_spec_ld_wakeup_0_bits = io_spec_ld_wakeup_0_bits; // @[issue-unit.scala 158:28 issue-unit.scala 163:37]
  assign slots_15_io_in_uop_valid = _GEN_37[1:0] == 2'h2 ? will_be_valid_17 : _GEN_2978; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 72:37]
  assign slots_15_io_in_uop_bits_switch = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_switch : io_dis_uops_0_bits_switch; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_switch_off = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_switch_off :
    io_dis_uops_0_bits_switch_off; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_unicore = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_is_unicore :
    io_dis_uops_0_bits_is_unicore; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_shift = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_shift : io_dis_uops_0_bits_shift; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_lrs3_rtype = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_lrs3_rtype :
    io_dis_uops_0_bits_lrs3_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_rflag = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_rflag : io_dis_uops_0_bits_rflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_wflag = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_wflag : io_dis_uops_0_bits_wflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_prflag = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_prflag : io_dis_uops_0_bits_prflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_pwflag = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_pwflag : io_dis_uops_0_bits_pwflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_pflag_busy = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_pflag_busy :
    io_dis_uops_0_bits_pflag_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_stale_pflag = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_stale_pflag :
    io_dis_uops_0_bits_stale_pflag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_op1_sel = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_op1_sel :
    io_dis_uops_0_bits_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_op2_sel = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_op2_sel :
    io_dis_uops_0_bits_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_split_num = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_split_num :
    io_dis_uops_0_bits_split_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_self_index = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_self_index :
    io_dis_uops_0_bits_self_index; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_rob_inst_idx = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_rob_inst_idx :
    io_dis_uops_0_bits_rob_inst_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_address_num = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_address_num :
    io_dis_uops_0_bits_address_num; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_uopc = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_uopc : io_dis_uops_0_bits_uopc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_inst = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_inst : io_dis_uops_0_bits_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_debug_inst = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_debug_inst :
    io_dis_uops_0_bits_debug_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_rvc = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_is_rvc : io_dis_uops_0_bits_is_rvc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_debug_pc = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_debug_pc :
    io_dis_uops_0_bits_debug_pc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_iq_type = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_iq_type :
    io_dis_uops_0_bits_iq_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_fu_code = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_fu_code :
    io_dis_uops_0_bits_fu_code; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_br_type = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_br_type :
    io_dis_uops_0_bits_ctrl_br_type; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_op1_sel = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_op1_sel :
    io_dis_uops_0_bits_ctrl_op1_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_op2_sel = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_op2_sel :
    io_dis_uops_0_bits_ctrl_op2_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_imm_sel = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_imm_sel :
    io_dis_uops_0_bits_ctrl_imm_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_op_fcn = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_op_fcn :
    io_dis_uops_0_bits_ctrl_op_fcn; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_fcn_dw = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_fcn_dw :
    io_dis_uops_0_bits_ctrl_fcn_dw; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_csr_cmd = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_csr_cmd :
    io_dis_uops_0_bits_ctrl_csr_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_is_load = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_is_load :
    io_dis_uops_0_bits_ctrl_is_load; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_is_sta = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_is_sta :
    io_dis_uops_0_bits_ctrl_is_sta; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_is_std = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_is_std :
    io_dis_uops_0_bits_ctrl_is_std; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ctrl_op3_sel = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_ctrl_op3_sel :
    io_dis_uops_0_bits_ctrl_op3_sel; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_iw_state = 2'h1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_iw_p1_poisoned = 1'h0; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_iw_p2_poisoned = 1'h0; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_br = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_is_br : io_dis_uops_0_bits_is_br; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_jalr = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_is_jalr :
    io_dis_uops_0_bits_is_jalr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_jal = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_is_jal : io_dis_uops_0_bits_is_jal; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_sfb = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_is_sfb : io_dis_uops_0_bits_is_sfb; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_br_mask = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_br_mask :
    io_dis_uops_0_bits_br_mask; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_br_tag = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_br_tag : io_dis_uops_0_bits_br_tag; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ftq_idx = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_ftq_idx :
    io_dis_uops_0_bits_ftq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_edge_inst = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_edge_inst :
    io_dis_uops_0_bits_edge_inst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_pc_lob = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_pc_lob : io_dis_uops_0_bits_pc_lob; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_taken = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_taken : io_dis_uops_0_bits_taken; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_imm_packed = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_imm_packed :
    io_dis_uops_0_bits_imm_packed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_csr_addr = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_csr_addr :
    io_dis_uops_0_bits_csr_addr; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_rob_idx = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_rob_idx :
    io_dis_uops_0_bits_rob_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ldq_idx = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_ldq_idx :
    io_dis_uops_0_bits_ldq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_stq_idx = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_stq_idx :
    io_dis_uops_0_bits_stq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_rxq_idx = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_rxq_idx :
    io_dis_uops_0_bits_rxq_idx; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_pdst = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_pdst : io_dis_uops_0_bits_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_prs1 = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_prs1 : io_dis_uops_0_bits_prs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_prs2 = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_prs2 : io_dis_uops_0_bits_prs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_prs3 = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_prs3 : io_dis_uops_0_bits_prs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ppred = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_ppred : io_dis_uops_0_bits_ppred; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_prs1_busy = _GEN_37[1:0] == 2'h2 ? uops_17_prs1_busy : uops_16_prs1_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_prs2_busy = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_prs2_busy :
    io_dis_uops_0_bits_prs2_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_prs3_busy = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_prs3_busy :
    io_dis_uops_0_bits_prs3_busy; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ppred_busy = 1'h0; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_stale_pdst = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_stale_pdst :
    io_dis_uops_0_bits_stale_pdst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_exception = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_exception :
    io_dis_uops_0_bits_exception; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_exc_cause = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_exc_cause :
    io_dis_uops_0_bits_exc_cause; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_bypassable = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_bypassable :
    io_dis_uops_0_bits_bypassable; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_mem_cmd = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_mem_cmd :
    io_dis_uops_0_bits_mem_cmd; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_mem_size = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_mem_size :
    io_dis_uops_0_bits_mem_size; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_mem_signed = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_mem_signed :
    io_dis_uops_0_bits_mem_signed; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_fence = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_is_fence :
    io_dis_uops_0_bits_is_fence; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_fencei = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_is_fencei :
    io_dis_uops_0_bits_is_fencei; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_amo = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_is_amo : io_dis_uops_0_bits_is_amo; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_uses_ldq = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_uses_ldq :
    io_dis_uops_0_bits_uses_ldq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_uses_stq = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_uses_stq :
    io_dis_uops_0_bits_uses_stq; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_sys_pc2epc = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_is_sys_pc2epc :
    io_dis_uops_0_bits_is_sys_pc2epc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_is_unique = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_is_unique :
    io_dis_uops_0_bits_is_unique; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_flush_on_commit = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_flush_on_commit :
    io_dis_uops_0_bits_flush_on_commit; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ldst_is_rs1 = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_ldst_is_rs1 :
    io_dis_uops_0_bits_ldst_is_rs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ldst = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_ldst : io_dis_uops_0_bits_ldst; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_lrs1 = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_lrs1 : io_dis_uops_0_bits_lrs1; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_lrs2 = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_lrs2 : io_dis_uops_0_bits_lrs2; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_lrs3 = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_lrs3 : io_dis_uops_0_bits_lrs3; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_ldst_val = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_ldst_val :
    io_dis_uops_0_bits_ldst_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_dst_rtype = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_dst_rtype :
    io_dis_uops_0_bits_dst_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_lrs1_rtype = _GEN_37[1:0] == 2'h2 ? uops_17_lrs1_rtype : uops_16_lrs1_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_lrs2_rtype = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_lrs2_rtype :
    io_dis_uops_0_bits_lrs2_rtype; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_frs3_en = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_frs3_en :
    io_dis_uops_0_bits_frs3_en; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_fp_val = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_fp_val : io_dis_uops_0_bits_fp_val; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_fp_single = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_fp_single :
    io_dis_uops_0_bits_fp_single; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_xcpt_pf_if = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_xcpt_pf_if :
    io_dis_uops_0_bits_xcpt_pf_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_xcpt_ae_if = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_xcpt_ae_if :
    io_dis_uops_0_bits_xcpt_ae_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_xcpt_ma_if = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_xcpt_ma_if :
    io_dis_uops_0_bits_xcpt_ma_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_bp_debug_if = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_bp_debug_if :
    io_dis_uops_0_bits_bp_debug_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_bp_xcpt_if = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_bp_xcpt_if :
    io_dis_uops_0_bits_bp_xcpt_if; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_debug_fsrc = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_debug_fsrc :
    io_dis_uops_0_bits_debug_fsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  assign slots_15_io_in_uop_bits_debug_tsrc = _GEN_37[1:0] == 2'h2 ? io_dis_uops_1_bits_debug_tsrc :
    io_dis_uops_0_bits_debug_tsrc; // @[issue-unit-age-ordered.scala 71:48 issue-unit-age-ordered.scala 73:37]
  always @(posedge clock) begin
    REG <= num_available > 5'h0; // @[issue-unit-age-ordered.scala 87:51]
    REG_1 <= num_available > 5'h1; // @[issue-unit-age-ordered.scala 87:51]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_dis_uops_0_bits_ppred_busy & io_dis_uops_0_valid) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at issue-unit.scala:149 assert(!(io.dis_uops(w).bits.ppred_busy && io.dis_uops(w).valid))\n"
            ); // @[issue-unit.scala 149:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_dis_uops_0_bits_ppred_busy & io_dis_uops_0_valid) | reset)) begin
          $fatal; // @[issue-unit.scala 149:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_dis_uops_1_bits_ppred_busy & io_dis_uops_1_valid) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at issue-unit.scala:149 assert(!(io.dis_uops(w).bits.ppred_busy && io.dis_uops(w).valid))\n"
            ); // @[issue-unit.scala 149:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_dis_uops_1_bits_ppred_busy & io_dis_uops_1_valid) | reset)) begin
          $fatal; // @[issue-unit.scala 149:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(_T_85 <= 5'h1 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: [issue] window giving out too many grants.\n    at issue-unit.scala:176 assert (PopCount(issue_slots.map(s => s.grant)) <= issueWidth.U, \"[issue] window giving out too many grants.\")\n"
            ); // @[issue-unit.scala 176:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(_T_85 <= 5'h1 | reset)) begin
          $fatal; // @[issue-unit.scala 176:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG_1 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
