module EnqTranBuff(
  input         clock,
  input         reset,
  input         io_enq_0_dec_uops_0_switch,
  input         io_enq_0_dec_uops_0_switch_off,
  input         io_enq_0_dec_uops_0_is_unicore,
  input  [2:0]  io_enq_0_dec_uops_0_shift,
  input  [1:0]  io_enq_0_dec_uops_0_lrs3_rtype,
  input         io_enq_0_dec_uops_0_rflag,
  input         io_enq_0_dec_uops_0_wflag,
  input  [3:0]  io_enq_0_dec_uops_0_prflag,
  input  [3:0]  io_enq_0_dec_uops_0_pwflag,
  input         io_enq_0_dec_uops_0_pflag_busy,
  input  [3:0]  io_enq_0_dec_uops_0_stale_pflag,
  input  [3:0]  io_enq_0_dec_uops_0_op1_sel,
  input  [3:0]  io_enq_0_dec_uops_0_op2_sel,
  input  [5:0]  io_enq_0_dec_uops_0_split_num,
  input  [5:0]  io_enq_0_dec_uops_0_self_index,
  input  [5:0]  io_enq_0_dec_uops_0_rob_inst_idx,
  input  [5:0]  io_enq_0_dec_uops_0_address_num,
  input  [6:0]  io_enq_0_dec_uops_0_uopc,
  input  [31:0] io_enq_0_dec_uops_0_inst,
  input  [31:0] io_enq_0_dec_uops_0_debug_inst,
  input         io_enq_0_dec_uops_0_is_rvc,
  input  [39:0] io_enq_0_dec_uops_0_debug_pc,
  input  [2:0]  io_enq_0_dec_uops_0_iq_type,
  input  [9:0]  io_enq_0_dec_uops_0_fu_code,
  input  [3:0]  io_enq_0_dec_uops_0_ctrl_br_type,
  input  [1:0]  io_enq_0_dec_uops_0_ctrl_op1_sel,
  input  [2:0]  io_enq_0_dec_uops_0_ctrl_op2_sel,
  input  [2:0]  io_enq_0_dec_uops_0_ctrl_imm_sel,
  input  [3:0]  io_enq_0_dec_uops_0_ctrl_op_fcn,
  input         io_enq_0_dec_uops_0_ctrl_fcn_dw,
  input  [2:0]  io_enq_0_dec_uops_0_ctrl_csr_cmd,
  input         io_enq_0_dec_uops_0_ctrl_is_load,
  input         io_enq_0_dec_uops_0_ctrl_is_sta,
  input         io_enq_0_dec_uops_0_ctrl_is_std,
  input  [1:0]  io_enq_0_dec_uops_0_ctrl_op3_sel,
  input  [1:0]  io_enq_0_dec_uops_0_iw_state,
  input         io_enq_0_dec_uops_0_iw_p1_poisoned,
  input         io_enq_0_dec_uops_0_iw_p2_poisoned,
  input         io_enq_0_dec_uops_0_is_br,
  input         io_enq_0_dec_uops_0_is_jalr,
  input         io_enq_0_dec_uops_0_is_jal,
  input         io_enq_0_dec_uops_0_is_sfb,
  input  [11:0] io_enq_0_dec_uops_0_br_mask,
  input  [3:0]  io_enq_0_dec_uops_0_br_tag,
  input  [4:0]  io_enq_0_dec_uops_0_ftq_idx,
  input         io_enq_0_dec_uops_0_edge_inst,
  input  [5:0]  io_enq_0_dec_uops_0_pc_lob,
  input         io_enq_0_dec_uops_0_taken,
  input  [19:0] io_enq_0_dec_uops_0_imm_packed,
  input  [11:0] io_enq_0_dec_uops_0_csr_addr,
  input  [5:0]  io_enq_0_dec_uops_0_rob_idx,
  input  [4:0]  io_enq_0_dec_uops_0_ldq_idx,
  input  [4:0]  io_enq_0_dec_uops_0_stq_idx,
  input  [1:0]  io_enq_0_dec_uops_0_rxq_idx,
  input  [6:0]  io_enq_0_dec_uops_0_pdst,
  input  [6:0]  io_enq_0_dec_uops_0_prs1,
  input  [6:0]  io_enq_0_dec_uops_0_prs2,
  input  [6:0]  io_enq_0_dec_uops_0_prs3,
  input  [4:0]  io_enq_0_dec_uops_0_ppred,
  input         io_enq_0_dec_uops_0_prs1_busy,
  input         io_enq_0_dec_uops_0_prs2_busy,
  input         io_enq_0_dec_uops_0_prs3_busy,
  input         io_enq_0_dec_uops_0_ppred_busy,
  input  [6:0]  io_enq_0_dec_uops_0_stale_pdst,
  input         io_enq_0_dec_uops_0_exception,
  input  [63:0] io_enq_0_dec_uops_0_exc_cause,
  input         io_enq_0_dec_uops_0_bypassable,
  input  [4:0]  io_enq_0_dec_uops_0_mem_cmd,
  input  [1:0]  io_enq_0_dec_uops_0_mem_size,
  input         io_enq_0_dec_uops_0_mem_signed,
  input         io_enq_0_dec_uops_0_is_fence,
  input         io_enq_0_dec_uops_0_is_fencei,
  input         io_enq_0_dec_uops_0_is_amo,
  input         io_enq_0_dec_uops_0_uses_ldq,
  input         io_enq_0_dec_uops_0_uses_stq,
  input         io_enq_0_dec_uops_0_is_sys_pc2epc,
  input         io_enq_0_dec_uops_0_is_unique,
  input         io_enq_0_dec_uops_0_flush_on_commit,
  input         io_enq_0_dec_uops_0_ldst_is_rs1,
  input  [5:0]  io_enq_0_dec_uops_0_ldst,
  input  [5:0]  io_enq_0_dec_uops_0_lrs1,
  input  [5:0]  io_enq_0_dec_uops_0_lrs2,
  input  [5:0]  io_enq_0_dec_uops_0_lrs3,
  input         io_enq_0_dec_uops_0_ldst_val,
  input  [1:0]  io_enq_0_dec_uops_0_dst_rtype,
  input  [1:0]  io_enq_0_dec_uops_0_lrs1_rtype,
  input  [1:0]  io_enq_0_dec_uops_0_lrs2_rtype,
  input         io_enq_0_dec_uops_0_frs3_en,
  input         io_enq_0_dec_uops_0_fp_val,
  input         io_enq_0_dec_uops_0_fp_single,
  input         io_enq_0_dec_uops_0_xcpt_pf_if,
  input         io_enq_0_dec_uops_0_xcpt_ae_if,
  input         io_enq_0_dec_uops_0_xcpt_ma_if,
  input         io_enq_0_dec_uops_0_bp_debug_if,
  input         io_enq_0_dec_uops_0_bp_xcpt_if,
  input  [1:0]  io_enq_0_dec_uops_0_debug_fsrc,
  input  [1:0]  io_enq_0_dec_uops_0_debug_tsrc,
  input         io_enq_0_dec_uops_1_switch,
  input         io_enq_0_dec_uops_1_switch_off,
  input         io_enq_0_dec_uops_1_is_unicore,
  input  [2:0]  io_enq_0_dec_uops_1_shift,
  input  [1:0]  io_enq_0_dec_uops_1_lrs3_rtype,
  input         io_enq_0_dec_uops_1_rflag,
  input         io_enq_0_dec_uops_1_wflag,
  input  [3:0]  io_enq_0_dec_uops_1_prflag,
  input  [3:0]  io_enq_0_dec_uops_1_pwflag,
  input         io_enq_0_dec_uops_1_pflag_busy,
  input  [3:0]  io_enq_0_dec_uops_1_stale_pflag,
  input  [3:0]  io_enq_0_dec_uops_1_op1_sel,
  input  [3:0]  io_enq_0_dec_uops_1_op2_sel,
  input  [5:0]  io_enq_0_dec_uops_1_split_num,
  input  [5:0]  io_enq_0_dec_uops_1_self_index,
  input  [5:0]  io_enq_0_dec_uops_1_rob_inst_idx,
  input  [5:0]  io_enq_0_dec_uops_1_address_num,
  input  [6:0]  io_enq_0_dec_uops_1_uopc,
  input  [31:0] io_enq_0_dec_uops_1_inst,
  input  [31:0] io_enq_0_dec_uops_1_debug_inst,
  input         io_enq_0_dec_uops_1_is_rvc,
  input  [39:0] io_enq_0_dec_uops_1_debug_pc,
  input  [2:0]  io_enq_0_dec_uops_1_iq_type,
  input  [9:0]  io_enq_0_dec_uops_1_fu_code,
  input  [3:0]  io_enq_0_dec_uops_1_ctrl_br_type,
  input  [1:0]  io_enq_0_dec_uops_1_ctrl_op1_sel,
  input  [2:0]  io_enq_0_dec_uops_1_ctrl_op2_sel,
  input  [2:0]  io_enq_0_dec_uops_1_ctrl_imm_sel,
  input  [3:0]  io_enq_0_dec_uops_1_ctrl_op_fcn,
  input         io_enq_0_dec_uops_1_ctrl_fcn_dw,
  input  [2:0]  io_enq_0_dec_uops_1_ctrl_csr_cmd,
  input         io_enq_0_dec_uops_1_ctrl_is_load,
  input         io_enq_0_dec_uops_1_ctrl_is_sta,
  input         io_enq_0_dec_uops_1_ctrl_is_std,
  input  [1:0]  io_enq_0_dec_uops_1_ctrl_op3_sel,
  input  [1:0]  io_enq_0_dec_uops_1_iw_state,
  input         io_enq_0_dec_uops_1_iw_p1_poisoned,
  input         io_enq_0_dec_uops_1_iw_p2_poisoned,
  input         io_enq_0_dec_uops_1_is_br,
  input         io_enq_0_dec_uops_1_is_jalr,
  input         io_enq_0_dec_uops_1_is_jal,
  input         io_enq_0_dec_uops_1_is_sfb,
  input  [11:0] io_enq_0_dec_uops_1_br_mask,
  input  [3:0]  io_enq_0_dec_uops_1_br_tag,
  input  [4:0]  io_enq_0_dec_uops_1_ftq_idx,
  input         io_enq_0_dec_uops_1_edge_inst,
  input  [5:0]  io_enq_0_dec_uops_1_pc_lob,
  input         io_enq_0_dec_uops_1_taken,
  input  [19:0] io_enq_0_dec_uops_1_imm_packed,
  input  [11:0] io_enq_0_dec_uops_1_csr_addr,
  input  [5:0]  io_enq_0_dec_uops_1_rob_idx,
  input  [4:0]  io_enq_0_dec_uops_1_ldq_idx,
  input  [4:0]  io_enq_0_dec_uops_1_stq_idx,
  input  [1:0]  io_enq_0_dec_uops_1_rxq_idx,
  input  [6:0]  io_enq_0_dec_uops_1_pdst,
  input  [6:0]  io_enq_0_dec_uops_1_prs1,
  input  [6:0]  io_enq_0_dec_uops_1_prs2,
  input  [6:0]  io_enq_0_dec_uops_1_prs3,
  input  [4:0]  io_enq_0_dec_uops_1_ppred,
  input         io_enq_0_dec_uops_1_prs1_busy,
  input         io_enq_0_dec_uops_1_prs2_busy,
  input         io_enq_0_dec_uops_1_prs3_busy,
  input         io_enq_0_dec_uops_1_ppred_busy,
  input  [6:0]  io_enq_0_dec_uops_1_stale_pdst,
  input         io_enq_0_dec_uops_1_exception,
  input  [63:0] io_enq_0_dec_uops_1_exc_cause,
  input         io_enq_0_dec_uops_1_bypassable,
  input  [4:0]  io_enq_0_dec_uops_1_mem_cmd,
  input  [1:0]  io_enq_0_dec_uops_1_mem_size,
  input         io_enq_0_dec_uops_1_mem_signed,
  input         io_enq_0_dec_uops_1_is_fence,
  input         io_enq_0_dec_uops_1_is_fencei,
  input         io_enq_0_dec_uops_1_is_amo,
  input         io_enq_0_dec_uops_1_uses_ldq,
  input         io_enq_0_dec_uops_1_uses_stq,
  input         io_enq_0_dec_uops_1_is_sys_pc2epc,
  input         io_enq_0_dec_uops_1_is_unique,
  input         io_enq_0_dec_uops_1_flush_on_commit,
  input         io_enq_0_dec_uops_1_ldst_is_rs1,
  input  [5:0]  io_enq_0_dec_uops_1_ldst,
  input  [5:0]  io_enq_0_dec_uops_1_lrs1,
  input  [5:0]  io_enq_0_dec_uops_1_lrs2,
  input  [5:0]  io_enq_0_dec_uops_1_lrs3,
  input         io_enq_0_dec_uops_1_ldst_val,
  input  [1:0]  io_enq_0_dec_uops_1_dst_rtype,
  input  [1:0]  io_enq_0_dec_uops_1_lrs1_rtype,
  input  [1:0]  io_enq_0_dec_uops_1_lrs2_rtype,
  input         io_enq_0_dec_uops_1_frs3_en,
  input         io_enq_0_dec_uops_1_fp_val,
  input         io_enq_0_dec_uops_1_fp_single,
  input         io_enq_0_dec_uops_1_xcpt_pf_if,
  input         io_enq_0_dec_uops_1_xcpt_ae_if,
  input         io_enq_0_dec_uops_1_xcpt_ma_if,
  input         io_enq_0_dec_uops_1_bp_debug_if,
  input         io_enq_0_dec_uops_1_bp_xcpt_if,
  input  [1:0]  io_enq_0_dec_uops_1_debug_fsrc,
  input  [1:0]  io_enq_0_dec_uops_1_debug_tsrc,
  input         io_enq_0_dec_uops_2_switch,
  input         io_enq_0_dec_uops_2_switch_off,
  input         io_enq_0_dec_uops_2_is_unicore,
  input  [2:0]  io_enq_0_dec_uops_2_shift,
  input  [1:0]  io_enq_0_dec_uops_2_lrs3_rtype,
  input         io_enq_0_dec_uops_2_rflag,
  input         io_enq_0_dec_uops_2_wflag,
  input  [3:0]  io_enq_0_dec_uops_2_prflag,
  input  [3:0]  io_enq_0_dec_uops_2_pwflag,
  input         io_enq_0_dec_uops_2_pflag_busy,
  input  [3:0]  io_enq_0_dec_uops_2_stale_pflag,
  input  [3:0]  io_enq_0_dec_uops_2_op1_sel,
  input  [3:0]  io_enq_0_dec_uops_2_op2_sel,
  input  [5:0]  io_enq_0_dec_uops_2_split_num,
  input  [5:0]  io_enq_0_dec_uops_2_self_index,
  input  [5:0]  io_enq_0_dec_uops_2_rob_inst_idx,
  input  [5:0]  io_enq_0_dec_uops_2_address_num,
  input  [6:0]  io_enq_0_dec_uops_2_uopc,
  input  [31:0] io_enq_0_dec_uops_2_inst,
  input  [31:0] io_enq_0_dec_uops_2_debug_inst,
  input         io_enq_0_dec_uops_2_is_rvc,
  input  [39:0] io_enq_0_dec_uops_2_debug_pc,
  input  [2:0]  io_enq_0_dec_uops_2_iq_type,
  input  [9:0]  io_enq_0_dec_uops_2_fu_code,
  input  [3:0]  io_enq_0_dec_uops_2_ctrl_br_type,
  input  [1:0]  io_enq_0_dec_uops_2_ctrl_op1_sel,
  input  [2:0]  io_enq_0_dec_uops_2_ctrl_op2_sel,
  input  [2:0]  io_enq_0_dec_uops_2_ctrl_imm_sel,
  input  [3:0]  io_enq_0_dec_uops_2_ctrl_op_fcn,
  input         io_enq_0_dec_uops_2_ctrl_fcn_dw,
  input  [2:0]  io_enq_0_dec_uops_2_ctrl_csr_cmd,
  input         io_enq_0_dec_uops_2_ctrl_is_load,
  input         io_enq_0_dec_uops_2_ctrl_is_sta,
  input         io_enq_0_dec_uops_2_ctrl_is_std,
  input  [1:0]  io_enq_0_dec_uops_2_ctrl_op3_sel,
  input  [1:0]  io_enq_0_dec_uops_2_iw_state,
  input         io_enq_0_dec_uops_2_iw_p1_poisoned,
  input         io_enq_0_dec_uops_2_iw_p2_poisoned,
  input         io_enq_0_dec_uops_2_is_br,
  input         io_enq_0_dec_uops_2_is_jalr,
  input         io_enq_0_dec_uops_2_is_jal,
  input         io_enq_0_dec_uops_2_is_sfb,
  input  [11:0] io_enq_0_dec_uops_2_br_mask,
  input  [3:0]  io_enq_0_dec_uops_2_br_tag,
  input  [4:0]  io_enq_0_dec_uops_2_ftq_idx,
  input         io_enq_0_dec_uops_2_edge_inst,
  input  [5:0]  io_enq_0_dec_uops_2_pc_lob,
  input         io_enq_0_dec_uops_2_taken,
  input  [19:0] io_enq_0_dec_uops_2_imm_packed,
  input  [11:0] io_enq_0_dec_uops_2_csr_addr,
  input  [5:0]  io_enq_0_dec_uops_2_rob_idx,
  input  [4:0]  io_enq_0_dec_uops_2_ldq_idx,
  input  [4:0]  io_enq_0_dec_uops_2_stq_idx,
  input  [1:0]  io_enq_0_dec_uops_2_rxq_idx,
  input  [6:0]  io_enq_0_dec_uops_2_pdst,
  input  [6:0]  io_enq_0_dec_uops_2_prs1,
  input  [6:0]  io_enq_0_dec_uops_2_prs2,
  input  [6:0]  io_enq_0_dec_uops_2_prs3,
  input  [4:0]  io_enq_0_dec_uops_2_ppred,
  input         io_enq_0_dec_uops_2_prs1_busy,
  input         io_enq_0_dec_uops_2_prs2_busy,
  input         io_enq_0_dec_uops_2_prs3_busy,
  input         io_enq_0_dec_uops_2_ppred_busy,
  input  [6:0]  io_enq_0_dec_uops_2_stale_pdst,
  input         io_enq_0_dec_uops_2_exception,
  input  [63:0] io_enq_0_dec_uops_2_exc_cause,
  input         io_enq_0_dec_uops_2_bypassable,
  input  [4:0]  io_enq_0_dec_uops_2_mem_cmd,
  input  [1:0]  io_enq_0_dec_uops_2_mem_size,
  input         io_enq_0_dec_uops_2_mem_signed,
  input         io_enq_0_dec_uops_2_is_fence,
  input         io_enq_0_dec_uops_2_is_fencei,
  input         io_enq_0_dec_uops_2_is_amo,
  input         io_enq_0_dec_uops_2_uses_ldq,
  input         io_enq_0_dec_uops_2_uses_stq,
  input         io_enq_0_dec_uops_2_is_sys_pc2epc,
  input         io_enq_0_dec_uops_2_is_unique,
  input         io_enq_0_dec_uops_2_flush_on_commit,
  input         io_enq_0_dec_uops_2_ldst_is_rs1,
  input  [5:0]  io_enq_0_dec_uops_2_ldst,
  input  [5:0]  io_enq_0_dec_uops_2_lrs1,
  input  [5:0]  io_enq_0_dec_uops_2_lrs2,
  input  [5:0]  io_enq_0_dec_uops_2_lrs3,
  input         io_enq_0_dec_uops_2_ldst_val,
  input  [1:0]  io_enq_0_dec_uops_2_dst_rtype,
  input  [1:0]  io_enq_0_dec_uops_2_lrs1_rtype,
  input  [1:0]  io_enq_0_dec_uops_2_lrs2_rtype,
  input         io_enq_0_dec_uops_2_frs3_en,
  input         io_enq_0_dec_uops_2_fp_val,
  input         io_enq_0_dec_uops_2_fp_single,
  input         io_enq_0_dec_uops_2_xcpt_pf_if,
  input         io_enq_0_dec_uops_2_xcpt_ae_if,
  input         io_enq_0_dec_uops_2_xcpt_ma_if,
  input         io_enq_0_dec_uops_2_bp_debug_if,
  input         io_enq_0_dec_uops_2_bp_xcpt_if,
  input  [1:0]  io_enq_0_dec_uops_2_debug_fsrc,
  input  [1:0]  io_enq_0_dec_uops_2_debug_tsrc,
  input         io_enq_0_dec_uops_3_switch,
  input         io_enq_0_dec_uops_3_switch_off,
  input         io_enq_0_dec_uops_3_is_unicore,
  input  [2:0]  io_enq_0_dec_uops_3_shift,
  input  [1:0]  io_enq_0_dec_uops_3_lrs3_rtype,
  input         io_enq_0_dec_uops_3_rflag,
  input         io_enq_0_dec_uops_3_wflag,
  input  [3:0]  io_enq_0_dec_uops_3_prflag,
  input  [3:0]  io_enq_0_dec_uops_3_pwflag,
  input         io_enq_0_dec_uops_3_pflag_busy,
  input  [3:0]  io_enq_0_dec_uops_3_stale_pflag,
  input  [3:0]  io_enq_0_dec_uops_3_op1_sel,
  input  [3:0]  io_enq_0_dec_uops_3_op2_sel,
  input  [5:0]  io_enq_0_dec_uops_3_split_num,
  input  [5:0]  io_enq_0_dec_uops_3_self_index,
  input  [5:0]  io_enq_0_dec_uops_3_rob_inst_idx,
  input  [5:0]  io_enq_0_dec_uops_3_address_num,
  input  [6:0]  io_enq_0_dec_uops_3_uopc,
  input  [31:0] io_enq_0_dec_uops_3_inst,
  input  [31:0] io_enq_0_dec_uops_3_debug_inst,
  input         io_enq_0_dec_uops_3_is_rvc,
  input  [39:0] io_enq_0_dec_uops_3_debug_pc,
  input  [2:0]  io_enq_0_dec_uops_3_iq_type,
  input  [9:0]  io_enq_0_dec_uops_3_fu_code,
  input  [3:0]  io_enq_0_dec_uops_3_ctrl_br_type,
  input  [1:0]  io_enq_0_dec_uops_3_ctrl_op1_sel,
  input  [2:0]  io_enq_0_dec_uops_3_ctrl_op2_sel,
  input  [2:0]  io_enq_0_dec_uops_3_ctrl_imm_sel,
  input  [3:0]  io_enq_0_dec_uops_3_ctrl_op_fcn,
  input         io_enq_0_dec_uops_3_ctrl_fcn_dw,
  input  [2:0]  io_enq_0_dec_uops_3_ctrl_csr_cmd,
  input         io_enq_0_dec_uops_3_ctrl_is_load,
  input         io_enq_0_dec_uops_3_ctrl_is_sta,
  input         io_enq_0_dec_uops_3_ctrl_is_std,
  input  [1:0]  io_enq_0_dec_uops_3_ctrl_op3_sel,
  input  [1:0]  io_enq_0_dec_uops_3_iw_state,
  input         io_enq_0_dec_uops_3_iw_p1_poisoned,
  input         io_enq_0_dec_uops_3_iw_p2_poisoned,
  input         io_enq_0_dec_uops_3_is_br,
  input         io_enq_0_dec_uops_3_is_jalr,
  input         io_enq_0_dec_uops_3_is_jal,
  input         io_enq_0_dec_uops_3_is_sfb,
  input  [11:0] io_enq_0_dec_uops_3_br_mask,
  input  [3:0]  io_enq_0_dec_uops_3_br_tag,
  input  [4:0]  io_enq_0_dec_uops_3_ftq_idx,
  input         io_enq_0_dec_uops_3_edge_inst,
  input  [5:0]  io_enq_0_dec_uops_3_pc_lob,
  input         io_enq_0_dec_uops_3_taken,
  input  [19:0] io_enq_0_dec_uops_3_imm_packed,
  input  [11:0] io_enq_0_dec_uops_3_csr_addr,
  input  [5:0]  io_enq_0_dec_uops_3_rob_idx,
  input  [4:0]  io_enq_0_dec_uops_3_ldq_idx,
  input  [4:0]  io_enq_0_dec_uops_3_stq_idx,
  input  [1:0]  io_enq_0_dec_uops_3_rxq_idx,
  input  [6:0]  io_enq_0_dec_uops_3_pdst,
  input  [6:0]  io_enq_0_dec_uops_3_prs1,
  input  [6:0]  io_enq_0_dec_uops_3_prs2,
  input  [6:0]  io_enq_0_dec_uops_3_prs3,
  input  [4:0]  io_enq_0_dec_uops_3_ppred,
  input         io_enq_0_dec_uops_3_prs1_busy,
  input         io_enq_0_dec_uops_3_prs2_busy,
  input         io_enq_0_dec_uops_3_prs3_busy,
  input         io_enq_0_dec_uops_3_ppred_busy,
  input  [6:0]  io_enq_0_dec_uops_3_stale_pdst,
  input         io_enq_0_dec_uops_3_exception,
  input  [63:0] io_enq_0_dec_uops_3_exc_cause,
  input         io_enq_0_dec_uops_3_bypassable,
  input  [4:0]  io_enq_0_dec_uops_3_mem_cmd,
  input  [1:0]  io_enq_0_dec_uops_3_mem_size,
  input         io_enq_0_dec_uops_3_mem_signed,
  input         io_enq_0_dec_uops_3_is_fence,
  input         io_enq_0_dec_uops_3_is_fencei,
  input         io_enq_0_dec_uops_3_is_amo,
  input         io_enq_0_dec_uops_3_uses_ldq,
  input         io_enq_0_dec_uops_3_uses_stq,
  input         io_enq_0_dec_uops_3_is_sys_pc2epc,
  input         io_enq_0_dec_uops_3_is_unique,
  input         io_enq_0_dec_uops_3_flush_on_commit,
  input         io_enq_0_dec_uops_3_ldst_is_rs1,
  input  [5:0]  io_enq_0_dec_uops_3_ldst,
  input  [5:0]  io_enq_0_dec_uops_3_lrs1,
  input  [5:0]  io_enq_0_dec_uops_3_lrs2,
  input  [5:0]  io_enq_0_dec_uops_3_lrs3,
  input         io_enq_0_dec_uops_3_ldst_val,
  input  [1:0]  io_enq_0_dec_uops_3_dst_rtype,
  input  [1:0]  io_enq_0_dec_uops_3_lrs1_rtype,
  input  [1:0]  io_enq_0_dec_uops_3_lrs2_rtype,
  input         io_enq_0_dec_uops_3_frs3_en,
  input         io_enq_0_dec_uops_3_fp_val,
  input         io_enq_0_dec_uops_3_fp_single,
  input         io_enq_0_dec_uops_3_xcpt_pf_if,
  input         io_enq_0_dec_uops_3_xcpt_ae_if,
  input         io_enq_0_dec_uops_3_xcpt_ma_if,
  input         io_enq_0_dec_uops_3_bp_debug_if,
  input         io_enq_0_dec_uops_3_bp_xcpt_if,
  input  [1:0]  io_enq_0_dec_uops_3_debug_fsrc,
  input  [1:0]  io_enq_0_dec_uops_3_debug_tsrc,
  input         io_enq_0_val_mask_0,
  input         io_enq_0_val_mask_1,
  input         io_enq_0_val_mask_2,
  input         io_enq_0_val_mask_3,
  input         io_enq_1_dec_uops_0_switch,
  input         io_enq_1_dec_uops_0_switch_off,
  input         io_enq_1_dec_uops_0_is_unicore,
  input  [2:0]  io_enq_1_dec_uops_0_shift,
  input  [1:0]  io_enq_1_dec_uops_0_lrs3_rtype,
  input         io_enq_1_dec_uops_0_rflag,
  input         io_enq_1_dec_uops_0_wflag,
  input  [3:0]  io_enq_1_dec_uops_0_prflag,
  input  [3:0]  io_enq_1_dec_uops_0_pwflag,
  input         io_enq_1_dec_uops_0_pflag_busy,
  input  [3:0]  io_enq_1_dec_uops_0_stale_pflag,
  input  [3:0]  io_enq_1_dec_uops_0_op1_sel,
  input  [3:0]  io_enq_1_dec_uops_0_op2_sel,
  input  [5:0]  io_enq_1_dec_uops_0_split_num,
  input  [5:0]  io_enq_1_dec_uops_0_self_index,
  input  [5:0]  io_enq_1_dec_uops_0_rob_inst_idx,
  input  [5:0]  io_enq_1_dec_uops_0_address_num,
  input  [6:0]  io_enq_1_dec_uops_0_uopc,
  input  [31:0] io_enq_1_dec_uops_0_inst,
  input  [31:0] io_enq_1_dec_uops_0_debug_inst,
  input         io_enq_1_dec_uops_0_is_rvc,
  input  [39:0] io_enq_1_dec_uops_0_debug_pc,
  input  [2:0]  io_enq_1_dec_uops_0_iq_type,
  input  [9:0]  io_enq_1_dec_uops_0_fu_code,
  input  [3:0]  io_enq_1_dec_uops_0_ctrl_br_type,
  input  [1:0]  io_enq_1_dec_uops_0_ctrl_op1_sel,
  input  [2:0]  io_enq_1_dec_uops_0_ctrl_op2_sel,
  input  [2:0]  io_enq_1_dec_uops_0_ctrl_imm_sel,
  input  [3:0]  io_enq_1_dec_uops_0_ctrl_op_fcn,
  input         io_enq_1_dec_uops_0_ctrl_fcn_dw,
  input  [2:0]  io_enq_1_dec_uops_0_ctrl_csr_cmd,
  input         io_enq_1_dec_uops_0_ctrl_is_load,
  input         io_enq_1_dec_uops_0_ctrl_is_sta,
  input         io_enq_1_dec_uops_0_ctrl_is_std,
  input  [1:0]  io_enq_1_dec_uops_0_ctrl_op3_sel,
  input  [1:0]  io_enq_1_dec_uops_0_iw_state,
  input         io_enq_1_dec_uops_0_iw_p1_poisoned,
  input         io_enq_1_dec_uops_0_iw_p2_poisoned,
  input         io_enq_1_dec_uops_0_is_br,
  input         io_enq_1_dec_uops_0_is_jalr,
  input         io_enq_1_dec_uops_0_is_jal,
  input         io_enq_1_dec_uops_0_is_sfb,
  input  [11:0] io_enq_1_dec_uops_0_br_mask,
  input  [3:0]  io_enq_1_dec_uops_0_br_tag,
  input  [4:0]  io_enq_1_dec_uops_0_ftq_idx,
  input         io_enq_1_dec_uops_0_edge_inst,
  input  [5:0]  io_enq_1_dec_uops_0_pc_lob,
  input         io_enq_1_dec_uops_0_taken,
  input  [19:0] io_enq_1_dec_uops_0_imm_packed,
  input  [11:0] io_enq_1_dec_uops_0_csr_addr,
  input  [5:0]  io_enq_1_dec_uops_0_rob_idx,
  input  [4:0]  io_enq_1_dec_uops_0_ldq_idx,
  input  [4:0]  io_enq_1_dec_uops_0_stq_idx,
  input  [1:0]  io_enq_1_dec_uops_0_rxq_idx,
  input  [6:0]  io_enq_1_dec_uops_0_pdst,
  input  [6:0]  io_enq_1_dec_uops_0_prs1,
  input  [6:0]  io_enq_1_dec_uops_0_prs2,
  input  [6:0]  io_enq_1_dec_uops_0_prs3,
  input  [4:0]  io_enq_1_dec_uops_0_ppred,
  input         io_enq_1_dec_uops_0_prs1_busy,
  input         io_enq_1_dec_uops_0_prs2_busy,
  input         io_enq_1_dec_uops_0_prs3_busy,
  input         io_enq_1_dec_uops_0_ppred_busy,
  input  [6:0]  io_enq_1_dec_uops_0_stale_pdst,
  input         io_enq_1_dec_uops_0_exception,
  input  [63:0] io_enq_1_dec_uops_0_exc_cause,
  input         io_enq_1_dec_uops_0_bypassable,
  input  [4:0]  io_enq_1_dec_uops_0_mem_cmd,
  input  [1:0]  io_enq_1_dec_uops_0_mem_size,
  input         io_enq_1_dec_uops_0_mem_signed,
  input         io_enq_1_dec_uops_0_is_fence,
  input         io_enq_1_dec_uops_0_is_fencei,
  input         io_enq_1_dec_uops_0_is_amo,
  input         io_enq_1_dec_uops_0_uses_ldq,
  input         io_enq_1_dec_uops_0_uses_stq,
  input         io_enq_1_dec_uops_0_is_sys_pc2epc,
  input         io_enq_1_dec_uops_0_is_unique,
  input         io_enq_1_dec_uops_0_flush_on_commit,
  input         io_enq_1_dec_uops_0_ldst_is_rs1,
  input  [5:0]  io_enq_1_dec_uops_0_ldst,
  input  [5:0]  io_enq_1_dec_uops_0_lrs1,
  input  [5:0]  io_enq_1_dec_uops_0_lrs2,
  input  [5:0]  io_enq_1_dec_uops_0_lrs3,
  input         io_enq_1_dec_uops_0_ldst_val,
  input  [1:0]  io_enq_1_dec_uops_0_dst_rtype,
  input  [1:0]  io_enq_1_dec_uops_0_lrs1_rtype,
  input  [1:0]  io_enq_1_dec_uops_0_lrs2_rtype,
  input         io_enq_1_dec_uops_0_frs3_en,
  input         io_enq_1_dec_uops_0_fp_val,
  input         io_enq_1_dec_uops_0_fp_single,
  input         io_enq_1_dec_uops_0_xcpt_pf_if,
  input         io_enq_1_dec_uops_0_xcpt_ae_if,
  input         io_enq_1_dec_uops_0_xcpt_ma_if,
  input         io_enq_1_dec_uops_0_bp_debug_if,
  input         io_enq_1_dec_uops_0_bp_xcpt_if,
  input  [1:0]  io_enq_1_dec_uops_0_debug_fsrc,
  input  [1:0]  io_enq_1_dec_uops_0_debug_tsrc,
  input         io_enq_1_dec_uops_1_switch,
  input         io_enq_1_dec_uops_1_switch_off,
  input         io_enq_1_dec_uops_1_is_unicore,
  input  [2:0]  io_enq_1_dec_uops_1_shift,
  input  [1:0]  io_enq_1_dec_uops_1_lrs3_rtype,
  input         io_enq_1_dec_uops_1_rflag,
  input         io_enq_1_dec_uops_1_wflag,
  input  [3:0]  io_enq_1_dec_uops_1_prflag,
  input  [3:0]  io_enq_1_dec_uops_1_pwflag,
  input         io_enq_1_dec_uops_1_pflag_busy,
  input  [3:0]  io_enq_1_dec_uops_1_stale_pflag,
  input  [3:0]  io_enq_1_dec_uops_1_op1_sel,
  input  [3:0]  io_enq_1_dec_uops_1_op2_sel,
  input  [5:0]  io_enq_1_dec_uops_1_split_num,
  input  [5:0]  io_enq_1_dec_uops_1_self_index,
  input  [5:0]  io_enq_1_dec_uops_1_rob_inst_idx,
  input  [5:0]  io_enq_1_dec_uops_1_address_num,
  input  [6:0]  io_enq_1_dec_uops_1_uopc,
  input  [31:0] io_enq_1_dec_uops_1_inst,
  input  [31:0] io_enq_1_dec_uops_1_debug_inst,
  input         io_enq_1_dec_uops_1_is_rvc,
  input  [39:0] io_enq_1_dec_uops_1_debug_pc,
  input  [2:0]  io_enq_1_dec_uops_1_iq_type,
  input  [9:0]  io_enq_1_dec_uops_1_fu_code,
  input  [3:0]  io_enq_1_dec_uops_1_ctrl_br_type,
  input  [1:0]  io_enq_1_dec_uops_1_ctrl_op1_sel,
  input  [2:0]  io_enq_1_dec_uops_1_ctrl_op2_sel,
  input  [2:0]  io_enq_1_dec_uops_1_ctrl_imm_sel,
  input  [3:0]  io_enq_1_dec_uops_1_ctrl_op_fcn,
  input         io_enq_1_dec_uops_1_ctrl_fcn_dw,
  input  [2:0]  io_enq_1_dec_uops_1_ctrl_csr_cmd,
  input         io_enq_1_dec_uops_1_ctrl_is_load,
  input         io_enq_1_dec_uops_1_ctrl_is_sta,
  input         io_enq_1_dec_uops_1_ctrl_is_std,
  input  [1:0]  io_enq_1_dec_uops_1_ctrl_op3_sel,
  input  [1:0]  io_enq_1_dec_uops_1_iw_state,
  input         io_enq_1_dec_uops_1_iw_p1_poisoned,
  input         io_enq_1_dec_uops_1_iw_p2_poisoned,
  input         io_enq_1_dec_uops_1_is_br,
  input         io_enq_1_dec_uops_1_is_jalr,
  input         io_enq_1_dec_uops_1_is_jal,
  input         io_enq_1_dec_uops_1_is_sfb,
  input  [11:0] io_enq_1_dec_uops_1_br_mask,
  input  [3:0]  io_enq_1_dec_uops_1_br_tag,
  input  [4:0]  io_enq_1_dec_uops_1_ftq_idx,
  input         io_enq_1_dec_uops_1_edge_inst,
  input  [5:0]  io_enq_1_dec_uops_1_pc_lob,
  input         io_enq_1_dec_uops_1_taken,
  input  [19:0] io_enq_1_dec_uops_1_imm_packed,
  input  [11:0] io_enq_1_dec_uops_1_csr_addr,
  input  [5:0]  io_enq_1_dec_uops_1_rob_idx,
  input  [4:0]  io_enq_1_dec_uops_1_ldq_idx,
  input  [4:0]  io_enq_1_dec_uops_1_stq_idx,
  input  [1:0]  io_enq_1_dec_uops_1_rxq_idx,
  input  [6:0]  io_enq_1_dec_uops_1_pdst,
  input  [6:0]  io_enq_1_dec_uops_1_prs1,
  input  [6:0]  io_enq_1_dec_uops_1_prs2,
  input  [6:0]  io_enq_1_dec_uops_1_prs3,
  input  [4:0]  io_enq_1_dec_uops_1_ppred,
  input         io_enq_1_dec_uops_1_prs1_busy,
  input         io_enq_1_dec_uops_1_prs2_busy,
  input         io_enq_1_dec_uops_1_prs3_busy,
  input         io_enq_1_dec_uops_1_ppred_busy,
  input  [6:0]  io_enq_1_dec_uops_1_stale_pdst,
  input         io_enq_1_dec_uops_1_exception,
  input  [63:0] io_enq_1_dec_uops_1_exc_cause,
  input         io_enq_1_dec_uops_1_bypassable,
  input  [4:0]  io_enq_1_dec_uops_1_mem_cmd,
  input  [1:0]  io_enq_1_dec_uops_1_mem_size,
  input         io_enq_1_dec_uops_1_mem_signed,
  input         io_enq_1_dec_uops_1_is_fence,
  input         io_enq_1_dec_uops_1_is_fencei,
  input         io_enq_1_dec_uops_1_is_amo,
  input         io_enq_1_dec_uops_1_uses_ldq,
  input         io_enq_1_dec_uops_1_uses_stq,
  input         io_enq_1_dec_uops_1_is_sys_pc2epc,
  input         io_enq_1_dec_uops_1_is_unique,
  input         io_enq_1_dec_uops_1_flush_on_commit,
  input         io_enq_1_dec_uops_1_ldst_is_rs1,
  input  [5:0]  io_enq_1_dec_uops_1_ldst,
  input  [5:0]  io_enq_1_dec_uops_1_lrs1,
  input  [5:0]  io_enq_1_dec_uops_1_lrs2,
  input  [5:0]  io_enq_1_dec_uops_1_lrs3,
  input         io_enq_1_dec_uops_1_ldst_val,
  input  [1:0]  io_enq_1_dec_uops_1_dst_rtype,
  input  [1:0]  io_enq_1_dec_uops_1_lrs1_rtype,
  input  [1:0]  io_enq_1_dec_uops_1_lrs2_rtype,
  input         io_enq_1_dec_uops_1_frs3_en,
  input         io_enq_1_dec_uops_1_fp_val,
  input         io_enq_1_dec_uops_1_fp_single,
  input         io_enq_1_dec_uops_1_xcpt_pf_if,
  input         io_enq_1_dec_uops_1_xcpt_ae_if,
  input         io_enq_1_dec_uops_1_xcpt_ma_if,
  input         io_enq_1_dec_uops_1_bp_debug_if,
  input         io_enq_1_dec_uops_1_bp_xcpt_if,
  input  [1:0]  io_enq_1_dec_uops_1_debug_fsrc,
  input  [1:0]  io_enq_1_dec_uops_1_debug_tsrc,
  input         io_enq_1_dec_uops_2_switch,
  input         io_enq_1_dec_uops_2_switch_off,
  input         io_enq_1_dec_uops_2_is_unicore,
  input  [2:0]  io_enq_1_dec_uops_2_shift,
  input  [1:0]  io_enq_1_dec_uops_2_lrs3_rtype,
  input         io_enq_1_dec_uops_2_rflag,
  input         io_enq_1_dec_uops_2_wflag,
  input  [3:0]  io_enq_1_dec_uops_2_prflag,
  input  [3:0]  io_enq_1_dec_uops_2_pwflag,
  input         io_enq_1_dec_uops_2_pflag_busy,
  input  [3:0]  io_enq_1_dec_uops_2_stale_pflag,
  input  [3:0]  io_enq_1_dec_uops_2_op1_sel,
  input  [3:0]  io_enq_1_dec_uops_2_op2_sel,
  input  [5:0]  io_enq_1_dec_uops_2_split_num,
  input  [5:0]  io_enq_1_dec_uops_2_self_index,
  input  [5:0]  io_enq_1_dec_uops_2_rob_inst_idx,
  input  [5:0]  io_enq_1_dec_uops_2_address_num,
  input  [6:0]  io_enq_1_dec_uops_2_uopc,
  input  [31:0] io_enq_1_dec_uops_2_inst,
  input  [31:0] io_enq_1_dec_uops_2_debug_inst,
  input         io_enq_1_dec_uops_2_is_rvc,
  input  [39:0] io_enq_1_dec_uops_2_debug_pc,
  input  [2:0]  io_enq_1_dec_uops_2_iq_type,
  input  [9:0]  io_enq_1_dec_uops_2_fu_code,
  input  [3:0]  io_enq_1_dec_uops_2_ctrl_br_type,
  input  [1:0]  io_enq_1_dec_uops_2_ctrl_op1_sel,
  input  [2:0]  io_enq_1_dec_uops_2_ctrl_op2_sel,
  input  [2:0]  io_enq_1_dec_uops_2_ctrl_imm_sel,
  input  [3:0]  io_enq_1_dec_uops_2_ctrl_op_fcn,
  input         io_enq_1_dec_uops_2_ctrl_fcn_dw,
  input  [2:0]  io_enq_1_dec_uops_2_ctrl_csr_cmd,
  input         io_enq_1_dec_uops_2_ctrl_is_load,
  input         io_enq_1_dec_uops_2_ctrl_is_sta,
  input         io_enq_1_dec_uops_2_ctrl_is_std,
  input  [1:0]  io_enq_1_dec_uops_2_ctrl_op3_sel,
  input  [1:0]  io_enq_1_dec_uops_2_iw_state,
  input         io_enq_1_dec_uops_2_iw_p1_poisoned,
  input         io_enq_1_dec_uops_2_iw_p2_poisoned,
  input         io_enq_1_dec_uops_2_is_br,
  input         io_enq_1_dec_uops_2_is_jalr,
  input         io_enq_1_dec_uops_2_is_jal,
  input         io_enq_1_dec_uops_2_is_sfb,
  input  [11:0] io_enq_1_dec_uops_2_br_mask,
  input  [3:0]  io_enq_1_dec_uops_2_br_tag,
  input  [4:0]  io_enq_1_dec_uops_2_ftq_idx,
  input         io_enq_1_dec_uops_2_edge_inst,
  input  [5:0]  io_enq_1_dec_uops_2_pc_lob,
  input         io_enq_1_dec_uops_2_taken,
  input  [19:0] io_enq_1_dec_uops_2_imm_packed,
  input  [11:0] io_enq_1_dec_uops_2_csr_addr,
  input  [5:0]  io_enq_1_dec_uops_2_rob_idx,
  input  [4:0]  io_enq_1_dec_uops_2_ldq_idx,
  input  [4:0]  io_enq_1_dec_uops_2_stq_idx,
  input  [1:0]  io_enq_1_dec_uops_2_rxq_idx,
  input  [6:0]  io_enq_1_dec_uops_2_pdst,
  input  [6:0]  io_enq_1_dec_uops_2_prs1,
  input  [6:0]  io_enq_1_dec_uops_2_prs2,
  input  [6:0]  io_enq_1_dec_uops_2_prs3,
  input  [4:0]  io_enq_1_dec_uops_2_ppred,
  input         io_enq_1_dec_uops_2_prs1_busy,
  input         io_enq_1_dec_uops_2_prs2_busy,
  input         io_enq_1_dec_uops_2_prs3_busy,
  input         io_enq_1_dec_uops_2_ppred_busy,
  input  [6:0]  io_enq_1_dec_uops_2_stale_pdst,
  input         io_enq_1_dec_uops_2_exception,
  input  [63:0] io_enq_1_dec_uops_2_exc_cause,
  input         io_enq_1_dec_uops_2_bypassable,
  input  [4:0]  io_enq_1_dec_uops_2_mem_cmd,
  input  [1:0]  io_enq_1_dec_uops_2_mem_size,
  input         io_enq_1_dec_uops_2_mem_signed,
  input         io_enq_1_dec_uops_2_is_fence,
  input         io_enq_1_dec_uops_2_is_fencei,
  input         io_enq_1_dec_uops_2_is_amo,
  input         io_enq_1_dec_uops_2_uses_ldq,
  input         io_enq_1_dec_uops_2_uses_stq,
  input         io_enq_1_dec_uops_2_is_sys_pc2epc,
  input         io_enq_1_dec_uops_2_is_unique,
  input         io_enq_1_dec_uops_2_flush_on_commit,
  input         io_enq_1_dec_uops_2_ldst_is_rs1,
  input  [5:0]  io_enq_1_dec_uops_2_ldst,
  input  [5:0]  io_enq_1_dec_uops_2_lrs1,
  input  [5:0]  io_enq_1_dec_uops_2_lrs2,
  input  [5:0]  io_enq_1_dec_uops_2_lrs3,
  input         io_enq_1_dec_uops_2_ldst_val,
  input  [1:0]  io_enq_1_dec_uops_2_dst_rtype,
  input  [1:0]  io_enq_1_dec_uops_2_lrs1_rtype,
  input  [1:0]  io_enq_1_dec_uops_2_lrs2_rtype,
  input         io_enq_1_dec_uops_2_frs3_en,
  input         io_enq_1_dec_uops_2_fp_val,
  input         io_enq_1_dec_uops_2_fp_single,
  input         io_enq_1_dec_uops_2_xcpt_pf_if,
  input         io_enq_1_dec_uops_2_xcpt_ae_if,
  input         io_enq_1_dec_uops_2_xcpt_ma_if,
  input         io_enq_1_dec_uops_2_bp_debug_if,
  input         io_enq_1_dec_uops_2_bp_xcpt_if,
  input  [1:0]  io_enq_1_dec_uops_2_debug_fsrc,
  input  [1:0]  io_enq_1_dec_uops_2_debug_tsrc,
  input         io_enq_1_dec_uops_3_switch,
  input         io_enq_1_dec_uops_3_switch_off,
  input         io_enq_1_dec_uops_3_is_unicore,
  input  [2:0]  io_enq_1_dec_uops_3_shift,
  input  [1:0]  io_enq_1_dec_uops_3_lrs3_rtype,
  input         io_enq_1_dec_uops_3_rflag,
  input         io_enq_1_dec_uops_3_wflag,
  input  [3:0]  io_enq_1_dec_uops_3_prflag,
  input  [3:0]  io_enq_1_dec_uops_3_pwflag,
  input         io_enq_1_dec_uops_3_pflag_busy,
  input  [3:0]  io_enq_1_dec_uops_3_stale_pflag,
  input  [3:0]  io_enq_1_dec_uops_3_op1_sel,
  input  [3:0]  io_enq_1_dec_uops_3_op2_sel,
  input  [5:0]  io_enq_1_dec_uops_3_split_num,
  input  [5:0]  io_enq_1_dec_uops_3_self_index,
  input  [5:0]  io_enq_1_dec_uops_3_rob_inst_idx,
  input  [5:0]  io_enq_1_dec_uops_3_address_num,
  input  [6:0]  io_enq_1_dec_uops_3_uopc,
  input  [31:0] io_enq_1_dec_uops_3_inst,
  input  [31:0] io_enq_1_dec_uops_3_debug_inst,
  input         io_enq_1_dec_uops_3_is_rvc,
  input  [39:0] io_enq_1_dec_uops_3_debug_pc,
  input  [2:0]  io_enq_1_dec_uops_3_iq_type,
  input  [9:0]  io_enq_1_dec_uops_3_fu_code,
  input  [3:0]  io_enq_1_dec_uops_3_ctrl_br_type,
  input  [1:0]  io_enq_1_dec_uops_3_ctrl_op1_sel,
  input  [2:0]  io_enq_1_dec_uops_3_ctrl_op2_sel,
  input  [2:0]  io_enq_1_dec_uops_3_ctrl_imm_sel,
  input  [3:0]  io_enq_1_dec_uops_3_ctrl_op_fcn,
  input         io_enq_1_dec_uops_3_ctrl_fcn_dw,
  input  [2:0]  io_enq_1_dec_uops_3_ctrl_csr_cmd,
  input         io_enq_1_dec_uops_3_ctrl_is_load,
  input         io_enq_1_dec_uops_3_ctrl_is_sta,
  input         io_enq_1_dec_uops_3_ctrl_is_std,
  input  [1:0]  io_enq_1_dec_uops_3_ctrl_op3_sel,
  input  [1:0]  io_enq_1_dec_uops_3_iw_state,
  input         io_enq_1_dec_uops_3_iw_p1_poisoned,
  input         io_enq_1_dec_uops_3_iw_p2_poisoned,
  input         io_enq_1_dec_uops_3_is_br,
  input         io_enq_1_dec_uops_3_is_jalr,
  input         io_enq_1_dec_uops_3_is_jal,
  input         io_enq_1_dec_uops_3_is_sfb,
  input  [11:0] io_enq_1_dec_uops_3_br_mask,
  input  [3:0]  io_enq_1_dec_uops_3_br_tag,
  input  [4:0]  io_enq_1_dec_uops_3_ftq_idx,
  input         io_enq_1_dec_uops_3_edge_inst,
  input  [5:0]  io_enq_1_dec_uops_3_pc_lob,
  input         io_enq_1_dec_uops_3_taken,
  input  [19:0] io_enq_1_dec_uops_3_imm_packed,
  input  [11:0] io_enq_1_dec_uops_3_csr_addr,
  input  [5:0]  io_enq_1_dec_uops_3_rob_idx,
  input  [4:0]  io_enq_1_dec_uops_3_ldq_idx,
  input  [4:0]  io_enq_1_dec_uops_3_stq_idx,
  input  [1:0]  io_enq_1_dec_uops_3_rxq_idx,
  input  [6:0]  io_enq_1_dec_uops_3_pdst,
  input  [6:0]  io_enq_1_dec_uops_3_prs1,
  input  [6:0]  io_enq_1_dec_uops_3_prs2,
  input  [6:0]  io_enq_1_dec_uops_3_prs3,
  input  [4:0]  io_enq_1_dec_uops_3_ppred,
  input         io_enq_1_dec_uops_3_prs1_busy,
  input         io_enq_1_dec_uops_3_prs2_busy,
  input         io_enq_1_dec_uops_3_prs3_busy,
  input         io_enq_1_dec_uops_3_ppred_busy,
  input  [6:0]  io_enq_1_dec_uops_3_stale_pdst,
  input         io_enq_1_dec_uops_3_exception,
  input  [63:0] io_enq_1_dec_uops_3_exc_cause,
  input         io_enq_1_dec_uops_3_bypassable,
  input  [4:0]  io_enq_1_dec_uops_3_mem_cmd,
  input  [1:0]  io_enq_1_dec_uops_3_mem_size,
  input         io_enq_1_dec_uops_3_mem_signed,
  input         io_enq_1_dec_uops_3_is_fence,
  input         io_enq_1_dec_uops_3_is_fencei,
  input         io_enq_1_dec_uops_3_is_amo,
  input         io_enq_1_dec_uops_3_uses_ldq,
  input         io_enq_1_dec_uops_3_uses_stq,
  input         io_enq_1_dec_uops_3_is_sys_pc2epc,
  input         io_enq_1_dec_uops_3_is_unique,
  input         io_enq_1_dec_uops_3_flush_on_commit,
  input         io_enq_1_dec_uops_3_ldst_is_rs1,
  input  [5:0]  io_enq_1_dec_uops_3_ldst,
  input  [5:0]  io_enq_1_dec_uops_3_lrs1,
  input  [5:0]  io_enq_1_dec_uops_3_lrs2,
  input  [5:0]  io_enq_1_dec_uops_3_lrs3,
  input         io_enq_1_dec_uops_3_ldst_val,
  input  [1:0]  io_enq_1_dec_uops_3_dst_rtype,
  input  [1:0]  io_enq_1_dec_uops_3_lrs1_rtype,
  input  [1:0]  io_enq_1_dec_uops_3_lrs2_rtype,
  input         io_enq_1_dec_uops_3_frs3_en,
  input         io_enq_1_dec_uops_3_fp_val,
  input         io_enq_1_dec_uops_3_fp_single,
  input         io_enq_1_dec_uops_3_xcpt_pf_if,
  input         io_enq_1_dec_uops_3_xcpt_ae_if,
  input         io_enq_1_dec_uops_3_xcpt_ma_if,
  input         io_enq_1_dec_uops_3_bp_debug_if,
  input         io_enq_1_dec_uops_3_bp_xcpt_if,
  input  [1:0]  io_enq_1_dec_uops_3_debug_fsrc,
  input  [1:0]  io_enq_1_dec_uops_3_debug_tsrc,
  input         io_enq_1_val_mask_0,
  input         io_enq_1_val_mask_1,
  input         io_enq_1_val_mask_2,
  input         io_enq_1_val_mask_3,
  input         io_enq_2_dec_uops_0_switch,
  input         io_enq_2_dec_uops_0_switch_off,
  input         io_enq_2_dec_uops_0_is_unicore,
  input  [2:0]  io_enq_2_dec_uops_0_shift,
  input  [1:0]  io_enq_2_dec_uops_0_lrs3_rtype,
  input         io_enq_2_dec_uops_0_rflag,
  input         io_enq_2_dec_uops_0_wflag,
  input  [3:0]  io_enq_2_dec_uops_0_prflag,
  input  [3:0]  io_enq_2_dec_uops_0_pwflag,
  input         io_enq_2_dec_uops_0_pflag_busy,
  input  [3:0]  io_enq_2_dec_uops_0_stale_pflag,
  input  [3:0]  io_enq_2_dec_uops_0_op1_sel,
  input  [3:0]  io_enq_2_dec_uops_0_op2_sel,
  input  [5:0]  io_enq_2_dec_uops_0_split_num,
  input  [5:0]  io_enq_2_dec_uops_0_self_index,
  input  [5:0]  io_enq_2_dec_uops_0_rob_inst_idx,
  input  [5:0]  io_enq_2_dec_uops_0_address_num,
  input  [6:0]  io_enq_2_dec_uops_0_uopc,
  input  [31:0] io_enq_2_dec_uops_0_inst,
  input  [31:0] io_enq_2_dec_uops_0_debug_inst,
  input         io_enq_2_dec_uops_0_is_rvc,
  input  [39:0] io_enq_2_dec_uops_0_debug_pc,
  input  [2:0]  io_enq_2_dec_uops_0_iq_type,
  input  [9:0]  io_enq_2_dec_uops_0_fu_code,
  input  [3:0]  io_enq_2_dec_uops_0_ctrl_br_type,
  input  [1:0]  io_enq_2_dec_uops_0_ctrl_op1_sel,
  input  [2:0]  io_enq_2_dec_uops_0_ctrl_op2_sel,
  input  [2:0]  io_enq_2_dec_uops_0_ctrl_imm_sel,
  input  [3:0]  io_enq_2_dec_uops_0_ctrl_op_fcn,
  input         io_enq_2_dec_uops_0_ctrl_fcn_dw,
  input  [2:0]  io_enq_2_dec_uops_0_ctrl_csr_cmd,
  input         io_enq_2_dec_uops_0_ctrl_is_load,
  input         io_enq_2_dec_uops_0_ctrl_is_sta,
  input         io_enq_2_dec_uops_0_ctrl_is_std,
  input  [1:0]  io_enq_2_dec_uops_0_ctrl_op3_sel,
  input  [1:0]  io_enq_2_dec_uops_0_iw_state,
  input         io_enq_2_dec_uops_0_iw_p1_poisoned,
  input         io_enq_2_dec_uops_0_iw_p2_poisoned,
  input         io_enq_2_dec_uops_0_is_br,
  input         io_enq_2_dec_uops_0_is_jalr,
  input         io_enq_2_dec_uops_0_is_jal,
  input         io_enq_2_dec_uops_0_is_sfb,
  input  [11:0] io_enq_2_dec_uops_0_br_mask,
  input  [3:0]  io_enq_2_dec_uops_0_br_tag,
  input  [4:0]  io_enq_2_dec_uops_0_ftq_idx,
  input         io_enq_2_dec_uops_0_edge_inst,
  input  [5:0]  io_enq_2_dec_uops_0_pc_lob,
  input         io_enq_2_dec_uops_0_taken,
  input  [19:0] io_enq_2_dec_uops_0_imm_packed,
  input  [11:0] io_enq_2_dec_uops_0_csr_addr,
  input  [5:0]  io_enq_2_dec_uops_0_rob_idx,
  input  [4:0]  io_enq_2_dec_uops_0_ldq_idx,
  input  [4:0]  io_enq_2_dec_uops_0_stq_idx,
  input  [1:0]  io_enq_2_dec_uops_0_rxq_idx,
  input  [6:0]  io_enq_2_dec_uops_0_pdst,
  input  [6:0]  io_enq_2_dec_uops_0_prs1,
  input  [6:0]  io_enq_2_dec_uops_0_prs2,
  input  [6:0]  io_enq_2_dec_uops_0_prs3,
  input  [4:0]  io_enq_2_dec_uops_0_ppred,
  input         io_enq_2_dec_uops_0_prs1_busy,
  input         io_enq_2_dec_uops_0_prs2_busy,
  input         io_enq_2_dec_uops_0_prs3_busy,
  input         io_enq_2_dec_uops_0_ppred_busy,
  input  [6:0]  io_enq_2_dec_uops_0_stale_pdst,
  input         io_enq_2_dec_uops_0_exception,
  input  [63:0] io_enq_2_dec_uops_0_exc_cause,
  input         io_enq_2_dec_uops_0_bypassable,
  input  [4:0]  io_enq_2_dec_uops_0_mem_cmd,
  input  [1:0]  io_enq_2_dec_uops_0_mem_size,
  input         io_enq_2_dec_uops_0_mem_signed,
  input         io_enq_2_dec_uops_0_is_fence,
  input         io_enq_2_dec_uops_0_is_fencei,
  input         io_enq_2_dec_uops_0_is_amo,
  input         io_enq_2_dec_uops_0_uses_ldq,
  input         io_enq_2_dec_uops_0_uses_stq,
  input         io_enq_2_dec_uops_0_is_sys_pc2epc,
  input         io_enq_2_dec_uops_0_is_unique,
  input         io_enq_2_dec_uops_0_flush_on_commit,
  input         io_enq_2_dec_uops_0_ldst_is_rs1,
  input  [5:0]  io_enq_2_dec_uops_0_ldst,
  input  [5:0]  io_enq_2_dec_uops_0_lrs1,
  input  [5:0]  io_enq_2_dec_uops_0_lrs2,
  input  [5:0]  io_enq_2_dec_uops_0_lrs3,
  input         io_enq_2_dec_uops_0_ldst_val,
  input  [1:0]  io_enq_2_dec_uops_0_dst_rtype,
  input  [1:0]  io_enq_2_dec_uops_0_lrs1_rtype,
  input  [1:0]  io_enq_2_dec_uops_0_lrs2_rtype,
  input         io_enq_2_dec_uops_0_frs3_en,
  input         io_enq_2_dec_uops_0_fp_val,
  input         io_enq_2_dec_uops_0_fp_single,
  input         io_enq_2_dec_uops_0_xcpt_pf_if,
  input         io_enq_2_dec_uops_0_xcpt_ae_if,
  input         io_enq_2_dec_uops_0_xcpt_ma_if,
  input         io_enq_2_dec_uops_0_bp_debug_if,
  input         io_enq_2_dec_uops_0_bp_xcpt_if,
  input  [1:0]  io_enq_2_dec_uops_0_debug_fsrc,
  input  [1:0]  io_enq_2_dec_uops_0_debug_tsrc,
  input         io_enq_2_dec_uops_1_switch,
  input         io_enq_2_dec_uops_1_switch_off,
  input         io_enq_2_dec_uops_1_is_unicore,
  input  [2:0]  io_enq_2_dec_uops_1_shift,
  input  [1:0]  io_enq_2_dec_uops_1_lrs3_rtype,
  input         io_enq_2_dec_uops_1_rflag,
  input         io_enq_2_dec_uops_1_wflag,
  input  [3:0]  io_enq_2_dec_uops_1_prflag,
  input  [3:0]  io_enq_2_dec_uops_1_pwflag,
  input         io_enq_2_dec_uops_1_pflag_busy,
  input  [3:0]  io_enq_2_dec_uops_1_stale_pflag,
  input  [3:0]  io_enq_2_dec_uops_1_op1_sel,
  input  [3:0]  io_enq_2_dec_uops_1_op2_sel,
  input  [5:0]  io_enq_2_dec_uops_1_split_num,
  input  [5:0]  io_enq_2_dec_uops_1_self_index,
  input  [5:0]  io_enq_2_dec_uops_1_rob_inst_idx,
  input  [5:0]  io_enq_2_dec_uops_1_address_num,
  input  [6:0]  io_enq_2_dec_uops_1_uopc,
  input  [31:0] io_enq_2_dec_uops_1_inst,
  input  [31:0] io_enq_2_dec_uops_1_debug_inst,
  input         io_enq_2_dec_uops_1_is_rvc,
  input  [39:0] io_enq_2_dec_uops_1_debug_pc,
  input  [2:0]  io_enq_2_dec_uops_1_iq_type,
  input  [9:0]  io_enq_2_dec_uops_1_fu_code,
  input  [3:0]  io_enq_2_dec_uops_1_ctrl_br_type,
  input  [1:0]  io_enq_2_dec_uops_1_ctrl_op1_sel,
  input  [2:0]  io_enq_2_dec_uops_1_ctrl_op2_sel,
  input  [2:0]  io_enq_2_dec_uops_1_ctrl_imm_sel,
  input  [3:0]  io_enq_2_dec_uops_1_ctrl_op_fcn,
  input         io_enq_2_dec_uops_1_ctrl_fcn_dw,
  input  [2:0]  io_enq_2_dec_uops_1_ctrl_csr_cmd,
  input         io_enq_2_dec_uops_1_ctrl_is_load,
  input         io_enq_2_dec_uops_1_ctrl_is_sta,
  input         io_enq_2_dec_uops_1_ctrl_is_std,
  input  [1:0]  io_enq_2_dec_uops_1_ctrl_op3_sel,
  input  [1:0]  io_enq_2_dec_uops_1_iw_state,
  input         io_enq_2_dec_uops_1_iw_p1_poisoned,
  input         io_enq_2_dec_uops_1_iw_p2_poisoned,
  input         io_enq_2_dec_uops_1_is_br,
  input         io_enq_2_dec_uops_1_is_jalr,
  input         io_enq_2_dec_uops_1_is_jal,
  input         io_enq_2_dec_uops_1_is_sfb,
  input  [11:0] io_enq_2_dec_uops_1_br_mask,
  input  [3:0]  io_enq_2_dec_uops_1_br_tag,
  input  [4:0]  io_enq_2_dec_uops_1_ftq_idx,
  input         io_enq_2_dec_uops_1_edge_inst,
  input  [5:0]  io_enq_2_dec_uops_1_pc_lob,
  input         io_enq_2_dec_uops_1_taken,
  input  [19:0] io_enq_2_dec_uops_1_imm_packed,
  input  [11:0] io_enq_2_dec_uops_1_csr_addr,
  input  [5:0]  io_enq_2_dec_uops_1_rob_idx,
  input  [4:0]  io_enq_2_dec_uops_1_ldq_idx,
  input  [4:0]  io_enq_2_dec_uops_1_stq_idx,
  input  [1:0]  io_enq_2_dec_uops_1_rxq_idx,
  input  [6:0]  io_enq_2_dec_uops_1_pdst,
  input  [6:0]  io_enq_2_dec_uops_1_prs1,
  input  [6:0]  io_enq_2_dec_uops_1_prs2,
  input  [6:0]  io_enq_2_dec_uops_1_prs3,
  input  [4:0]  io_enq_2_dec_uops_1_ppred,
  input         io_enq_2_dec_uops_1_prs1_busy,
  input         io_enq_2_dec_uops_1_prs2_busy,
  input         io_enq_2_dec_uops_1_prs3_busy,
  input         io_enq_2_dec_uops_1_ppred_busy,
  input  [6:0]  io_enq_2_dec_uops_1_stale_pdst,
  input         io_enq_2_dec_uops_1_exception,
  input  [63:0] io_enq_2_dec_uops_1_exc_cause,
  input         io_enq_2_dec_uops_1_bypassable,
  input  [4:0]  io_enq_2_dec_uops_1_mem_cmd,
  input  [1:0]  io_enq_2_dec_uops_1_mem_size,
  input         io_enq_2_dec_uops_1_mem_signed,
  input         io_enq_2_dec_uops_1_is_fence,
  input         io_enq_2_dec_uops_1_is_fencei,
  input         io_enq_2_dec_uops_1_is_amo,
  input         io_enq_2_dec_uops_1_uses_ldq,
  input         io_enq_2_dec_uops_1_uses_stq,
  input         io_enq_2_dec_uops_1_is_sys_pc2epc,
  input         io_enq_2_dec_uops_1_is_unique,
  input         io_enq_2_dec_uops_1_flush_on_commit,
  input         io_enq_2_dec_uops_1_ldst_is_rs1,
  input  [5:0]  io_enq_2_dec_uops_1_ldst,
  input  [5:0]  io_enq_2_dec_uops_1_lrs1,
  input  [5:0]  io_enq_2_dec_uops_1_lrs2,
  input  [5:0]  io_enq_2_dec_uops_1_lrs3,
  input         io_enq_2_dec_uops_1_ldst_val,
  input  [1:0]  io_enq_2_dec_uops_1_dst_rtype,
  input  [1:0]  io_enq_2_dec_uops_1_lrs1_rtype,
  input  [1:0]  io_enq_2_dec_uops_1_lrs2_rtype,
  input         io_enq_2_dec_uops_1_frs3_en,
  input         io_enq_2_dec_uops_1_fp_val,
  input         io_enq_2_dec_uops_1_fp_single,
  input         io_enq_2_dec_uops_1_xcpt_pf_if,
  input         io_enq_2_dec_uops_1_xcpt_ae_if,
  input         io_enq_2_dec_uops_1_xcpt_ma_if,
  input         io_enq_2_dec_uops_1_bp_debug_if,
  input         io_enq_2_dec_uops_1_bp_xcpt_if,
  input  [1:0]  io_enq_2_dec_uops_1_debug_fsrc,
  input  [1:0]  io_enq_2_dec_uops_1_debug_tsrc,
  input         io_enq_2_dec_uops_2_switch,
  input         io_enq_2_dec_uops_2_switch_off,
  input         io_enq_2_dec_uops_2_is_unicore,
  input  [2:0]  io_enq_2_dec_uops_2_shift,
  input  [1:0]  io_enq_2_dec_uops_2_lrs3_rtype,
  input         io_enq_2_dec_uops_2_rflag,
  input         io_enq_2_dec_uops_2_wflag,
  input  [3:0]  io_enq_2_dec_uops_2_prflag,
  input  [3:0]  io_enq_2_dec_uops_2_pwflag,
  input         io_enq_2_dec_uops_2_pflag_busy,
  input  [3:0]  io_enq_2_dec_uops_2_stale_pflag,
  input  [3:0]  io_enq_2_dec_uops_2_op1_sel,
  input  [3:0]  io_enq_2_dec_uops_2_op2_sel,
  input  [5:0]  io_enq_2_dec_uops_2_split_num,
  input  [5:0]  io_enq_2_dec_uops_2_self_index,
  input  [5:0]  io_enq_2_dec_uops_2_rob_inst_idx,
  input  [5:0]  io_enq_2_dec_uops_2_address_num,
  input  [6:0]  io_enq_2_dec_uops_2_uopc,
  input  [31:0] io_enq_2_dec_uops_2_inst,
  input  [31:0] io_enq_2_dec_uops_2_debug_inst,
  input         io_enq_2_dec_uops_2_is_rvc,
  input  [39:0] io_enq_2_dec_uops_2_debug_pc,
  input  [2:0]  io_enq_2_dec_uops_2_iq_type,
  input  [9:0]  io_enq_2_dec_uops_2_fu_code,
  input  [3:0]  io_enq_2_dec_uops_2_ctrl_br_type,
  input  [1:0]  io_enq_2_dec_uops_2_ctrl_op1_sel,
  input  [2:0]  io_enq_2_dec_uops_2_ctrl_op2_sel,
  input  [2:0]  io_enq_2_dec_uops_2_ctrl_imm_sel,
  input  [3:0]  io_enq_2_dec_uops_2_ctrl_op_fcn,
  input         io_enq_2_dec_uops_2_ctrl_fcn_dw,
  input  [2:0]  io_enq_2_dec_uops_2_ctrl_csr_cmd,
  input         io_enq_2_dec_uops_2_ctrl_is_load,
  input         io_enq_2_dec_uops_2_ctrl_is_sta,
  input         io_enq_2_dec_uops_2_ctrl_is_std,
  input  [1:0]  io_enq_2_dec_uops_2_ctrl_op3_sel,
  input  [1:0]  io_enq_2_dec_uops_2_iw_state,
  input         io_enq_2_dec_uops_2_iw_p1_poisoned,
  input         io_enq_2_dec_uops_2_iw_p2_poisoned,
  input         io_enq_2_dec_uops_2_is_br,
  input         io_enq_2_dec_uops_2_is_jalr,
  input         io_enq_2_dec_uops_2_is_jal,
  input         io_enq_2_dec_uops_2_is_sfb,
  input  [11:0] io_enq_2_dec_uops_2_br_mask,
  input  [3:0]  io_enq_2_dec_uops_2_br_tag,
  input  [4:0]  io_enq_2_dec_uops_2_ftq_idx,
  input         io_enq_2_dec_uops_2_edge_inst,
  input  [5:0]  io_enq_2_dec_uops_2_pc_lob,
  input         io_enq_2_dec_uops_2_taken,
  input  [19:0] io_enq_2_dec_uops_2_imm_packed,
  input  [11:0] io_enq_2_dec_uops_2_csr_addr,
  input  [5:0]  io_enq_2_dec_uops_2_rob_idx,
  input  [4:0]  io_enq_2_dec_uops_2_ldq_idx,
  input  [4:0]  io_enq_2_dec_uops_2_stq_idx,
  input  [1:0]  io_enq_2_dec_uops_2_rxq_idx,
  input  [6:0]  io_enq_2_dec_uops_2_pdst,
  input  [6:0]  io_enq_2_dec_uops_2_prs1,
  input  [6:0]  io_enq_2_dec_uops_2_prs2,
  input  [6:0]  io_enq_2_dec_uops_2_prs3,
  input  [4:0]  io_enq_2_dec_uops_2_ppred,
  input         io_enq_2_dec_uops_2_prs1_busy,
  input         io_enq_2_dec_uops_2_prs2_busy,
  input         io_enq_2_dec_uops_2_prs3_busy,
  input         io_enq_2_dec_uops_2_ppred_busy,
  input  [6:0]  io_enq_2_dec_uops_2_stale_pdst,
  input         io_enq_2_dec_uops_2_exception,
  input  [63:0] io_enq_2_dec_uops_2_exc_cause,
  input         io_enq_2_dec_uops_2_bypassable,
  input  [4:0]  io_enq_2_dec_uops_2_mem_cmd,
  input  [1:0]  io_enq_2_dec_uops_2_mem_size,
  input         io_enq_2_dec_uops_2_mem_signed,
  input         io_enq_2_dec_uops_2_is_fence,
  input         io_enq_2_dec_uops_2_is_fencei,
  input         io_enq_2_dec_uops_2_is_amo,
  input         io_enq_2_dec_uops_2_uses_ldq,
  input         io_enq_2_dec_uops_2_uses_stq,
  input         io_enq_2_dec_uops_2_is_sys_pc2epc,
  input         io_enq_2_dec_uops_2_is_unique,
  input         io_enq_2_dec_uops_2_flush_on_commit,
  input         io_enq_2_dec_uops_2_ldst_is_rs1,
  input  [5:0]  io_enq_2_dec_uops_2_ldst,
  input  [5:0]  io_enq_2_dec_uops_2_lrs1,
  input  [5:0]  io_enq_2_dec_uops_2_lrs2,
  input  [5:0]  io_enq_2_dec_uops_2_lrs3,
  input         io_enq_2_dec_uops_2_ldst_val,
  input  [1:0]  io_enq_2_dec_uops_2_dst_rtype,
  input  [1:0]  io_enq_2_dec_uops_2_lrs1_rtype,
  input  [1:0]  io_enq_2_dec_uops_2_lrs2_rtype,
  input         io_enq_2_dec_uops_2_frs3_en,
  input         io_enq_2_dec_uops_2_fp_val,
  input         io_enq_2_dec_uops_2_fp_single,
  input         io_enq_2_dec_uops_2_xcpt_pf_if,
  input         io_enq_2_dec_uops_2_xcpt_ae_if,
  input         io_enq_2_dec_uops_2_xcpt_ma_if,
  input         io_enq_2_dec_uops_2_bp_debug_if,
  input         io_enq_2_dec_uops_2_bp_xcpt_if,
  input  [1:0]  io_enq_2_dec_uops_2_debug_fsrc,
  input  [1:0]  io_enq_2_dec_uops_2_debug_tsrc,
  input         io_enq_2_dec_uops_3_switch,
  input         io_enq_2_dec_uops_3_switch_off,
  input         io_enq_2_dec_uops_3_is_unicore,
  input  [2:0]  io_enq_2_dec_uops_3_shift,
  input  [1:0]  io_enq_2_dec_uops_3_lrs3_rtype,
  input         io_enq_2_dec_uops_3_rflag,
  input         io_enq_2_dec_uops_3_wflag,
  input  [3:0]  io_enq_2_dec_uops_3_prflag,
  input  [3:0]  io_enq_2_dec_uops_3_pwflag,
  input         io_enq_2_dec_uops_3_pflag_busy,
  input  [3:0]  io_enq_2_dec_uops_3_stale_pflag,
  input  [3:0]  io_enq_2_dec_uops_3_op1_sel,
  input  [3:0]  io_enq_2_dec_uops_3_op2_sel,
  input  [5:0]  io_enq_2_dec_uops_3_split_num,
  input  [5:0]  io_enq_2_dec_uops_3_self_index,
  input  [5:0]  io_enq_2_dec_uops_3_rob_inst_idx,
  input  [5:0]  io_enq_2_dec_uops_3_address_num,
  input  [6:0]  io_enq_2_dec_uops_3_uopc,
  input  [31:0] io_enq_2_dec_uops_3_inst,
  input  [31:0] io_enq_2_dec_uops_3_debug_inst,
  input         io_enq_2_dec_uops_3_is_rvc,
  input  [39:0] io_enq_2_dec_uops_3_debug_pc,
  input  [2:0]  io_enq_2_dec_uops_3_iq_type,
  input  [9:0]  io_enq_2_dec_uops_3_fu_code,
  input  [3:0]  io_enq_2_dec_uops_3_ctrl_br_type,
  input  [1:0]  io_enq_2_dec_uops_3_ctrl_op1_sel,
  input  [2:0]  io_enq_2_dec_uops_3_ctrl_op2_sel,
  input  [2:0]  io_enq_2_dec_uops_3_ctrl_imm_sel,
  input  [3:0]  io_enq_2_dec_uops_3_ctrl_op_fcn,
  input         io_enq_2_dec_uops_3_ctrl_fcn_dw,
  input  [2:0]  io_enq_2_dec_uops_3_ctrl_csr_cmd,
  input         io_enq_2_dec_uops_3_ctrl_is_load,
  input         io_enq_2_dec_uops_3_ctrl_is_sta,
  input         io_enq_2_dec_uops_3_ctrl_is_std,
  input  [1:0]  io_enq_2_dec_uops_3_ctrl_op3_sel,
  input  [1:0]  io_enq_2_dec_uops_3_iw_state,
  input         io_enq_2_dec_uops_3_iw_p1_poisoned,
  input         io_enq_2_dec_uops_3_iw_p2_poisoned,
  input         io_enq_2_dec_uops_3_is_br,
  input         io_enq_2_dec_uops_3_is_jalr,
  input         io_enq_2_dec_uops_3_is_jal,
  input         io_enq_2_dec_uops_3_is_sfb,
  input  [11:0] io_enq_2_dec_uops_3_br_mask,
  input  [3:0]  io_enq_2_dec_uops_3_br_tag,
  input  [4:0]  io_enq_2_dec_uops_3_ftq_idx,
  input         io_enq_2_dec_uops_3_edge_inst,
  input  [5:0]  io_enq_2_dec_uops_3_pc_lob,
  input         io_enq_2_dec_uops_3_taken,
  input  [19:0] io_enq_2_dec_uops_3_imm_packed,
  input  [11:0] io_enq_2_dec_uops_3_csr_addr,
  input  [5:0]  io_enq_2_dec_uops_3_rob_idx,
  input  [4:0]  io_enq_2_dec_uops_3_ldq_idx,
  input  [4:0]  io_enq_2_dec_uops_3_stq_idx,
  input  [1:0]  io_enq_2_dec_uops_3_rxq_idx,
  input  [6:0]  io_enq_2_dec_uops_3_pdst,
  input  [6:0]  io_enq_2_dec_uops_3_prs1,
  input  [6:0]  io_enq_2_dec_uops_3_prs2,
  input  [6:0]  io_enq_2_dec_uops_3_prs3,
  input  [4:0]  io_enq_2_dec_uops_3_ppred,
  input         io_enq_2_dec_uops_3_prs1_busy,
  input         io_enq_2_dec_uops_3_prs2_busy,
  input         io_enq_2_dec_uops_3_prs3_busy,
  input         io_enq_2_dec_uops_3_ppred_busy,
  input  [6:0]  io_enq_2_dec_uops_3_stale_pdst,
  input         io_enq_2_dec_uops_3_exception,
  input  [63:0] io_enq_2_dec_uops_3_exc_cause,
  input         io_enq_2_dec_uops_3_bypassable,
  input  [4:0]  io_enq_2_dec_uops_3_mem_cmd,
  input  [1:0]  io_enq_2_dec_uops_3_mem_size,
  input         io_enq_2_dec_uops_3_mem_signed,
  input         io_enq_2_dec_uops_3_is_fence,
  input         io_enq_2_dec_uops_3_is_fencei,
  input         io_enq_2_dec_uops_3_is_amo,
  input         io_enq_2_dec_uops_3_uses_ldq,
  input         io_enq_2_dec_uops_3_uses_stq,
  input         io_enq_2_dec_uops_3_is_sys_pc2epc,
  input         io_enq_2_dec_uops_3_is_unique,
  input         io_enq_2_dec_uops_3_flush_on_commit,
  input         io_enq_2_dec_uops_3_ldst_is_rs1,
  input  [5:0]  io_enq_2_dec_uops_3_ldst,
  input  [5:0]  io_enq_2_dec_uops_3_lrs1,
  input  [5:0]  io_enq_2_dec_uops_3_lrs2,
  input  [5:0]  io_enq_2_dec_uops_3_lrs3,
  input         io_enq_2_dec_uops_3_ldst_val,
  input  [1:0]  io_enq_2_dec_uops_3_dst_rtype,
  input  [1:0]  io_enq_2_dec_uops_3_lrs1_rtype,
  input  [1:0]  io_enq_2_dec_uops_3_lrs2_rtype,
  input         io_enq_2_dec_uops_3_frs3_en,
  input         io_enq_2_dec_uops_3_fp_val,
  input         io_enq_2_dec_uops_3_fp_single,
  input         io_enq_2_dec_uops_3_xcpt_pf_if,
  input         io_enq_2_dec_uops_3_xcpt_ae_if,
  input         io_enq_2_dec_uops_3_xcpt_ma_if,
  input         io_enq_2_dec_uops_3_bp_debug_if,
  input         io_enq_2_dec_uops_3_bp_xcpt_if,
  input  [1:0]  io_enq_2_dec_uops_3_debug_fsrc,
  input  [1:0]  io_enq_2_dec_uops_3_debug_tsrc,
  input         io_enq_2_val_mask_0,
  input         io_enq_2_val_mask_1,
  input         io_enq_2_val_mask_2,
  input         io_enq_2_val_mask_3,
  input         io_enq_3_dec_uops_0_switch,
  input         io_enq_3_dec_uops_0_switch_off,
  input         io_enq_3_dec_uops_0_is_unicore,
  input  [2:0]  io_enq_3_dec_uops_0_shift,
  input  [1:0]  io_enq_3_dec_uops_0_lrs3_rtype,
  input         io_enq_3_dec_uops_0_rflag,
  input         io_enq_3_dec_uops_0_wflag,
  input  [3:0]  io_enq_3_dec_uops_0_prflag,
  input  [3:0]  io_enq_3_dec_uops_0_pwflag,
  input         io_enq_3_dec_uops_0_pflag_busy,
  input  [3:0]  io_enq_3_dec_uops_0_stale_pflag,
  input  [3:0]  io_enq_3_dec_uops_0_op1_sel,
  input  [3:0]  io_enq_3_dec_uops_0_op2_sel,
  input  [5:0]  io_enq_3_dec_uops_0_split_num,
  input  [5:0]  io_enq_3_dec_uops_0_self_index,
  input  [5:0]  io_enq_3_dec_uops_0_rob_inst_idx,
  input  [5:0]  io_enq_3_dec_uops_0_address_num,
  input  [6:0]  io_enq_3_dec_uops_0_uopc,
  input  [31:0] io_enq_3_dec_uops_0_inst,
  input  [31:0] io_enq_3_dec_uops_0_debug_inst,
  input         io_enq_3_dec_uops_0_is_rvc,
  input  [39:0] io_enq_3_dec_uops_0_debug_pc,
  input  [2:0]  io_enq_3_dec_uops_0_iq_type,
  input  [9:0]  io_enq_3_dec_uops_0_fu_code,
  input  [3:0]  io_enq_3_dec_uops_0_ctrl_br_type,
  input  [1:0]  io_enq_3_dec_uops_0_ctrl_op1_sel,
  input  [2:0]  io_enq_3_dec_uops_0_ctrl_op2_sel,
  input  [2:0]  io_enq_3_dec_uops_0_ctrl_imm_sel,
  input  [3:0]  io_enq_3_dec_uops_0_ctrl_op_fcn,
  input         io_enq_3_dec_uops_0_ctrl_fcn_dw,
  input  [2:0]  io_enq_3_dec_uops_0_ctrl_csr_cmd,
  input         io_enq_3_dec_uops_0_ctrl_is_load,
  input         io_enq_3_dec_uops_0_ctrl_is_sta,
  input         io_enq_3_dec_uops_0_ctrl_is_std,
  input  [1:0]  io_enq_3_dec_uops_0_ctrl_op3_sel,
  input  [1:0]  io_enq_3_dec_uops_0_iw_state,
  input         io_enq_3_dec_uops_0_iw_p1_poisoned,
  input         io_enq_3_dec_uops_0_iw_p2_poisoned,
  input         io_enq_3_dec_uops_0_is_br,
  input         io_enq_3_dec_uops_0_is_jalr,
  input         io_enq_3_dec_uops_0_is_jal,
  input         io_enq_3_dec_uops_0_is_sfb,
  input  [11:0] io_enq_3_dec_uops_0_br_mask,
  input  [3:0]  io_enq_3_dec_uops_0_br_tag,
  input  [4:0]  io_enq_3_dec_uops_0_ftq_idx,
  input         io_enq_3_dec_uops_0_edge_inst,
  input  [5:0]  io_enq_3_dec_uops_0_pc_lob,
  input         io_enq_3_dec_uops_0_taken,
  input  [19:0] io_enq_3_dec_uops_0_imm_packed,
  input  [11:0] io_enq_3_dec_uops_0_csr_addr,
  input  [5:0]  io_enq_3_dec_uops_0_rob_idx,
  input  [4:0]  io_enq_3_dec_uops_0_ldq_idx,
  input  [4:0]  io_enq_3_dec_uops_0_stq_idx,
  input  [1:0]  io_enq_3_dec_uops_0_rxq_idx,
  input  [6:0]  io_enq_3_dec_uops_0_pdst,
  input  [6:0]  io_enq_3_dec_uops_0_prs1,
  input  [6:0]  io_enq_3_dec_uops_0_prs2,
  input  [6:0]  io_enq_3_dec_uops_0_prs3,
  input  [4:0]  io_enq_3_dec_uops_0_ppred,
  input         io_enq_3_dec_uops_0_prs1_busy,
  input         io_enq_3_dec_uops_0_prs2_busy,
  input         io_enq_3_dec_uops_0_prs3_busy,
  input         io_enq_3_dec_uops_0_ppred_busy,
  input  [6:0]  io_enq_3_dec_uops_0_stale_pdst,
  input         io_enq_3_dec_uops_0_exception,
  input  [63:0] io_enq_3_dec_uops_0_exc_cause,
  input         io_enq_3_dec_uops_0_bypassable,
  input  [4:0]  io_enq_3_dec_uops_0_mem_cmd,
  input  [1:0]  io_enq_3_dec_uops_0_mem_size,
  input         io_enq_3_dec_uops_0_mem_signed,
  input         io_enq_3_dec_uops_0_is_fence,
  input         io_enq_3_dec_uops_0_is_fencei,
  input         io_enq_3_dec_uops_0_is_amo,
  input         io_enq_3_dec_uops_0_uses_ldq,
  input         io_enq_3_dec_uops_0_uses_stq,
  input         io_enq_3_dec_uops_0_is_sys_pc2epc,
  input         io_enq_3_dec_uops_0_is_unique,
  input         io_enq_3_dec_uops_0_flush_on_commit,
  input         io_enq_3_dec_uops_0_ldst_is_rs1,
  input  [5:0]  io_enq_3_dec_uops_0_ldst,
  input  [5:0]  io_enq_3_dec_uops_0_lrs1,
  input  [5:0]  io_enq_3_dec_uops_0_lrs2,
  input  [5:0]  io_enq_3_dec_uops_0_lrs3,
  input         io_enq_3_dec_uops_0_ldst_val,
  input  [1:0]  io_enq_3_dec_uops_0_dst_rtype,
  input  [1:0]  io_enq_3_dec_uops_0_lrs1_rtype,
  input  [1:0]  io_enq_3_dec_uops_0_lrs2_rtype,
  input         io_enq_3_dec_uops_0_frs3_en,
  input         io_enq_3_dec_uops_0_fp_val,
  input         io_enq_3_dec_uops_0_fp_single,
  input         io_enq_3_dec_uops_0_xcpt_pf_if,
  input         io_enq_3_dec_uops_0_xcpt_ae_if,
  input         io_enq_3_dec_uops_0_xcpt_ma_if,
  input         io_enq_3_dec_uops_0_bp_debug_if,
  input         io_enq_3_dec_uops_0_bp_xcpt_if,
  input  [1:0]  io_enq_3_dec_uops_0_debug_fsrc,
  input  [1:0]  io_enq_3_dec_uops_0_debug_tsrc,
  input         io_enq_3_dec_uops_1_switch,
  input         io_enq_3_dec_uops_1_switch_off,
  input         io_enq_3_dec_uops_1_is_unicore,
  input  [2:0]  io_enq_3_dec_uops_1_shift,
  input  [1:0]  io_enq_3_dec_uops_1_lrs3_rtype,
  input         io_enq_3_dec_uops_1_rflag,
  input         io_enq_3_dec_uops_1_wflag,
  input  [3:0]  io_enq_3_dec_uops_1_prflag,
  input  [3:0]  io_enq_3_dec_uops_1_pwflag,
  input         io_enq_3_dec_uops_1_pflag_busy,
  input  [3:0]  io_enq_3_dec_uops_1_stale_pflag,
  input  [3:0]  io_enq_3_dec_uops_1_op1_sel,
  input  [3:0]  io_enq_3_dec_uops_1_op2_sel,
  input  [5:0]  io_enq_3_dec_uops_1_split_num,
  input  [5:0]  io_enq_3_dec_uops_1_self_index,
  input  [5:0]  io_enq_3_dec_uops_1_rob_inst_idx,
  input  [5:0]  io_enq_3_dec_uops_1_address_num,
  input  [6:0]  io_enq_3_dec_uops_1_uopc,
  input  [31:0] io_enq_3_dec_uops_1_inst,
  input  [31:0] io_enq_3_dec_uops_1_debug_inst,
  input         io_enq_3_dec_uops_1_is_rvc,
  input  [39:0] io_enq_3_dec_uops_1_debug_pc,
  input  [2:0]  io_enq_3_dec_uops_1_iq_type,
  input  [9:0]  io_enq_3_dec_uops_1_fu_code,
  input  [3:0]  io_enq_3_dec_uops_1_ctrl_br_type,
  input  [1:0]  io_enq_3_dec_uops_1_ctrl_op1_sel,
  input  [2:0]  io_enq_3_dec_uops_1_ctrl_op2_sel,
  input  [2:0]  io_enq_3_dec_uops_1_ctrl_imm_sel,
  input  [3:0]  io_enq_3_dec_uops_1_ctrl_op_fcn,
  input         io_enq_3_dec_uops_1_ctrl_fcn_dw,
  input  [2:0]  io_enq_3_dec_uops_1_ctrl_csr_cmd,
  input         io_enq_3_dec_uops_1_ctrl_is_load,
  input         io_enq_3_dec_uops_1_ctrl_is_sta,
  input         io_enq_3_dec_uops_1_ctrl_is_std,
  input  [1:0]  io_enq_3_dec_uops_1_ctrl_op3_sel,
  input  [1:0]  io_enq_3_dec_uops_1_iw_state,
  input         io_enq_3_dec_uops_1_iw_p1_poisoned,
  input         io_enq_3_dec_uops_1_iw_p2_poisoned,
  input         io_enq_3_dec_uops_1_is_br,
  input         io_enq_3_dec_uops_1_is_jalr,
  input         io_enq_3_dec_uops_1_is_jal,
  input         io_enq_3_dec_uops_1_is_sfb,
  input  [11:0] io_enq_3_dec_uops_1_br_mask,
  input  [3:0]  io_enq_3_dec_uops_1_br_tag,
  input  [4:0]  io_enq_3_dec_uops_1_ftq_idx,
  input         io_enq_3_dec_uops_1_edge_inst,
  input  [5:0]  io_enq_3_dec_uops_1_pc_lob,
  input         io_enq_3_dec_uops_1_taken,
  input  [19:0] io_enq_3_dec_uops_1_imm_packed,
  input  [11:0] io_enq_3_dec_uops_1_csr_addr,
  input  [5:0]  io_enq_3_dec_uops_1_rob_idx,
  input  [4:0]  io_enq_3_dec_uops_1_ldq_idx,
  input  [4:0]  io_enq_3_dec_uops_1_stq_idx,
  input  [1:0]  io_enq_3_dec_uops_1_rxq_idx,
  input  [6:0]  io_enq_3_dec_uops_1_pdst,
  input  [6:0]  io_enq_3_dec_uops_1_prs1,
  input  [6:0]  io_enq_3_dec_uops_1_prs2,
  input  [6:0]  io_enq_3_dec_uops_1_prs3,
  input  [4:0]  io_enq_3_dec_uops_1_ppred,
  input         io_enq_3_dec_uops_1_prs1_busy,
  input         io_enq_3_dec_uops_1_prs2_busy,
  input         io_enq_3_dec_uops_1_prs3_busy,
  input         io_enq_3_dec_uops_1_ppred_busy,
  input  [6:0]  io_enq_3_dec_uops_1_stale_pdst,
  input         io_enq_3_dec_uops_1_exception,
  input  [63:0] io_enq_3_dec_uops_1_exc_cause,
  input         io_enq_3_dec_uops_1_bypassable,
  input  [4:0]  io_enq_3_dec_uops_1_mem_cmd,
  input  [1:0]  io_enq_3_dec_uops_1_mem_size,
  input         io_enq_3_dec_uops_1_mem_signed,
  input         io_enq_3_dec_uops_1_is_fence,
  input         io_enq_3_dec_uops_1_is_fencei,
  input         io_enq_3_dec_uops_1_is_amo,
  input         io_enq_3_dec_uops_1_uses_ldq,
  input         io_enq_3_dec_uops_1_uses_stq,
  input         io_enq_3_dec_uops_1_is_sys_pc2epc,
  input         io_enq_3_dec_uops_1_is_unique,
  input         io_enq_3_dec_uops_1_flush_on_commit,
  input         io_enq_3_dec_uops_1_ldst_is_rs1,
  input  [5:0]  io_enq_3_dec_uops_1_ldst,
  input  [5:0]  io_enq_3_dec_uops_1_lrs1,
  input  [5:0]  io_enq_3_dec_uops_1_lrs2,
  input  [5:0]  io_enq_3_dec_uops_1_lrs3,
  input         io_enq_3_dec_uops_1_ldst_val,
  input  [1:0]  io_enq_3_dec_uops_1_dst_rtype,
  input  [1:0]  io_enq_3_dec_uops_1_lrs1_rtype,
  input  [1:0]  io_enq_3_dec_uops_1_lrs2_rtype,
  input         io_enq_3_dec_uops_1_frs3_en,
  input         io_enq_3_dec_uops_1_fp_val,
  input         io_enq_3_dec_uops_1_fp_single,
  input         io_enq_3_dec_uops_1_xcpt_pf_if,
  input         io_enq_3_dec_uops_1_xcpt_ae_if,
  input         io_enq_3_dec_uops_1_xcpt_ma_if,
  input         io_enq_3_dec_uops_1_bp_debug_if,
  input         io_enq_3_dec_uops_1_bp_xcpt_if,
  input  [1:0]  io_enq_3_dec_uops_1_debug_fsrc,
  input  [1:0]  io_enq_3_dec_uops_1_debug_tsrc,
  input         io_enq_3_dec_uops_2_switch,
  input         io_enq_3_dec_uops_2_switch_off,
  input         io_enq_3_dec_uops_2_is_unicore,
  input  [2:0]  io_enq_3_dec_uops_2_shift,
  input  [1:0]  io_enq_3_dec_uops_2_lrs3_rtype,
  input         io_enq_3_dec_uops_2_rflag,
  input         io_enq_3_dec_uops_2_wflag,
  input  [3:0]  io_enq_3_dec_uops_2_prflag,
  input  [3:0]  io_enq_3_dec_uops_2_pwflag,
  input         io_enq_3_dec_uops_2_pflag_busy,
  input  [3:0]  io_enq_3_dec_uops_2_stale_pflag,
  input  [3:0]  io_enq_3_dec_uops_2_op1_sel,
  input  [3:0]  io_enq_3_dec_uops_2_op2_sel,
  input  [5:0]  io_enq_3_dec_uops_2_split_num,
  input  [5:0]  io_enq_3_dec_uops_2_self_index,
  input  [5:0]  io_enq_3_dec_uops_2_rob_inst_idx,
  input  [5:0]  io_enq_3_dec_uops_2_address_num,
  input  [6:0]  io_enq_3_dec_uops_2_uopc,
  input  [31:0] io_enq_3_dec_uops_2_inst,
  input  [31:0] io_enq_3_dec_uops_2_debug_inst,
  input         io_enq_3_dec_uops_2_is_rvc,
  input  [39:0] io_enq_3_dec_uops_2_debug_pc,
  input  [2:0]  io_enq_3_dec_uops_2_iq_type,
  input  [9:0]  io_enq_3_dec_uops_2_fu_code,
  input  [3:0]  io_enq_3_dec_uops_2_ctrl_br_type,
  input  [1:0]  io_enq_3_dec_uops_2_ctrl_op1_sel,
  input  [2:0]  io_enq_3_dec_uops_2_ctrl_op2_sel,
  input  [2:0]  io_enq_3_dec_uops_2_ctrl_imm_sel,
  input  [3:0]  io_enq_3_dec_uops_2_ctrl_op_fcn,
  input         io_enq_3_dec_uops_2_ctrl_fcn_dw,
  input  [2:0]  io_enq_3_dec_uops_2_ctrl_csr_cmd,
  input         io_enq_3_dec_uops_2_ctrl_is_load,
  input         io_enq_3_dec_uops_2_ctrl_is_sta,
  input         io_enq_3_dec_uops_2_ctrl_is_std,
  input  [1:0]  io_enq_3_dec_uops_2_ctrl_op3_sel,
  input  [1:0]  io_enq_3_dec_uops_2_iw_state,
  input         io_enq_3_dec_uops_2_iw_p1_poisoned,
  input         io_enq_3_dec_uops_2_iw_p2_poisoned,
  input         io_enq_3_dec_uops_2_is_br,
  input         io_enq_3_dec_uops_2_is_jalr,
  input         io_enq_3_dec_uops_2_is_jal,
  input         io_enq_3_dec_uops_2_is_sfb,
  input  [11:0] io_enq_3_dec_uops_2_br_mask,
  input  [3:0]  io_enq_3_dec_uops_2_br_tag,
  input  [4:0]  io_enq_3_dec_uops_2_ftq_idx,
  input         io_enq_3_dec_uops_2_edge_inst,
  input  [5:0]  io_enq_3_dec_uops_2_pc_lob,
  input         io_enq_3_dec_uops_2_taken,
  input  [19:0] io_enq_3_dec_uops_2_imm_packed,
  input  [11:0] io_enq_3_dec_uops_2_csr_addr,
  input  [5:0]  io_enq_3_dec_uops_2_rob_idx,
  input  [4:0]  io_enq_3_dec_uops_2_ldq_idx,
  input  [4:0]  io_enq_3_dec_uops_2_stq_idx,
  input  [1:0]  io_enq_3_dec_uops_2_rxq_idx,
  input  [6:0]  io_enq_3_dec_uops_2_pdst,
  input  [6:0]  io_enq_3_dec_uops_2_prs1,
  input  [6:0]  io_enq_3_dec_uops_2_prs2,
  input  [6:0]  io_enq_3_dec_uops_2_prs3,
  input  [4:0]  io_enq_3_dec_uops_2_ppred,
  input         io_enq_3_dec_uops_2_prs1_busy,
  input         io_enq_3_dec_uops_2_prs2_busy,
  input         io_enq_3_dec_uops_2_prs3_busy,
  input         io_enq_3_dec_uops_2_ppred_busy,
  input  [6:0]  io_enq_3_dec_uops_2_stale_pdst,
  input         io_enq_3_dec_uops_2_exception,
  input  [63:0] io_enq_3_dec_uops_2_exc_cause,
  input         io_enq_3_dec_uops_2_bypassable,
  input  [4:0]  io_enq_3_dec_uops_2_mem_cmd,
  input  [1:0]  io_enq_3_dec_uops_2_mem_size,
  input         io_enq_3_dec_uops_2_mem_signed,
  input         io_enq_3_dec_uops_2_is_fence,
  input         io_enq_3_dec_uops_2_is_fencei,
  input         io_enq_3_dec_uops_2_is_amo,
  input         io_enq_3_dec_uops_2_uses_ldq,
  input         io_enq_3_dec_uops_2_uses_stq,
  input         io_enq_3_dec_uops_2_is_sys_pc2epc,
  input         io_enq_3_dec_uops_2_is_unique,
  input         io_enq_3_dec_uops_2_flush_on_commit,
  input         io_enq_3_dec_uops_2_ldst_is_rs1,
  input  [5:0]  io_enq_3_dec_uops_2_ldst,
  input  [5:0]  io_enq_3_dec_uops_2_lrs1,
  input  [5:0]  io_enq_3_dec_uops_2_lrs2,
  input  [5:0]  io_enq_3_dec_uops_2_lrs3,
  input         io_enq_3_dec_uops_2_ldst_val,
  input  [1:0]  io_enq_3_dec_uops_2_dst_rtype,
  input  [1:0]  io_enq_3_dec_uops_2_lrs1_rtype,
  input  [1:0]  io_enq_3_dec_uops_2_lrs2_rtype,
  input         io_enq_3_dec_uops_2_frs3_en,
  input         io_enq_3_dec_uops_2_fp_val,
  input         io_enq_3_dec_uops_2_fp_single,
  input         io_enq_3_dec_uops_2_xcpt_pf_if,
  input         io_enq_3_dec_uops_2_xcpt_ae_if,
  input         io_enq_3_dec_uops_2_xcpt_ma_if,
  input         io_enq_3_dec_uops_2_bp_debug_if,
  input         io_enq_3_dec_uops_2_bp_xcpt_if,
  input  [1:0]  io_enq_3_dec_uops_2_debug_fsrc,
  input  [1:0]  io_enq_3_dec_uops_2_debug_tsrc,
  input         io_enq_3_dec_uops_3_switch,
  input         io_enq_3_dec_uops_3_switch_off,
  input         io_enq_3_dec_uops_3_is_unicore,
  input  [2:0]  io_enq_3_dec_uops_3_shift,
  input  [1:0]  io_enq_3_dec_uops_3_lrs3_rtype,
  input         io_enq_3_dec_uops_3_rflag,
  input         io_enq_3_dec_uops_3_wflag,
  input  [3:0]  io_enq_3_dec_uops_3_prflag,
  input  [3:0]  io_enq_3_dec_uops_3_pwflag,
  input         io_enq_3_dec_uops_3_pflag_busy,
  input  [3:0]  io_enq_3_dec_uops_3_stale_pflag,
  input  [3:0]  io_enq_3_dec_uops_3_op1_sel,
  input  [3:0]  io_enq_3_dec_uops_3_op2_sel,
  input  [5:0]  io_enq_3_dec_uops_3_split_num,
  input  [5:0]  io_enq_3_dec_uops_3_self_index,
  input  [5:0]  io_enq_3_dec_uops_3_rob_inst_idx,
  input  [5:0]  io_enq_3_dec_uops_3_address_num,
  input  [6:0]  io_enq_3_dec_uops_3_uopc,
  input  [31:0] io_enq_3_dec_uops_3_inst,
  input  [31:0] io_enq_3_dec_uops_3_debug_inst,
  input         io_enq_3_dec_uops_3_is_rvc,
  input  [39:0] io_enq_3_dec_uops_3_debug_pc,
  input  [2:0]  io_enq_3_dec_uops_3_iq_type,
  input  [9:0]  io_enq_3_dec_uops_3_fu_code,
  input  [3:0]  io_enq_3_dec_uops_3_ctrl_br_type,
  input  [1:0]  io_enq_3_dec_uops_3_ctrl_op1_sel,
  input  [2:0]  io_enq_3_dec_uops_3_ctrl_op2_sel,
  input  [2:0]  io_enq_3_dec_uops_3_ctrl_imm_sel,
  input  [3:0]  io_enq_3_dec_uops_3_ctrl_op_fcn,
  input         io_enq_3_dec_uops_3_ctrl_fcn_dw,
  input  [2:0]  io_enq_3_dec_uops_3_ctrl_csr_cmd,
  input         io_enq_3_dec_uops_3_ctrl_is_load,
  input         io_enq_3_dec_uops_3_ctrl_is_sta,
  input         io_enq_3_dec_uops_3_ctrl_is_std,
  input  [1:0]  io_enq_3_dec_uops_3_ctrl_op3_sel,
  input  [1:0]  io_enq_3_dec_uops_3_iw_state,
  input         io_enq_3_dec_uops_3_iw_p1_poisoned,
  input         io_enq_3_dec_uops_3_iw_p2_poisoned,
  input         io_enq_3_dec_uops_3_is_br,
  input         io_enq_3_dec_uops_3_is_jalr,
  input         io_enq_3_dec_uops_3_is_jal,
  input         io_enq_3_dec_uops_3_is_sfb,
  input  [11:0] io_enq_3_dec_uops_3_br_mask,
  input  [3:0]  io_enq_3_dec_uops_3_br_tag,
  input  [4:0]  io_enq_3_dec_uops_3_ftq_idx,
  input         io_enq_3_dec_uops_3_edge_inst,
  input  [5:0]  io_enq_3_dec_uops_3_pc_lob,
  input         io_enq_3_dec_uops_3_taken,
  input  [19:0] io_enq_3_dec_uops_3_imm_packed,
  input  [11:0] io_enq_3_dec_uops_3_csr_addr,
  input  [5:0]  io_enq_3_dec_uops_3_rob_idx,
  input  [4:0]  io_enq_3_dec_uops_3_ldq_idx,
  input  [4:0]  io_enq_3_dec_uops_3_stq_idx,
  input  [1:0]  io_enq_3_dec_uops_3_rxq_idx,
  input  [6:0]  io_enq_3_dec_uops_3_pdst,
  input  [6:0]  io_enq_3_dec_uops_3_prs1,
  input  [6:0]  io_enq_3_dec_uops_3_prs2,
  input  [6:0]  io_enq_3_dec_uops_3_prs3,
  input  [4:0]  io_enq_3_dec_uops_3_ppred,
  input         io_enq_3_dec_uops_3_prs1_busy,
  input         io_enq_3_dec_uops_3_prs2_busy,
  input         io_enq_3_dec_uops_3_prs3_busy,
  input         io_enq_3_dec_uops_3_ppred_busy,
  input  [6:0]  io_enq_3_dec_uops_3_stale_pdst,
  input         io_enq_3_dec_uops_3_exception,
  input  [63:0] io_enq_3_dec_uops_3_exc_cause,
  input         io_enq_3_dec_uops_3_bypassable,
  input  [4:0]  io_enq_3_dec_uops_3_mem_cmd,
  input  [1:0]  io_enq_3_dec_uops_3_mem_size,
  input         io_enq_3_dec_uops_3_mem_signed,
  input         io_enq_3_dec_uops_3_is_fence,
  input         io_enq_3_dec_uops_3_is_fencei,
  input         io_enq_3_dec_uops_3_is_amo,
  input         io_enq_3_dec_uops_3_uses_ldq,
  input         io_enq_3_dec_uops_3_uses_stq,
  input         io_enq_3_dec_uops_3_is_sys_pc2epc,
  input         io_enq_3_dec_uops_3_is_unique,
  input         io_enq_3_dec_uops_3_flush_on_commit,
  input         io_enq_3_dec_uops_3_ldst_is_rs1,
  input  [5:0]  io_enq_3_dec_uops_3_ldst,
  input  [5:0]  io_enq_3_dec_uops_3_lrs1,
  input  [5:0]  io_enq_3_dec_uops_3_lrs2,
  input  [5:0]  io_enq_3_dec_uops_3_lrs3,
  input         io_enq_3_dec_uops_3_ldst_val,
  input  [1:0]  io_enq_3_dec_uops_3_dst_rtype,
  input  [1:0]  io_enq_3_dec_uops_3_lrs1_rtype,
  input  [1:0]  io_enq_3_dec_uops_3_lrs2_rtype,
  input         io_enq_3_dec_uops_3_frs3_en,
  input         io_enq_3_dec_uops_3_fp_val,
  input         io_enq_3_dec_uops_3_fp_single,
  input         io_enq_3_dec_uops_3_xcpt_pf_if,
  input         io_enq_3_dec_uops_3_xcpt_ae_if,
  input         io_enq_3_dec_uops_3_xcpt_ma_if,
  input         io_enq_3_dec_uops_3_bp_debug_if,
  input         io_enq_3_dec_uops_3_bp_xcpt_if,
  input  [1:0]  io_enq_3_dec_uops_3_debug_fsrc,
  input  [1:0]  io_enq_3_dec_uops_3_debug_tsrc,
  input         io_enq_3_val_mask_0,
  input         io_enq_3_val_mask_1,
  input         io_enq_3_val_mask_2,
  input         io_enq_3_val_mask_3,
  input         io_enq_4_dec_uops_0_switch,
  input         io_enq_4_dec_uops_0_switch_off,
  input         io_enq_4_dec_uops_0_is_unicore,
  input  [2:0]  io_enq_4_dec_uops_0_shift,
  input  [1:0]  io_enq_4_dec_uops_0_lrs3_rtype,
  input         io_enq_4_dec_uops_0_rflag,
  input         io_enq_4_dec_uops_0_wflag,
  input  [3:0]  io_enq_4_dec_uops_0_prflag,
  input  [3:0]  io_enq_4_dec_uops_0_pwflag,
  input         io_enq_4_dec_uops_0_pflag_busy,
  input  [3:0]  io_enq_4_dec_uops_0_stale_pflag,
  input  [3:0]  io_enq_4_dec_uops_0_op1_sel,
  input  [3:0]  io_enq_4_dec_uops_0_op2_sel,
  input  [5:0]  io_enq_4_dec_uops_0_split_num,
  input  [5:0]  io_enq_4_dec_uops_0_self_index,
  input  [5:0]  io_enq_4_dec_uops_0_rob_inst_idx,
  input  [5:0]  io_enq_4_dec_uops_0_address_num,
  input  [6:0]  io_enq_4_dec_uops_0_uopc,
  input  [31:0] io_enq_4_dec_uops_0_inst,
  input  [31:0] io_enq_4_dec_uops_0_debug_inst,
  input         io_enq_4_dec_uops_0_is_rvc,
  input  [39:0] io_enq_4_dec_uops_0_debug_pc,
  input  [2:0]  io_enq_4_dec_uops_0_iq_type,
  input  [9:0]  io_enq_4_dec_uops_0_fu_code,
  input  [3:0]  io_enq_4_dec_uops_0_ctrl_br_type,
  input  [1:0]  io_enq_4_dec_uops_0_ctrl_op1_sel,
  input  [2:0]  io_enq_4_dec_uops_0_ctrl_op2_sel,
  input  [2:0]  io_enq_4_dec_uops_0_ctrl_imm_sel,
  input  [3:0]  io_enq_4_dec_uops_0_ctrl_op_fcn,
  input         io_enq_4_dec_uops_0_ctrl_fcn_dw,
  input  [2:0]  io_enq_4_dec_uops_0_ctrl_csr_cmd,
  input         io_enq_4_dec_uops_0_ctrl_is_load,
  input         io_enq_4_dec_uops_0_ctrl_is_sta,
  input         io_enq_4_dec_uops_0_ctrl_is_std,
  input  [1:0]  io_enq_4_dec_uops_0_ctrl_op3_sel,
  input  [1:0]  io_enq_4_dec_uops_0_iw_state,
  input         io_enq_4_dec_uops_0_iw_p1_poisoned,
  input         io_enq_4_dec_uops_0_iw_p2_poisoned,
  input         io_enq_4_dec_uops_0_is_br,
  input         io_enq_4_dec_uops_0_is_jalr,
  input         io_enq_4_dec_uops_0_is_jal,
  input         io_enq_4_dec_uops_0_is_sfb,
  input  [11:0] io_enq_4_dec_uops_0_br_mask,
  input  [3:0]  io_enq_4_dec_uops_0_br_tag,
  input  [4:0]  io_enq_4_dec_uops_0_ftq_idx,
  input         io_enq_4_dec_uops_0_edge_inst,
  input  [5:0]  io_enq_4_dec_uops_0_pc_lob,
  input         io_enq_4_dec_uops_0_taken,
  input  [19:0] io_enq_4_dec_uops_0_imm_packed,
  input  [11:0] io_enq_4_dec_uops_0_csr_addr,
  input  [5:0]  io_enq_4_dec_uops_0_rob_idx,
  input  [4:0]  io_enq_4_dec_uops_0_ldq_idx,
  input  [4:0]  io_enq_4_dec_uops_0_stq_idx,
  input  [1:0]  io_enq_4_dec_uops_0_rxq_idx,
  input  [6:0]  io_enq_4_dec_uops_0_pdst,
  input  [6:0]  io_enq_4_dec_uops_0_prs1,
  input  [6:0]  io_enq_4_dec_uops_0_prs2,
  input  [6:0]  io_enq_4_dec_uops_0_prs3,
  input  [4:0]  io_enq_4_dec_uops_0_ppred,
  input         io_enq_4_dec_uops_0_prs1_busy,
  input         io_enq_4_dec_uops_0_prs2_busy,
  input         io_enq_4_dec_uops_0_prs3_busy,
  input         io_enq_4_dec_uops_0_ppred_busy,
  input  [6:0]  io_enq_4_dec_uops_0_stale_pdst,
  input         io_enq_4_dec_uops_0_exception,
  input  [63:0] io_enq_4_dec_uops_0_exc_cause,
  input         io_enq_4_dec_uops_0_bypassable,
  input  [4:0]  io_enq_4_dec_uops_0_mem_cmd,
  input  [1:0]  io_enq_4_dec_uops_0_mem_size,
  input         io_enq_4_dec_uops_0_mem_signed,
  input         io_enq_4_dec_uops_0_is_fence,
  input         io_enq_4_dec_uops_0_is_fencei,
  input         io_enq_4_dec_uops_0_is_amo,
  input         io_enq_4_dec_uops_0_uses_ldq,
  input         io_enq_4_dec_uops_0_uses_stq,
  input         io_enq_4_dec_uops_0_is_sys_pc2epc,
  input         io_enq_4_dec_uops_0_is_unique,
  input         io_enq_4_dec_uops_0_flush_on_commit,
  input         io_enq_4_dec_uops_0_ldst_is_rs1,
  input  [5:0]  io_enq_4_dec_uops_0_ldst,
  input  [5:0]  io_enq_4_dec_uops_0_lrs1,
  input  [5:0]  io_enq_4_dec_uops_0_lrs2,
  input  [5:0]  io_enq_4_dec_uops_0_lrs3,
  input         io_enq_4_dec_uops_0_ldst_val,
  input  [1:0]  io_enq_4_dec_uops_0_dst_rtype,
  input  [1:0]  io_enq_4_dec_uops_0_lrs1_rtype,
  input  [1:0]  io_enq_4_dec_uops_0_lrs2_rtype,
  input         io_enq_4_dec_uops_0_frs3_en,
  input         io_enq_4_dec_uops_0_fp_val,
  input         io_enq_4_dec_uops_0_fp_single,
  input         io_enq_4_dec_uops_0_xcpt_pf_if,
  input         io_enq_4_dec_uops_0_xcpt_ae_if,
  input         io_enq_4_dec_uops_0_xcpt_ma_if,
  input         io_enq_4_dec_uops_0_bp_debug_if,
  input         io_enq_4_dec_uops_0_bp_xcpt_if,
  input  [1:0]  io_enq_4_dec_uops_0_debug_fsrc,
  input  [1:0]  io_enq_4_dec_uops_0_debug_tsrc,
  input         io_enq_4_dec_uops_1_switch,
  input         io_enq_4_dec_uops_1_switch_off,
  input         io_enq_4_dec_uops_1_is_unicore,
  input  [2:0]  io_enq_4_dec_uops_1_shift,
  input  [1:0]  io_enq_4_dec_uops_1_lrs3_rtype,
  input         io_enq_4_dec_uops_1_rflag,
  input         io_enq_4_dec_uops_1_wflag,
  input  [3:0]  io_enq_4_dec_uops_1_prflag,
  input  [3:0]  io_enq_4_dec_uops_1_pwflag,
  input         io_enq_4_dec_uops_1_pflag_busy,
  input  [3:0]  io_enq_4_dec_uops_1_stale_pflag,
  input  [3:0]  io_enq_4_dec_uops_1_op1_sel,
  input  [3:0]  io_enq_4_dec_uops_1_op2_sel,
  input  [5:0]  io_enq_4_dec_uops_1_split_num,
  input  [5:0]  io_enq_4_dec_uops_1_self_index,
  input  [5:0]  io_enq_4_dec_uops_1_rob_inst_idx,
  input  [5:0]  io_enq_4_dec_uops_1_address_num,
  input  [6:0]  io_enq_4_dec_uops_1_uopc,
  input  [31:0] io_enq_4_dec_uops_1_inst,
  input  [31:0] io_enq_4_dec_uops_1_debug_inst,
  input         io_enq_4_dec_uops_1_is_rvc,
  input  [39:0] io_enq_4_dec_uops_1_debug_pc,
  input  [2:0]  io_enq_4_dec_uops_1_iq_type,
  input  [9:0]  io_enq_4_dec_uops_1_fu_code,
  input  [3:0]  io_enq_4_dec_uops_1_ctrl_br_type,
  input  [1:0]  io_enq_4_dec_uops_1_ctrl_op1_sel,
  input  [2:0]  io_enq_4_dec_uops_1_ctrl_op2_sel,
  input  [2:0]  io_enq_4_dec_uops_1_ctrl_imm_sel,
  input  [3:0]  io_enq_4_dec_uops_1_ctrl_op_fcn,
  input         io_enq_4_dec_uops_1_ctrl_fcn_dw,
  input  [2:0]  io_enq_4_dec_uops_1_ctrl_csr_cmd,
  input         io_enq_4_dec_uops_1_ctrl_is_load,
  input         io_enq_4_dec_uops_1_ctrl_is_sta,
  input         io_enq_4_dec_uops_1_ctrl_is_std,
  input  [1:0]  io_enq_4_dec_uops_1_ctrl_op3_sel,
  input  [1:0]  io_enq_4_dec_uops_1_iw_state,
  input         io_enq_4_dec_uops_1_iw_p1_poisoned,
  input         io_enq_4_dec_uops_1_iw_p2_poisoned,
  input         io_enq_4_dec_uops_1_is_br,
  input         io_enq_4_dec_uops_1_is_jalr,
  input         io_enq_4_dec_uops_1_is_jal,
  input         io_enq_4_dec_uops_1_is_sfb,
  input  [11:0] io_enq_4_dec_uops_1_br_mask,
  input  [3:0]  io_enq_4_dec_uops_1_br_tag,
  input  [4:0]  io_enq_4_dec_uops_1_ftq_idx,
  input         io_enq_4_dec_uops_1_edge_inst,
  input  [5:0]  io_enq_4_dec_uops_1_pc_lob,
  input         io_enq_4_dec_uops_1_taken,
  input  [19:0] io_enq_4_dec_uops_1_imm_packed,
  input  [11:0] io_enq_4_dec_uops_1_csr_addr,
  input  [5:0]  io_enq_4_dec_uops_1_rob_idx,
  input  [4:0]  io_enq_4_dec_uops_1_ldq_idx,
  input  [4:0]  io_enq_4_dec_uops_1_stq_idx,
  input  [1:0]  io_enq_4_dec_uops_1_rxq_idx,
  input  [6:0]  io_enq_4_dec_uops_1_pdst,
  input  [6:0]  io_enq_4_dec_uops_1_prs1,
  input  [6:0]  io_enq_4_dec_uops_1_prs2,
  input  [6:0]  io_enq_4_dec_uops_1_prs3,
  input  [4:0]  io_enq_4_dec_uops_1_ppred,
  input         io_enq_4_dec_uops_1_prs1_busy,
  input         io_enq_4_dec_uops_1_prs2_busy,
  input         io_enq_4_dec_uops_1_prs3_busy,
  input         io_enq_4_dec_uops_1_ppred_busy,
  input  [6:0]  io_enq_4_dec_uops_1_stale_pdst,
  input         io_enq_4_dec_uops_1_exception,
  input  [63:0] io_enq_4_dec_uops_1_exc_cause,
  input         io_enq_4_dec_uops_1_bypassable,
  input  [4:0]  io_enq_4_dec_uops_1_mem_cmd,
  input  [1:0]  io_enq_4_dec_uops_1_mem_size,
  input         io_enq_4_dec_uops_1_mem_signed,
  input         io_enq_4_dec_uops_1_is_fence,
  input         io_enq_4_dec_uops_1_is_fencei,
  input         io_enq_4_dec_uops_1_is_amo,
  input         io_enq_4_dec_uops_1_uses_ldq,
  input         io_enq_4_dec_uops_1_uses_stq,
  input         io_enq_4_dec_uops_1_is_sys_pc2epc,
  input         io_enq_4_dec_uops_1_is_unique,
  input         io_enq_4_dec_uops_1_flush_on_commit,
  input         io_enq_4_dec_uops_1_ldst_is_rs1,
  input  [5:0]  io_enq_4_dec_uops_1_ldst,
  input  [5:0]  io_enq_4_dec_uops_1_lrs1,
  input  [5:0]  io_enq_4_dec_uops_1_lrs2,
  input  [5:0]  io_enq_4_dec_uops_1_lrs3,
  input         io_enq_4_dec_uops_1_ldst_val,
  input  [1:0]  io_enq_4_dec_uops_1_dst_rtype,
  input  [1:0]  io_enq_4_dec_uops_1_lrs1_rtype,
  input  [1:0]  io_enq_4_dec_uops_1_lrs2_rtype,
  input         io_enq_4_dec_uops_1_frs3_en,
  input         io_enq_4_dec_uops_1_fp_val,
  input         io_enq_4_dec_uops_1_fp_single,
  input         io_enq_4_dec_uops_1_xcpt_pf_if,
  input         io_enq_4_dec_uops_1_xcpt_ae_if,
  input         io_enq_4_dec_uops_1_xcpt_ma_if,
  input         io_enq_4_dec_uops_1_bp_debug_if,
  input         io_enq_4_dec_uops_1_bp_xcpt_if,
  input  [1:0]  io_enq_4_dec_uops_1_debug_fsrc,
  input  [1:0]  io_enq_4_dec_uops_1_debug_tsrc,
  input         io_enq_4_dec_uops_2_switch,
  input         io_enq_4_dec_uops_2_switch_off,
  input         io_enq_4_dec_uops_2_is_unicore,
  input  [2:0]  io_enq_4_dec_uops_2_shift,
  input  [1:0]  io_enq_4_dec_uops_2_lrs3_rtype,
  input         io_enq_4_dec_uops_2_rflag,
  input         io_enq_4_dec_uops_2_wflag,
  input  [3:0]  io_enq_4_dec_uops_2_prflag,
  input  [3:0]  io_enq_4_dec_uops_2_pwflag,
  input         io_enq_4_dec_uops_2_pflag_busy,
  input  [3:0]  io_enq_4_dec_uops_2_stale_pflag,
  input  [3:0]  io_enq_4_dec_uops_2_op1_sel,
  input  [3:0]  io_enq_4_dec_uops_2_op2_sel,
  input  [5:0]  io_enq_4_dec_uops_2_split_num,
  input  [5:0]  io_enq_4_dec_uops_2_self_index,
  input  [5:0]  io_enq_4_dec_uops_2_rob_inst_idx,
  input  [5:0]  io_enq_4_dec_uops_2_address_num,
  input  [6:0]  io_enq_4_dec_uops_2_uopc,
  input  [31:0] io_enq_4_dec_uops_2_inst,
  input  [31:0] io_enq_4_dec_uops_2_debug_inst,
  input         io_enq_4_dec_uops_2_is_rvc,
  input  [39:0] io_enq_4_dec_uops_2_debug_pc,
  input  [2:0]  io_enq_4_dec_uops_2_iq_type,
  input  [9:0]  io_enq_4_dec_uops_2_fu_code,
  input  [3:0]  io_enq_4_dec_uops_2_ctrl_br_type,
  input  [1:0]  io_enq_4_dec_uops_2_ctrl_op1_sel,
  input  [2:0]  io_enq_4_dec_uops_2_ctrl_op2_sel,
  input  [2:0]  io_enq_4_dec_uops_2_ctrl_imm_sel,
  input  [3:0]  io_enq_4_dec_uops_2_ctrl_op_fcn,
  input         io_enq_4_dec_uops_2_ctrl_fcn_dw,
  input  [2:0]  io_enq_4_dec_uops_2_ctrl_csr_cmd,
  input         io_enq_4_dec_uops_2_ctrl_is_load,
  input         io_enq_4_dec_uops_2_ctrl_is_sta,
  input         io_enq_4_dec_uops_2_ctrl_is_std,
  input  [1:0]  io_enq_4_dec_uops_2_ctrl_op3_sel,
  input  [1:0]  io_enq_4_dec_uops_2_iw_state,
  input         io_enq_4_dec_uops_2_iw_p1_poisoned,
  input         io_enq_4_dec_uops_2_iw_p2_poisoned,
  input         io_enq_4_dec_uops_2_is_br,
  input         io_enq_4_dec_uops_2_is_jalr,
  input         io_enq_4_dec_uops_2_is_jal,
  input         io_enq_4_dec_uops_2_is_sfb,
  input  [11:0] io_enq_4_dec_uops_2_br_mask,
  input  [3:0]  io_enq_4_dec_uops_2_br_tag,
  input  [4:0]  io_enq_4_dec_uops_2_ftq_idx,
  input         io_enq_4_dec_uops_2_edge_inst,
  input  [5:0]  io_enq_4_dec_uops_2_pc_lob,
  input         io_enq_4_dec_uops_2_taken,
  input  [19:0] io_enq_4_dec_uops_2_imm_packed,
  input  [11:0] io_enq_4_dec_uops_2_csr_addr,
  input  [5:0]  io_enq_4_dec_uops_2_rob_idx,
  input  [4:0]  io_enq_4_dec_uops_2_ldq_idx,
  input  [4:0]  io_enq_4_dec_uops_2_stq_idx,
  input  [1:0]  io_enq_4_dec_uops_2_rxq_idx,
  input  [6:0]  io_enq_4_dec_uops_2_pdst,
  input  [6:0]  io_enq_4_dec_uops_2_prs1,
  input  [6:0]  io_enq_4_dec_uops_2_prs2,
  input  [6:0]  io_enq_4_dec_uops_2_prs3,
  input  [4:0]  io_enq_4_dec_uops_2_ppred,
  input         io_enq_4_dec_uops_2_prs1_busy,
  input         io_enq_4_dec_uops_2_prs2_busy,
  input         io_enq_4_dec_uops_2_prs3_busy,
  input         io_enq_4_dec_uops_2_ppred_busy,
  input  [6:0]  io_enq_4_dec_uops_2_stale_pdst,
  input         io_enq_4_dec_uops_2_exception,
  input  [63:0] io_enq_4_dec_uops_2_exc_cause,
  input         io_enq_4_dec_uops_2_bypassable,
  input  [4:0]  io_enq_4_dec_uops_2_mem_cmd,
  input  [1:0]  io_enq_4_dec_uops_2_mem_size,
  input         io_enq_4_dec_uops_2_mem_signed,
  input         io_enq_4_dec_uops_2_is_fence,
  input         io_enq_4_dec_uops_2_is_fencei,
  input         io_enq_4_dec_uops_2_is_amo,
  input         io_enq_4_dec_uops_2_uses_ldq,
  input         io_enq_4_dec_uops_2_uses_stq,
  input         io_enq_4_dec_uops_2_is_sys_pc2epc,
  input         io_enq_4_dec_uops_2_is_unique,
  input         io_enq_4_dec_uops_2_flush_on_commit,
  input         io_enq_4_dec_uops_2_ldst_is_rs1,
  input  [5:0]  io_enq_4_dec_uops_2_ldst,
  input  [5:0]  io_enq_4_dec_uops_2_lrs1,
  input  [5:0]  io_enq_4_dec_uops_2_lrs2,
  input  [5:0]  io_enq_4_dec_uops_2_lrs3,
  input         io_enq_4_dec_uops_2_ldst_val,
  input  [1:0]  io_enq_4_dec_uops_2_dst_rtype,
  input  [1:0]  io_enq_4_dec_uops_2_lrs1_rtype,
  input  [1:0]  io_enq_4_dec_uops_2_lrs2_rtype,
  input         io_enq_4_dec_uops_2_frs3_en,
  input         io_enq_4_dec_uops_2_fp_val,
  input         io_enq_4_dec_uops_2_fp_single,
  input         io_enq_4_dec_uops_2_xcpt_pf_if,
  input         io_enq_4_dec_uops_2_xcpt_ae_if,
  input         io_enq_4_dec_uops_2_xcpt_ma_if,
  input         io_enq_4_dec_uops_2_bp_debug_if,
  input         io_enq_4_dec_uops_2_bp_xcpt_if,
  input  [1:0]  io_enq_4_dec_uops_2_debug_fsrc,
  input  [1:0]  io_enq_4_dec_uops_2_debug_tsrc,
  input         io_enq_4_dec_uops_3_switch,
  input         io_enq_4_dec_uops_3_switch_off,
  input         io_enq_4_dec_uops_3_is_unicore,
  input  [2:0]  io_enq_4_dec_uops_3_shift,
  input  [1:0]  io_enq_4_dec_uops_3_lrs3_rtype,
  input         io_enq_4_dec_uops_3_rflag,
  input         io_enq_4_dec_uops_3_wflag,
  input  [3:0]  io_enq_4_dec_uops_3_prflag,
  input  [3:0]  io_enq_4_dec_uops_3_pwflag,
  input         io_enq_4_dec_uops_3_pflag_busy,
  input  [3:0]  io_enq_4_dec_uops_3_stale_pflag,
  input  [3:0]  io_enq_4_dec_uops_3_op1_sel,
  input  [3:0]  io_enq_4_dec_uops_3_op2_sel,
  input  [5:0]  io_enq_4_dec_uops_3_split_num,
  input  [5:0]  io_enq_4_dec_uops_3_self_index,
  input  [5:0]  io_enq_4_dec_uops_3_rob_inst_idx,
  input  [5:0]  io_enq_4_dec_uops_3_address_num,
  input  [6:0]  io_enq_4_dec_uops_3_uopc,
  input  [31:0] io_enq_4_dec_uops_3_inst,
  input  [31:0] io_enq_4_dec_uops_3_debug_inst,
  input         io_enq_4_dec_uops_3_is_rvc,
  input  [39:0] io_enq_4_dec_uops_3_debug_pc,
  input  [2:0]  io_enq_4_dec_uops_3_iq_type,
  input  [9:0]  io_enq_4_dec_uops_3_fu_code,
  input  [3:0]  io_enq_4_dec_uops_3_ctrl_br_type,
  input  [1:0]  io_enq_4_dec_uops_3_ctrl_op1_sel,
  input  [2:0]  io_enq_4_dec_uops_3_ctrl_op2_sel,
  input  [2:0]  io_enq_4_dec_uops_3_ctrl_imm_sel,
  input  [3:0]  io_enq_4_dec_uops_3_ctrl_op_fcn,
  input         io_enq_4_dec_uops_3_ctrl_fcn_dw,
  input  [2:0]  io_enq_4_dec_uops_3_ctrl_csr_cmd,
  input         io_enq_4_dec_uops_3_ctrl_is_load,
  input         io_enq_4_dec_uops_3_ctrl_is_sta,
  input         io_enq_4_dec_uops_3_ctrl_is_std,
  input  [1:0]  io_enq_4_dec_uops_3_ctrl_op3_sel,
  input  [1:0]  io_enq_4_dec_uops_3_iw_state,
  input         io_enq_4_dec_uops_3_iw_p1_poisoned,
  input         io_enq_4_dec_uops_3_iw_p2_poisoned,
  input         io_enq_4_dec_uops_3_is_br,
  input         io_enq_4_dec_uops_3_is_jalr,
  input         io_enq_4_dec_uops_3_is_jal,
  input         io_enq_4_dec_uops_3_is_sfb,
  input  [11:0] io_enq_4_dec_uops_3_br_mask,
  input  [3:0]  io_enq_4_dec_uops_3_br_tag,
  input  [4:0]  io_enq_4_dec_uops_3_ftq_idx,
  input         io_enq_4_dec_uops_3_edge_inst,
  input  [5:0]  io_enq_4_dec_uops_3_pc_lob,
  input         io_enq_4_dec_uops_3_taken,
  input  [19:0] io_enq_4_dec_uops_3_imm_packed,
  input  [11:0] io_enq_4_dec_uops_3_csr_addr,
  input  [5:0]  io_enq_4_dec_uops_3_rob_idx,
  input  [4:0]  io_enq_4_dec_uops_3_ldq_idx,
  input  [4:0]  io_enq_4_dec_uops_3_stq_idx,
  input  [1:0]  io_enq_4_dec_uops_3_rxq_idx,
  input  [6:0]  io_enq_4_dec_uops_3_pdst,
  input  [6:0]  io_enq_4_dec_uops_3_prs1,
  input  [6:0]  io_enq_4_dec_uops_3_prs2,
  input  [6:0]  io_enq_4_dec_uops_3_prs3,
  input  [4:0]  io_enq_4_dec_uops_3_ppred,
  input         io_enq_4_dec_uops_3_prs1_busy,
  input         io_enq_4_dec_uops_3_prs2_busy,
  input         io_enq_4_dec_uops_3_prs3_busy,
  input         io_enq_4_dec_uops_3_ppred_busy,
  input  [6:0]  io_enq_4_dec_uops_3_stale_pdst,
  input         io_enq_4_dec_uops_3_exception,
  input  [63:0] io_enq_4_dec_uops_3_exc_cause,
  input         io_enq_4_dec_uops_3_bypassable,
  input  [4:0]  io_enq_4_dec_uops_3_mem_cmd,
  input  [1:0]  io_enq_4_dec_uops_3_mem_size,
  input         io_enq_4_dec_uops_3_mem_signed,
  input         io_enq_4_dec_uops_3_is_fence,
  input         io_enq_4_dec_uops_3_is_fencei,
  input         io_enq_4_dec_uops_3_is_amo,
  input         io_enq_4_dec_uops_3_uses_ldq,
  input         io_enq_4_dec_uops_3_uses_stq,
  input         io_enq_4_dec_uops_3_is_sys_pc2epc,
  input         io_enq_4_dec_uops_3_is_unique,
  input         io_enq_4_dec_uops_3_flush_on_commit,
  input         io_enq_4_dec_uops_3_ldst_is_rs1,
  input  [5:0]  io_enq_4_dec_uops_3_ldst,
  input  [5:0]  io_enq_4_dec_uops_3_lrs1,
  input  [5:0]  io_enq_4_dec_uops_3_lrs2,
  input  [5:0]  io_enq_4_dec_uops_3_lrs3,
  input         io_enq_4_dec_uops_3_ldst_val,
  input  [1:0]  io_enq_4_dec_uops_3_dst_rtype,
  input  [1:0]  io_enq_4_dec_uops_3_lrs1_rtype,
  input  [1:0]  io_enq_4_dec_uops_3_lrs2_rtype,
  input         io_enq_4_dec_uops_3_frs3_en,
  input         io_enq_4_dec_uops_3_fp_val,
  input         io_enq_4_dec_uops_3_fp_single,
  input         io_enq_4_dec_uops_3_xcpt_pf_if,
  input         io_enq_4_dec_uops_3_xcpt_ae_if,
  input         io_enq_4_dec_uops_3_xcpt_ma_if,
  input         io_enq_4_dec_uops_3_bp_debug_if,
  input         io_enq_4_dec_uops_3_bp_xcpt_if,
  input  [1:0]  io_enq_4_dec_uops_3_debug_fsrc,
  input  [1:0]  io_enq_4_dec_uops_3_debug_tsrc,
  input         io_enq_4_val_mask_0,
  input         io_enq_4_val_mask_1,
  input         io_enq_4_val_mask_2,
  input         io_enq_4_val_mask_3,
  input         io_enq_5_dec_uops_0_switch,
  input         io_enq_5_dec_uops_0_switch_off,
  input         io_enq_5_dec_uops_0_is_unicore,
  input  [2:0]  io_enq_5_dec_uops_0_shift,
  input  [1:0]  io_enq_5_dec_uops_0_lrs3_rtype,
  input         io_enq_5_dec_uops_0_rflag,
  input         io_enq_5_dec_uops_0_wflag,
  input  [3:0]  io_enq_5_dec_uops_0_prflag,
  input  [3:0]  io_enq_5_dec_uops_0_pwflag,
  input         io_enq_5_dec_uops_0_pflag_busy,
  input  [3:0]  io_enq_5_dec_uops_0_stale_pflag,
  input  [3:0]  io_enq_5_dec_uops_0_op1_sel,
  input  [3:0]  io_enq_5_dec_uops_0_op2_sel,
  input  [5:0]  io_enq_5_dec_uops_0_split_num,
  input  [5:0]  io_enq_5_dec_uops_0_self_index,
  input  [5:0]  io_enq_5_dec_uops_0_rob_inst_idx,
  input  [5:0]  io_enq_5_dec_uops_0_address_num,
  input  [6:0]  io_enq_5_dec_uops_0_uopc,
  input  [31:0] io_enq_5_dec_uops_0_inst,
  input  [31:0] io_enq_5_dec_uops_0_debug_inst,
  input         io_enq_5_dec_uops_0_is_rvc,
  input  [39:0] io_enq_5_dec_uops_0_debug_pc,
  input  [2:0]  io_enq_5_dec_uops_0_iq_type,
  input  [9:0]  io_enq_5_dec_uops_0_fu_code,
  input  [3:0]  io_enq_5_dec_uops_0_ctrl_br_type,
  input  [1:0]  io_enq_5_dec_uops_0_ctrl_op1_sel,
  input  [2:0]  io_enq_5_dec_uops_0_ctrl_op2_sel,
  input  [2:0]  io_enq_5_dec_uops_0_ctrl_imm_sel,
  input  [3:0]  io_enq_5_dec_uops_0_ctrl_op_fcn,
  input         io_enq_5_dec_uops_0_ctrl_fcn_dw,
  input  [2:0]  io_enq_5_dec_uops_0_ctrl_csr_cmd,
  input         io_enq_5_dec_uops_0_ctrl_is_load,
  input         io_enq_5_dec_uops_0_ctrl_is_sta,
  input         io_enq_5_dec_uops_0_ctrl_is_std,
  input  [1:0]  io_enq_5_dec_uops_0_ctrl_op3_sel,
  input  [1:0]  io_enq_5_dec_uops_0_iw_state,
  input         io_enq_5_dec_uops_0_iw_p1_poisoned,
  input         io_enq_5_dec_uops_0_iw_p2_poisoned,
  input         io_enq_5_dec_uops_0_is_br,
  input         io_enq_5_dec_uops_0_is_jalr,
  input         io_enq_5_dec_uops_0_is_jal,
  input         io_enq_5_dec_uops_0_is_sfb,
  input  [11:0] io_enq_5_dec_uops_0_br_mask,
  input  [3:0]  io_enq_5_dec_uops_0_br_tag,
  input  [4:0]  io_enq_5_dec_uops_0_ftq_idx,
  input         io_enq_5_dec_uops_0_edge_inst,
  input  [5:0]  io_enq_5_dec_uops_0_pc_lob,
  input         io_enq_5_dec_uops_0_taken,
  input  [19:0] io_enq_5_dec_uops_0_imm_packed,
  input  [11:0] io_enq_5_dec_uops_0_csr_addr,
  input  [5:0]  io_enq_5_dec_uops_0_rob_idx,
  input  [4:0]  io_enq_5_dec_uops_0_ldq_idx,
  input  [4:0]  io_enq_5_dec_uops_0_stq_idx,
  input  [1:0]  io_enq_5_dec_uops_0_rxq_idx,
  input  [6:0]  io_enq_5_dec_uops_0_pdst,
  input  [6:0]  io_enq_5_dec_uops_0_prs1,
  input  [6:0]  io_enq_5_dec_uops_0_prs2,
  input  [6:0]  io_enq_5_dec_uops_0_prs3,
  input  [4:0]  io_enq_5_dec_uops_0_ppred,
  input         io_enq_5_dec_uops_0_prs1_busy,
  input         io_enq_5_dec_uops_0_prs2_busy,
  input         io_enq_5_dec_uops_0_prs3_busy,
  input         io_enq_5_dec_uops_0_ppred_busy,
  input  [6:0]  io_enq_5_dec_uops_0_stale_pdst,
  input         io_enq_5_dec_uops_0_exception,
  input  [63:0] io_enq_5_dec_uops_0_exc_cause,
  input         io_enq_5_dec_uops_0_bypassable,
  input  [4:0]  io_enq_5_dec_uops_0_mem_cmd,
  input  [1:0]  io_enq_5_dec_uops_0_mem_size,
  input         io_enq_5_dec_uops_0_mem_signed,
  input         io_enq_5_dec_uops_0_is_fence,
  input         io_enq_5_dec_uops_0_is_fencei,
  input         io_enq_5_dec_uops_0_is_amo,
  input         io_enq_5_dec_uops_0_uses_ldq,
  input         io_enq_5_dec_uops_0_uses_stq,
  input         io_enq_5_dec_uops_0_is_sys_pc2epc,
  input         io_enq_5_dec_uops_0_is_unique,
  input         io_enq_5_dec_uops_0_flush_on_commit,
  input         io_enq_5_dec_uops_0_ldst_is_rs1,
  input  [5:0]  io_enq_5_dec_uops_0_ldst,
  input  [5:0]  io_enq_5_dec_uops_0_lrs1,
  input  [5:0]  io_enq_5_dec_uops_0_lrs2,
  input  [5:0]  io_enq_5_dec_uops_0_lrs3,
  input         io_enq_5_dec_uops_0_ldst_val,
  input  [1:0]  io_enq_5_dec_uops_0_dst_rtype,
  input  [1:0]  io_enq_5_dec_uops_0_lrs1_rtype,
  input  [1:0]  io_enq_5_dec_uops_0_lrs2_rtype,
  input         io_enq_5_dec_uops_0_frs3_en,
  input         io_enq_5_dec_uops_0_fp_val,
  input         io_enq_5_dec_uops_0_fp_single,
  input         io_enq_5_dec_uops_0_xcpt_pf_if,
  input         io_enq_5_dec_uops_0_xcpt_ae_if,
  input         io_enq_5_dec_uops_0_xcpt_ma_if,
  input         io_enq_5_dec_uops_0_bp_debug_if,
  input         io_enq_5_dec_uops_0_bp_xcpt_if,
  input  [1:0]  io_enq_5_dec_uops_0_debug_fsrc,
  input  [1:0]  io_enq_5_dec_uops_0_debug_tsrc,
  input         io_enq_5_dec_uops_1_switch,
  input         io_enq_5_dec_uops_1_switch_off,
  input         io_enq_5_dec_uops_1_is_unicore,
  input  [2:0]  io_enq_5_dec_uops_1_shift,
  input  [1:0]  io_enq_5_dec_uops_1_lrs3_rtype,
  input         io_enq_5_dec_uops_1_rflag,
  input         io_enq_5_dec_uops_1_wflag,
  input  [3:0]  io_enq_5_dec_uops_1_prflag,
  input  [3:0]  io_enq_5_dec_uops_1_pwflag,
  input         io_enq_5_dec_uops_1_pflag_busy,
  input  [3:0]  io_enq_5_dec_uops_1_stale_pflag,
  input  [3:0]  io_enq_5_dec_uops_1_op1_sel,
  input  [3:0]  io_enq_5_dec_uops_1_op2_sel,
  input  [5:0]  io_enq_5_dec_uops_1_split_num,
  input  [5:0]  io_enq_5_dec_uops_1_self_index,
  input  [5:0]  io_enq_5_dec_uops_1_rob_inst_idx,
  input  [5:0]  io_enq_5_dec_uops_1_address_num,
  input  [6:0]  io_enq_5_dec_uops_1_uopc,
  input  [31:0] io_enq_5_dec_uops_1_inst,
  input  [31:0] io_enq_5_dec_uops_1_debug_inst,
  input         io_enq_5_dec_uops_1_is_rvc,
  input  [39:0] io_enq_5_dec_uops_1_debug_pc,
  input  [2:0]  io_enq_5_dec_uops_1_iq_type,
  input  [9:0]  io_enq_5_dec_uops_1_fu_code,
  input  [3:0]  io_enq_5_dec_uops_1_ctrl_br_type,
  input  [1:0]  io_enq_5_dec_uops_1_ctrl_op1_sel,
  input  [2:0]  io_enq_5_dec_uops_1_ctrl_op2_sel,
  input  [2:0]  io_enq_5_dec_uops_1_ctrl_imm_sel,
  input  [3:0]  io_enq_5_dec_uops_1_ctrl_op_fcn,
  input         io_enq_5_dec_uops_1_ctrl_fcn_dw,
  input  [2:0]  io_enq_5_dec_uops_1_ctrl_csr_cmd,
  input         io_enq_5_dec_uops_1_ctrl_is_load,
  input         io_enq_5_dec_uops_1_ctrl_is_sta,
  input         io_enq_5_dec_uops_1_ctrl_is_std,
  input  [1:0]  io_enq_5_dec_uops_1_ctrl_op3_sel,
  input  [1:0]  io_enq_5_dec_uops_1_iw_state,
  input         io_enq_5_dec_uops_1_iw_p1_poisoned,
  input         io_enq_5_dec_uops_1_iw_p2_poisoned,
  input         io_enq_5_dec_uops_1_is_br,
  input         io_enq_5_dec_uops_1_is_jalr,
  input         io_enq_5_dec_uops_1_is_jal,
  input         io_enq_5_dec_uops_1_is_sfb,
  input  [11:0] io_enq_5_dec_uops_1_br_mask,
  input  [3:0]  io_enq_5_dec_uops_1_br_tag,
  input  [4:0]  io_enq_5_dec_uops_1_ftq_idx,
  input         io_enq_5_dec_uops_1_edge_inst,
  input  [5:0]  io_enq_5_dec_uops_1_pc_lob,
  input         io_enq_5_dec_uops_1_taken,
  input  [19:0] io_enq_5_dec_uops_1_imm_packed,
  input  [11:0] io_enq_5_dec_uops_1_csr_addr,
  input  [5:0]  io_enq_5_dec_uops_1_rob_idx,
  input  [4:0]  io_enq_5_dec_uops_1_ldq_idx,
  input  [4:0]  io_enq_5_dec_uops_1_stq_idx,
  input  [1:0]  io_enq_5_dec_uops_1_rxq_idx,
  input  [6:0]  io_enq_5_dec_uops_1_pdst,
  input  [6:0]  io_enq_5_dec_uops_1_prs1,
  input  [6:0]  io_enq_5_dec_uops_1_prs2,
  input  [6:0]  io_enq_5_dec_uops_1_prs3,
  input  [4:0]  io_enq_5_dec_uops_1_ppred,
  input         io_enq_5_dec_uops_1_prs1_busy,
  input         io_enq_5_dec_uops_1_prs2_busy,
  input         io_enq_5_dec_uops_1_prs3_busy,
  input         io_enq_5_dec_uops_1_ppred_busy,
  input  [6:0]  io_enq_5_dec_uops_1_stale_pdst,
  input         io_enq_5_dec_uops_1_exception,
  input  [63:0] io_enq_5_dec_uops_1_exc_cause,
  input         io_enq_5_dec_uops_1_bypassable,
  input  [4:0]  io_enq_5_dec_uops_1_mem_cmd,
  input  [1:0]  io_enq_5_dec_uops_1_mem_size,
  input         io_enq_5_dec_uops_1_mem_signed,
  input         io_enq_5_dec_uops_1_is_fence,
  input         io_enq_5_dec_uops_1_is_fencei,
  input         io_enq_5_dec_uops_1_is_amo,
  input         io_enq_5_dec_uops_1_uses_ldq,
  input         io_enq_5_dec_uops_1_uses_stq,
  input         io_enq_5_dec_uops_1_is_sys_pc2epc,
  input         io_enq_5_dec_uops_1_is_unique,
  input         io_enq_5_dec_uops_1_flush_on_commit,
  input         io_enq_5_dec_uops_1_ldst_is_rs1,
  input  [5:0]  io_enq_5_dec_uops_1_ldst,
  input  [5:0]  io_enq_5_dec_uops_1_lrs1,
  input  [5:0]  io_enq_5_dec_uops_1_lrs2,
  input  [5:0]  io_enq_5_dec_uops_1_lrs3,
  input         io_enq_5_dec_uops_1_ldst_val,
  input  [1:0]  io_enq_5_dec_uops_1_dst_rtype,
  input  [1:0]  io_enq_5_dec_uops_1_lrs1_rtype,
  input  [1:0]  io_enq_5_dec_uops_1_lrs2_rtype,
  input         io_enq_5_dec_uops_1_frs3_en,
  input         io_enq_5_dec_uops_1_fp_val,
  input         io_enq_5_dec_uops_1_fp_single,
  input         io_enq_5_dec_uops_1_xcpt_pf_if,
  input         io_enq_5_dec_uops_1_xcpt_ae_if,
  input         io_enq_5_dec_uops_1_xcpt_ma_if,
  input         io_enq_5_dec_uops_1_bp_debug_if,
  input         io_enq_5_dec_uops_1_bp_xcpt_if,
  input  [1:0]  io_enq_5_dec_uops_1_debug_fsrc,
  input  [1:0]  io_enq_5_dec_uops_1_debug_tsrc,
  input         io_enq_5_dec_uops_2_switch,
  input         io_enq_5_dec_uops_2_switch_off,
  input         io_enq_5_dec_uops_2_is_unicore,
  input  [2:0]  io_enq_5_dec_uops_2_shift,
  input  [1:0]  io_enq_5_dec_uops_2_lrs3_rtype,
  input         io_enq_5_dec_uops_2_rflag,
  input         io_enq_5_dec_uops_2_wflag,
  input  [3:0]  io_enq_5_dec_uops_2_prflag,
  input  [3:0]  io_enq_5_dec_uops_2_pwflag,
  input         io_enq_5_dec_uops_2_pflag_busy,
  input  [3:0]  io_enq_5_dec_uops_2_stale_pflag,
  input  [3:0]  io_enq_5_dec_uops_2_op1_sel,
  input  [3:0]  io_enq_5_dec_uops_2_op2_sel,
  input  [5:0]  io_enq_5_dec_uops_2_split_num,
  input  [5:0]  io_enq_5_dec_uops_2_self_index,
  input  [5:0]  io_enq_5_dec_uops_2_rob_inst_idx,
  input  [5:0]  io_enq_5_dec_uops_2_address_num,
  input  [6:0]  io_enq_5_dec_uops_2_uopc,
  input  [31:0] io_enq_5_dec_uops_2_inst,
  input  [31:0] io_enq_5_dec_uops_2_debug_inst,
  input         io_enq_5_dec_uops_2_is_rvc,
  input  [39:0] io_enq_5_dec_uops_2_debug_pc,
  input  [2:0]  io_enq_5_dec_uops_2_iq_type,
  input  [9:0]  io_enq_5_dec_uops_2_fu_code,
  input  [3:0]  io_enq_5_dec_uops_2_ctrl_br_type,
  input  [1:0]  io_enq_5_dec_uops_2_ctrl_op1_sel,
  input  [2:0]  io_enq_5_dec_uops_2_ctrl_op2_sel,
  input  [2:0]  io_enq_5_dec_uops_2_ctrl_imm_sel,
  input  [3:0]  io_enq_5_dec_uops_2_ctrl_op_fcn,
  input         io_enq_5_dec_uops_2_ctrl_fcn_dw,
  input  [2:0]  io_enq_5_dec_uops_2_ctrl_csr_cmd,
  input         io_enq_5_dec_uops_2_ctrl_is_load,
  input         io_enq_5_dec_uops_2_ctrl_is_sta,
  input         io_enq_5_dec_uops_2_ctrl_is_std,
  input  [1:0]  io_enq_5_dec_uops_2_ctrl_op3_sel,
  input  [1:0]  io_enq_5_dec_uops_2_iw_state,
  input         io_enq_5_dec_uops_2_iw_p1_poisoned,
  input         io_enq_5_dec_uops_2_iw_p2_poisoned,
  input         io_enq_5_dec_uops_2_is_br,
  input         io_enq_5_dec_uops_2_is_jalr,
  input         io_enq_5_dec_uops_2_is_jal,
  input         io_enq_5_dec_uops_2_is_sfb,
  input  [11:0] io_enq_5_dec_uops_2_br_mask,
  input  [3:0]  io_enq_5_dec_uops_2_br_tag,
  input  [4:0]  io_enq_5_dec_uops_2_ftq_idx,
  input         io_enq_5_dec_uops_2_edge_inst,
  input  [5:0]  io_enq_5_dec_uops_2_pc_lob,
  input         io_enq_5_dec_uops_2_taken,
  input  [19:0] io_enq_5_dec_uops_2_imm_packed,
  input  [11:0] io_enq_5_dec_uops_2_csr_addr,
  input  [5:0]  io_enq_5_dec_uops_2_rob_idx,
  input  [4:0]  io_enq_5_dec_uops_2_ldq_idx,
  input  [4:0]  io_enq_5_dec_uops_2_stq_idx,
  input  [1:0]  io_enq_5_dec_uops_2_rxq_idx,
  input  [6:0]  io_enq_5_dec_uops_2_pdst,
  input  [6:0]  io_enq_5_dec_uops_2_prs1,
  input  [6:0]  io_enq_5_dec_uops_2_prs2,
  input  [6:0]  io_enq_5_dec_uops_2_prs3,
  input  [4:0]  io_enq_5_dec_uops_2_ppred,
  input         io_enq_5_dec_uops_2_prs1_busy,
  input         io_enq_5_dec_uops_2_prs2_busy,
  input         io_enq_5_dec_uops_2_prs3_busy,
  input         io_enq_5_dec_uops_2_ppred_busy,
  input  [6:0]  io_enq_5_dec_uops_2_stale_pdst,
  input         io_enq_5_dec_uops_2_exception,
  input  [63:0] io_enq_5_dec_uops_2_exc_cause,
  input         io_enq_5_dec_uops_2_bypassable,
  input  [4:0]  io_enq_5_dec_uops_2_mem_cmd,
  input  [1:0]  io_enq_5_dec_uops_2_mem_size,
  input         io_enq_5_dec_uops_2_mem_signed,
  input         io_enq_5_dec_uops_2_is_fence,
  input         io_enq_5_dec_uops_2_is_fencei,
  input         io_enq_5_dec_uops_2_is_amo,
  input         io_enq_5_dec_uops_2_uses_ldq,
  input         io_enq_5_dec_uops_2_uses_stq,
  input         io_enq_5_dec_uops_2_is_sys_pc2epc,
  input         io_enq_5_dec_uops_2_is_unique,
  input         io_enq_5_dec_uops_2_flush_on_commit,
  input         io_enq_5_dec_uops_2_ldst_is_rs1,
  input  [5:0]  io_enq_5_dec_uops_2_ldst,
  input  [5:0]  io_enq_5_dec_uops_2_lrs1,
  input  [5:0]  io_enq_5_dec_uops_2_lrs2,
  input  [5:0]  io_enq_5_dec_uops_2_lrs3,
  input         io_enq_5_dec_uops_2_ldst_val,
  input  [1:0]  io_enq_5_dec_uops_2_dst_rtype,
  input  [1:0]  io_enq_5_dec_uops_2_lrs1_rtype,
  input  [1:0]  io_enq_5_dec_uops_2_lrs2_rtype,
  input         io_enq_5_dec_uops_2_frs3_en,
  input         io_enq_5_dec_uops_2_fp_val,
  input         io_enq_5_dec_uops_2_fp_single,
  input         io_enq_5_dec_uops_2_xcpt_pf_if,
  input         io_enq_5_dec_uops_2_xcpt_ae_if,
  input         io_enq_5_dec_uops_2_xcpt_ma_if,
  input         io_enq_5_dec_uops_2_bp_debug_if,
  input         io_enq_5_dec_uops_2_bp_xcpt_if,
  input  [1:0]  io_enq_5_dec_uops_2_debug_fsrc,
  input  [1:0]  io_enq_5_dec_uops_2_debug_tsrc,
  input         io_enq_5_dec_uops_3_switch,
  input         io_enq_5_dec_uops_3_switch_off,
  input         io_enq_5_dec_uops_3_is_unicore,
  input  [2:0]  io_enq_5_dec_uops_3_shift,
  input  [1:0]  io_enq_5_dec_uops_3_lrs3_rtype,
  input         io_enq_5_dec_uops_3_rflag,
  input         io_enq_5_dec_uops_3_wflag,
  input  [3:0]  io_enq_5_dec_uops_3_prflag,
  input  [3:0]  io_enq_5_dec_uops_3_pwflag,
  input         io_enq_5_dec_uops_3_pflag_busy,
  input  [3:0]  io_enq_5_dec_uops_3_stale_pflag,
  input  [3:0]  io_enq_5_dec_uops_3_op1_sel,
  input  [3:0]  io_enq_5_dec_uops_3_op2_sel,
  input  [5:0]  io_enq_5_dec_uops_3_split_num,
  input  [5:0]  io_enq_5_dec_uops_3_self_index,
  input  [5:0]  io_enq_5_dec_uops_3_rob_inst_idx,
  input  [5:0]  io_enq_5_dec_uops_3_address_num,
  input  [6:0]  io_enq_5_dec_uops_3_uopc,
  input  [31:0] io_enq_5_dec_uops_3_inst,
  input  [31:0] io_enq_5_dec_uops_3_debug_inst,
  input         io_enq_5_dec_uops_3_is_rvc,
  input  [39:0] io_enq_5_dec_uops_3_debug_pc,
  input  [2:0]  io_enq_5_dec_uops_3_iq_type,
  input  [9:0]  io_enq_5_dec_uops_3_fu_code,
  input  [3:0]  io_enq_5_dec_uops_3_ctrl_br_type,
  input  [1:0]  io_enq_5_dec_uops_3_ctrl_op1_sel,
  input  [2:0]  io_enq_5_dec_uops_3_ctrl_op2_sel,
  input  [2:0]  io_enq_5_dec_uops_3_ctrl_imm_sel,
  input  [3:0]  io_enq_5_dec_uops_3_ctrl_op_fcn,
  input         io_enq_5_dec_uops_3_ctrl_fcn_dw,
  input  [2:0]  io_enq_5_dec_uops_3_ctrl_csr_cmd,
  input         io_enq_5_dec_uops_3_ctrl_is_load,
  input         io_enq_5_dec_uops_3_ctrl_is_sta,
  input         io_enq_5_dec_uops_3_ctrl_is_std,
  input  [1:0]  io_enq_5_dec_uops_3_ctrl_op3_sel,
  input  [1:0]  io_enq_5_dec_uops_3_iw_state,
  input         io_enq_5_dec_uops_3_iw_p1_poisoned,
  input         io_enq_5_dec_uops_3_iw_p2_poisoned,
  input         io_enq_5_dec_uops_3_is_br,
  input         io_enq_5_dec_uops_3_is_jalr,
  input         io_enq_5_dec_uops_3_is_jal,
  input         io_enq_5_dec_uops_3_is_sfb,
  input  [11:0] io_enq_5_dec_uops_3_br_mask,
  input  [3:0]  io_enq_5_dec_uops_3_br_tag,
  input  [4:0]  io_enq_5_dec_uops_3_ftq_idx,
  input         io_enq_5_dec_uops_3_edge_inst,
  input  [5:0]  io_enq_5_dec_uops_3_pc_lob,
  input         io_enq_5_dec_uops_3_taken,
  input  [19:0] io_enq_5_dec_uops_3_imm_packed,
  input  [11:0] io_enq_5_dec_uops_3_csr_addr,
  input  [5:0]  io_enq_5_dec_uops_3_rob_idx,
  input  [4:0]  io_enq_5_dec_uops_3_ldq_idx,
  input  [4:0]  io_enq_5_dec_uops_3_stq_idx,
  input  [1:0]  io_enq_5_dec_uops_3_rxq_idx,
  input  [6:0]  io_enq_5_dec_uops_3_pdst,
  input  [6:0]  io_enq_5_dec_uops_3_prs1,
  input  [6:0]  io_enq_5_dec_uops_3_prs2,
  input  [6:0]  io_enq_5_dec_uops_3_prs3,
  input  [4:0]  io_enq_5_dec_uops_3_ppred,
  input         io_enq_5_dec_uops_3_prs1_busy,
  input         io_enq_5_dec_uops_3_prs2_busy,
  input         io_enq_5_dec_uops_3_prs3_busy,
  input         io_enq_5_dec_uops_3_ppred_busy,
  input  [6:0]  io_enq_5_dec_uops_3_stale_pdst,
  input         io_enq_5_dec_uops_3_exception,
  input  [63:0] io_enq_5_dec_uops_3_exc_cause,
  input         io_enq_5_dec_uops_3_bypassable,
  input  [4:0]  io_enq_5_dec_uops_3_mem_cmd,
  input  [1:0]  io_enq_5_dec_uops_3_mem_size,
  input         io_enq_5_dec_uops_3_mem_signed,
  input         io_enq_5_dec_uops_3_is_fence,
  input         io_enq_5_dec_uops_3_is_fencei,
  input         io_enq_5_dec_uops_3_is_amo,
  input         io_enq_5_dec_uops_3_uses_ldq,
  input         io_enq_5_dec_uops_3_uses_stq,
  input         io_enq_5_dec_uops_3_is_sys_pc2epc,
  input         io_enq_5_dec_uops_3_is_unique,
  input         io_enq_5_dec_uops_3_flush_on_commit,
  input         io_enq_5_dec_uops_3_ldst_is_rs1,
  input  [5:0]  io_enq_5_dec_uops_3_ldst,
  input  [5:0]  io_enq_5_dec_uops_3_lrs1,
  input  [5:0]  io_enq_5_dec_uops_3_lrs2,
  input  [5:0]  io_enq_5_dec_uops_3_lrs3,
  input         io_enq_5_dec_uops_3_ldst_val,
  input  [1:0]  io_enq_5_dec_uops_3_dst_rtype,
  input  [1:0]  io_enq_5_dec_uops_3_lrs1_rtype,
  input  [1:0]  io_enq_5_dec_uops_3_lrs2_rtype,
  input         io_enq_5_dec_uops_3_frs3_en,
  input         io_enq_5_dec_uops_3_fp_val,
  input         io_enq_5_dec_uops_3_fp_single,
  input         io_enq_5_dec_uops_3_xcpt_pf_if,
  input         io_enq_5_dec_uops_3_xcpt_ae_if,
  input         io_enq_5_dec_uops_3_xcpt_ma_if,
  input         io_enq_5_dec_uops_3_bp_debug_if,
  input         io_enq_5_dec_uops_3_bp_xcpt_if,
  input  [1:0]  io_enq_5_dec_uops_3_debug_fsrc,
  input  [1:0]  io_enq_5_dec_uops_3_debug_tsrc,
  input         io_enq_5_val_mask_0,
  input         io_enq_5_val_mask_1,
  input         io_enq_5_val_mask_2,
  input         io_enq_5_val_mask_3,
  input         io_enq_6_dec_uops_0_switch,
  input         io_enq_6_dec_uops_0_switch_off,
  input         io_enq_6_dec_uops_0_is_unicore,
  input  [2:0]  io_enq_6_dec_uops_0_shift,
  input  [1:0]  io_enq_6_dec_uops_0_lrs3_rtype,
  input         io_enq_6_dec_uops_0_rflag,
  input         io_enq_6_dec_uops_0_wflag,
  input  [3:0]  io_enq_6_dec_uops_0_prflag,
  input  [3:0]  io_enq_6_dec_uops_0_pwflag,
  input         io_enq_6_dec_uops_0_pflag_busy,
  input  [3:0]  io_enq_6_dec_uops_0_stale_pflag,
  input  [3:0]  io_enq_6_dec_uops_0_op1_sel,
  input  [3:0]  io_enq_6_dec_uops_0_op2_sel,
  input  [5:0]  io_enq_6_dec_uops_0_split_num,
  input  [5:0]  io_enq_6_dec_uops_0_self_index,
  input  [5:0]  io_enq_6_dec_uops_0_rob_inst_idx,
  input  [5:0]  io_enq_6_dec_uops_0_address_num,
  input  [6:0]  io_enq_6_dec_uops_0_uopc,
  input  [31:0] io_enq_6_dec_uops_0_inst,
  input  [31:0] io_enq_6_dec_uops_0_debug_inst,
  input         io_enq_6_dec_uops_0_is_rvc,
  input  [39:0] io_enq_6_dec_uops_0_debug_pc,
  input  [2:0]  io_enq_6_dec_uops_0_iq_type,
  input  [9:0]  io_enq_6_dec_uops_0_fu_code,
  input  [3:0]  io_enq_6_dec_uops_0_ctrl_br_type,
  input  [1:0]  io_enq_6_dec_uops_0_ctrl_op1_sel,
  input  [2:0]  io_enq_6_dec_uops_0_ctrl_op2_sel,
  input  [2:0]  io_enq_6_dec_uops_0_ctrl_imm_sel,
  input  [3:0]  io_enq_6_dec_uops_0_ctrl_op_fcn,
  input         io_enq_6_dec_uops_0_ctrl_fcn_dw,
  input  [2:0]  io_enq_6_dec_uops_0_ctrl_csr_cmd,
  input         io_enq_6_dec_uops_0_ctrl_is_load,
  input         io_enq_6_dec_uops_0_ctrl_is_sta,
  input         io_enq_6_dec_uops_0_ctrl_is_std,
  input  [1:0]  io_enq_6_dec_uops_0_ctrl_op3_sel,
  input  [1:0]  io_enq_6_dec_uops_0_iw_state,
  input         io_enq_6_dec_uops_0_iw_p1_poisoned,
  input         io_enq_6_dec_uops_0_iw_p2_poisoned,
  input         io_enq_6_dec_uops_0_is_br,
  input         io_enq_6_dec_uops_0_is_jalr,
  input         io_enq_6_dec_uops_0_is_jal,
  input         io_enq_6_dec_uops_0_is_sfb,
  input  [11:0] io_enq_6_dec_uops_0_br_mask,
  input  [3:0]  io_enq_6_dec_uops_0_br_tag,
  input  [4:0]  io_enq_6_dec_uops_0_ftq_idx,
  input         io_enq_6_dec_uops_0_edge_inst,
  input  [5:0]  io_enq_6_dec_uops_0_pc_lob,
  input         io_enq_6_dec_uops_0_taken,
  input  [19:0] io_enq_6_dec_uops_0_imm_packed,
  input  [11:0] io_enq_6_dec_uops_0_csr_addr,
  input  [5:0]  io_enq_6_dec_uops_0_rob_idx,
  input  [4:0]  io_enq_6_dec_uops_0_ldq_idx,
  input  [4:0]  io_enq_6_dec_uops_0_stq_idx,
  input  [1:0]  io_enq_6_dec_uops_0_rxq_idx,
  input  [6:0]  io_enq_6_dec_uops_0_pdst,
  input  [6:0]  io_enq_6_dec_uops_0_prs1,
  input  [6:0]  io_enq_6_dec_uops_0_prs2,
  input  [6:0]  io_enq_6_dec_uops_0_prs3,
  input  [4:0]  io_enq_6_dec_uops_0_ppred,
  input         io_enq_6_dec_uops_0_prs1_busy,
  input         io_enq_6_dec_uops_0_prs2_busy,
  input         io_enq_6_dec_uops_0_prs3_busy,
  input         io_enq_6_dec_uops_0_ppred_busy,
  input  [6:0]  io_enq_6_dec_uops_0_stale_pdst,
  input         io_enq_6_dec_uops_0_exception,
  input  [63:0] io_enq_6_dec_uops_0_exc_cause,
  input         io_enq_6_dec_uops_0_bypassable,
  input  [4:0]  io_enq_6_dec_uops_0_mem_cmd,
  input  [1:0]  io_enq_6_dec_uops_0_mem_size,
  input         io_enq_6_dec_uops_0_mem_signed,
  input         io_enq_6_dec_uops_0_is_fence,
  input         io_enq_6_dec_uops_0_is_fencei,
  input         io_enq_6_dec_uops_0_is_amo,
  input         io_enq_6_dec_uops_0_uses_ldq,
  input         io_enq_6_dec_uops_0_uses_stq,
  input         io_enq_6_dec_uops_0_is_sys_pc2epc,
  input         io_enq_6_dec_uops_0_is_unique,
  input         io_enq_6_dec_uops_0_flush_on_commit,
  input         io_enq_6_dec_uops_0_ldst_is_rs1,
  input  [5:0]  io_enq_6_dec_uops_0_ldst,
  input  [5:0]  io_enq_6_dec_uops_0_lrs1,
  input  [5:0]  io_enq_6_dec_uops_0_lrs2,
  input  [5:0]  io_enq_6_dec_uops_0_lrs3,
  input         io_enq_6_dec_uops_0_ldst_val,
  input  [1:0]  io_enq_6_dec_uops_0_dst_rtype,
  input  [1:0]  io_enq_6_dec_uops_0_lrs1_rtype,
  input  [1:0]  io_enq_6_dec_uops_0_lrs2_rtype,
  input         io_enq_6_dec_uops_0_frs3_en,
  input         io_enq_6_dec_uops_0_fp_val,
  input         io_enq_6_dec_uops_0_fp_single,
  input         io_enq_6_dec_uops_0_xcpt_pf_if,
  input         io_enq_6_dec_uops_0_xcpt_ae_if,
  input         io_enq_6_dec_uops_0_xcpt_ma_if,
  input         io_enq_6_dec_uops_0_bp_debug_if,
  input         io_enq_6_dec_uops_0_bp_xcpt_if,
  input  [1:0]  io_enq_6_dec_uops_0_debug_fsrc,
  input  [1:0]  io_enq_6_dec_uops_0_debug_tsrc,
  input         io_enq_6_dec_uops_1_switch,
  input         io_enq_6_dec_uops_1_switch_off,
  input         io_enq_6_dec_uops_1_is_unicore,
  input  [2:0]  io_enq_6_dec_uops_1_shift,
  input  [1:0]  io_enq_6_dec_uops_1_lrs3_rtype,
  input         io_enq_6_dec_uops_1_rflag,
  input         io_enq_6_dec_uops_1_wflag,
  input  [3:0]  io_enq_6_dec_uops_1_prflag,
  input  [3:0]  io_enq_6_dec_uops_1_pwflag,
  input         io_enq_6_dec_uops_1_pflag_busy,
  input  [3:0]  io_enq_6_dec_uops_1_stale_pflag,
  input  [3:0]  io_enq_6_dec_uops_1_op1_sel,
  input  [3:0]  io_enq_6_dec_uops_1_op2_sel,
  input  [5:0]  io_enq_6_dec_uops_1_split_num,
  input  [5:0]  io_enq_6_dec_uops_1_self_index,
  input  [5:0]  io_enq_6_dec_uops_1_rob_inst_idx,
  input  [5:0]  io_enq_6_dec_uops_1_address_num,
  input  [6:0]  io_enq_6_dec_uops_1_uopc,
  input  [31:0] io_enq_6_dec_uops_1_inst,
  input  [31:0] io_enq_6_dec_uops_1_debug_inst,
  input         io_enq_6_dec_uops_1_is_rvc,
  input  [39:0] io_enq_6_dec_uops_1_debug_pc,
  input  [2:0]  io_enq_6_dec_uops_1_iq_type,
  input  [9:0]  io_enq_6_dec_uops_1_fu_code,
  input  [3:0]  io_enq_6_dec_uops_1_ctrl_br_type,
  input  [1:0]  io_enq_6_dec_uops_1_ctrl_op1_sel,
  input  [2:0]  io_enq_6_dec_uops_1_ctrl_op2_sel,
  input  [2:0]  io_enq_6_dec_uops_1_ctrl_imm_sel,
  input  [3:0]  io_enq_6_dec_uops_1_ctrl_op_fcn,
  input         io_enq_6_dec_uops_1_ctrl_fcn_dw,
  input  [2:0]  io_enq_6_dec_uops_1_ctrl_csr_cmd,
  input         io_enq_6_dec_uops_1_ctrl_is_load,
  input         io_enq_6_dec_uops_1_ctrl_is_sta,
  input         io_enq_6_dec_uops_1_ctrl_is_std,
  input  [1:0]  io_enq_6_dec_uops_1_ctrl_op3_sel,
  input  [1:0]  io_enq_6_dec_uops_1_iw_state,
  input         io_enq_6_dec_uops_1_iw_p1_poisoned,
  input         io_enq_6_dec_uops_1_iw_p2_poisoned,
  input         io_enq_6_dec_uops_1_is_br,
  input         io_enq_6_dec_uops_1_is_jalr,
  input         io_enq_6_dec_uops_1_is_jal,
  input         io_enq_6_dec_uops_1_is_sfb,
  input  [11:0] io_enq_6_dec_uops_1_br_mask,
  input  [3:0]  io_enq_6_dec_uops_1_br_tag,
  input  [4:0]  io_enq_6_dec_uops_1_ftq_idx,
  input         io_enq_6_dec_uops_1_edge_inst,
  input  [5:0]  io_enq_6_dec_uops_1_pc_lob,
  input         io_enq_6_dec_uops_1_taken,
  input  [19:0] io_enq_6_dec_uops_1_imm_packed,
  input  [11:0] io_enq_6_dec_uops_1_csr_addr,
  input  [5:0]  io_enq_6_dec_uops_1_rob_idx,
  input  [4:0]  io_enq_6_dec_uops_1_ldq_idx,
  input  [4:0]  io_enq_6_dec_uops_1_stq_idx,
  input  [1:0]  io_enq_6_dec_uops_1_rxq_idx,
  input  [6:0]  io_enq_6_dec_uops_1_pdst,
  input  [6:0]  io_enq_6_dec_uops_1_prs1,
  input  [6:0]  io_enq_6_dec_uops_1_prs2,
  input  [6:0]  io_enq_6_dec_uops_1_prs3,
  input  [4:0]  io_enq_6_dec_uops_1_ppred,
  input         io_enq_6_dec_uops_1_prs1_busy,
  input         io_enq_6_dec_uops_1_prs2_busy,
  input         io_enq_6_dec_uops_1_prs3_busy,
  input         io_enq_6_dec_uops_1_ppred_busy,
  input  [6:0]  io_enq_6_dec_uops_1_stale_pdst,
  input         io_enq_6_dec_uops_1_exception,
  input  [63:0] io_enq_6_dec_uops_1_exc_cause,
  input         io_enq_6_dec_uops_1_bypassable,
  input  [4:0]  io_enq_6_dec_uops_1_mem_cmd,
  input  [1:0]  io_enq_6_dec_uops_1_mem_size,
  input         io_enq_6_dec_uops_1_mem_signed,
  input         io_enq_6_dec_uops_1_is_fence,
  input         io_enq_6_dec_uops_1_is_fencei,
  input         io_enq_6_dec_uops_1_is_amo,
  input         io_enq_6_dec_uops_1_uses_ldq,
  input         io_enq_6_dec_uops_1_uses_stq,
  input         io_enq_6_dec_uops_1_is_sys_pc2epc,
  input         io_enq_6_dec_uops_1_is_unique,
  input         io_enq_6_dec_uops_1_flush_on_commit,
  input         io_enq_6_dec_uops_1_ldst_is_rs1,
  input  [5:0]  io_enq_6_dec_uops_1_ldst,
  input  [5:0]  io_enq_6_dec_uops_1_lrs1,
  input  [5:0]  io_enq_6_dec_uops_1_lrs2,
  input  [5:0]  io_enq_6_dec_uops_1_lrs3,
  input         io_enq_6_dec_uops_1_ldst_val,
  input  [1:0]  io_enq_6_dec_uops_1_dst_rtype,
  input  [1:0]  io_enq_6_dec_uops_1_lrs1_rtype,
  input  [1:0]  io_enq_6_dec_uops_1_lrs2_rtype,
  input         io_enq_6_dec_uops_1_frs3_en,
  input         io_enq_6_dec_uops_1_fp_val,
  input         io_enq_6_dec_uops_1_fp_single,
  input         io_enq_6_dec_uops_1_xcpt_pf_if,
  input         io_enq_6_dec_uops_1_xcpt_ae_if,
  input         io_enq_6_dec_uops_1_xcpt_ma_if,
  input         io_enq_6_dec_uops_1_bp_debug_if,
  input         io_enq_6_dec_uops_1_bp_xcpt_if,
  input  [1:0]  io_enq_6_dec_uops_1_debug_fsrc,
  input  [1:0]  io_enq_6_dec_uops_1_debug_tsrc,
  input         io_enq_6_dec_uops_2_switch,
  input         io_enq_6_dec_uops_2_switch_off,
  input         io_enq_6_dec_uops_2_is_unicore,
  input  [2:0]  io_enq_6_dec_uops_2_shift,
  input  [1:0]  io_enq_6_dec_uops_2_lrs3_rtype,
  input         io_enq_6_dec_uops_2_rflag,
  input         io_enq_6_dec_uops_2_wflag,
  input  [3:0]  io_enq_6_dec_uops_2_prflag,
  input  [3:0]  io_enq_6_dec_uops_2_pwflag,
  input         io_enq_6_dec_uops_2_pflag_busy,
  input  [3:0]  io_enq_6_dec_uops_2_stale_pflag,
  input  [3:0]  io_enq_6_dec_uops_2_op1_sel,
  input  [3:0]  io_enq_6_dec_uops_2_op2_sel,
  input  [5:0]  io_enq_6_dec_uops_2_split_num,
  input  [5:0]  io_enq_6_dec_uops_2_self_index,
  input  [5:0]  io_enq_6_dec_uops_2_rob_inst_idx,
  input  [5:0]  io_enq_6_dec_uops_2_address_num,
  input  [6:0]  io_enq_6_dec_uops_2_uopc,
  input  [31:0] io_enq_6_dec_uops_2_inst,
  input  [31:0] io_enq_6_dec_uops_2_debug_inst,
  input         io_enq_6_dec_uops_2_is_rvc,
  input  [39:0] io_enq_6_dec_uops_2_debug_pc,
  input  [2:0]  io_enq_6_dec_uops_2_iq_type,
  input  [9:0]  io_enq_6_dec_uops_2_fu_code,
  input  [3:0]  io_enq_6_dec_uops_2_ctrl_br_type,
  input  [1:0]  io_enq_6_dec_uops_2_ctrl_op1_sel,
  input  [2:0]  io_enq_6_dec_uops_2_ctrl_op2_sel,
  input  [2:0]  io_enq_6_dec_uops_2_ctrl_imm_sel,
  input  [3:0]  io_enq_6_dec_uops_2_ctrl_op_fcn,
  input         io_enq_6_dec_uops_2_ctrl_fcn_dw,
  input  [2:0]  io_enq_6_dec_uops_2_ctrl_csr_cmd,
  input         io_enq_6_dec_uops_2_ctrl_is_load,
  input         io_enq_6_dec_uops_2_ctrl_is_sta,
  input         io_enq_6_dec_uops_2_ctrl_is_std,
  input  [1:0]  io_enq_6_dec_uops_2_ctrl_op3_sel,
  input  [1:0]  io_enq_6_dec_uops_2_iw_state,
  input         io_enq_6_dec_uops_2_iw_p1_poisoned,
  input         io_enq_6_dec_uops_2_iw_p2_poisoned,
  input         io_enq_6_dec_uops_2_is_br,
  input         io_enq_6_dec_uops_2_is_jalr,
  input         io_enq_6_dec_uops_2_is_jal,
  input         io_enq_6_dec_uops_2_is_sfb,
  input  [11:0] io_enq_6_dec_uops_2_br_mask,
  input  [3:0]  io_enq_6_dec_uops_2_br_tag,
  input  [4:0]  io_enq_6_dec_uops_2_ftq_idx,
  input         io_enq_6_dec_uops_2_edge_inst,
  input  [5:0]  io_enq_6_dec_uops_2_pc_lob,
  input         io_enq_6_dec_uops_2_taken,
  input  [19:0] io_enq_6_dec_uops_2_imm_packed,
  input  [11:0] io_enq_6_dec_uops_2_csr_addr,
  input  [5:0]  io_enq_6_dec_uops_2_rob_idx,
  input  [4:0]  io_enq_6_dec_uops_2_ldq_idx,
  input  [4:0]  io_enq_6_dec_uops_2_stq_idx,
  input  [1:0]  io_enq_6_dec_uops_2_rxq_idx,
  input  [6:0]  io_enq_6_dec_uops_2_pdst,
  input  [6:0]  io_enq_6_dec_uops_2_prs1,
  input  [6:0]  io_enq_6_dec_uops_2_prs2,
  input  [6:0]  io_enq_6_dec_uops_2_prs3,
  input  [4:0]  io_enq_6_dec_uops_2_ppred,
  input         io_enq_6_dec_uops_2_prs1_busy,
  input         io_enq_6_dec_uops_2_prs2_busy,
  input         io_enq_6_dec_uops_2_prs3_busy,
  input         io_enq_6_dec_uops_2_ppred_busy,
  input  [6:0]  io_enq_6_dec_uops_2_stale_pdst,
  input         io_enq_6_dec_uops_2_exception,
  input  [63:0] io_enq_6_dec_uops_2_exc_cause,
  input         io_enq_6_dec_uops_2_bypassable,
  input  [4:0]  io_enq_6_dec_uops_2_mem_cmd,
  input  [1:0]  io_enq_6_dec_uops_2_mem_size,
  input         io_enq_6_dec_uops_2_mem_signed,
  input         io_enq_6_dec_uops_2_is_fence,
  input         io_enq_6_dec_uops_2_is_fencei,
  input         io_enq_6_dec_uops_2_is_amo,
  input         io_enq_6_dec_uops_2_uses_ldq,
  input         io_enq_6_dec_uops_2_uses_stq,
  input         io_enq_6_dec_uops_2_is_sys_pc2epc,
  input         io_enq_6_dec_uops_2_is_unique,
  input         io_enq_6_dec_uops_2_flush_on_commit,
  input         io_enq_6_dec_uops_2_ldst_is_rs1,
  input  [5:0]  io_enq_6_dec_uops_2_ldst,
  input  [5:0]  io_enq_6_dec_uops_2_lrs1,
  input  [5:0]  io_enq_6_dec_uops_2_lrs2,
  input  [5:0]  io_enq_6_dec_uops_2_lrs3,
  input         io_enq_6_dec_uops_2_ldst_val,
  input  [1:0]  io_enq_6_dec_uops_2_dst_rtype,
  input  [1:0]  io_enq_6_dec_uops_2_lrs1_rtype,
  input  [1:0]  io_enq_6_dec_uops_2_lrs2_rtype,
  input         io_enq_6_dec_uops_2_frs3_en,
  input         io_enq_6_dec_uops_2_fp_val,
  input         io_enq_6_dec_uops_2_fp_single,
  input         io_enq_6_dec_uops_2_xcpt_pf_if,
  input         io_enq_6_dec_uops_2_xcpt_ae_if,
  input         io_enq_6_dec_uops_2_xcpt_ma_if,
  input         io_enq_6_dec_uops_2_bp_debug_if,
  input         io_enq_6_dec_uops_2_bp_xcpt_if,
  input  [1:0]  io_enq_6_dec_uops_2_debug_fsrc,
  input  [1:0]  io_enq_6_dec_uops_2_debug_tsrc,
  input         io_enq_6_dec_uops_3_switch,
  input         io_enq_6_dec_uops_3_switch_off,
  input         io_enq_6_dec_uops_3_is_unicore,
  input  [2:0]  io_enq_6_dec_uops_3_shift,
  input  [1:0]  io_enq_6_dec_uops_3_lrs3_rtype,
  input         io_enq_6_dec_uops_3_rflag,
  input         io_enq_6_dec_uops_3_wflag,
  input  [3:0]  io_enq_6_dec_uops_3_prflag,
  input  [3:0]  io_enq_6_dec_uops_3_pwflag,
  input         io_enq_6_dec_uops_3_pflag_busy,
  input  [3:0]  io_enq_6_dec_uops_3_stale_pflag,
  input  [3:0]  io_enq_6_dec_uops_3_op1_sel,
  input  [3:0]  io_enq_6_dec_uops_3_op2_sel,
  input  [5:0]  io_enq_6_dec_uops_3_split_num,
  input  [5:0]  io_enq_6_dec_uops_3_self_index,
  input  [5:0]  io_enq_6_dec_uops_3_rob_inst_idx,
  input  [5:0]  io_enq_6_dec_uops_3_address_num,
  input  [6:0]  io_enq_6_dec_uops_3_uopc,
  input  [31:0] io_enq_6_dec_uops_3_inst,
  input  [31:0] io_enq_6_dec_uops_3_debug_inst,
  input         io_enq_6_dec_uops_3_is_rvc,
  input  [39:0] io_enq_6_dec_uops_3_debug_pc,
  input  [2:0]  io_enq_6_dec_uops_3_iq_type,
  input  [9:0]  io_enq_6_dec_uops_3_fu_code,
  input  [3:0]  io_enq_6_dec_uops_3_ctrl_br_type,
  input  [1:0]  io_enq_6_dec_uops_3_ctrl_op1_sel,
  input  [2:0]  io_enq_6_dec_uops_3_ctrl_op2_sel,
  input  [2:0]  io_enq_6_dec_uops_3_ctrl_imm_sel,
  input  [3:0]  io_enq_6_dec_uops_3_ctrl_op_fcn,
  input         io_enq_6_dec_uops_3_ctrl_fcn_dw,
  input  [2:0]  io_enq_6_dec_uops_3_ctrl_csr_cmd,
  input         io_enq_6_dec_uops_3_ctrl_is_load,
  input         io_enq_6_dec_uops_3_ctrl_is_sta,
  input         io_enq_6_dec_uops_3_ctrl_is_std,
  input  [1:0]  io_enq_6_dec_uops_3_ctrl_op3_sel,
  input  [1:0]  io_enq_6_dec_uops_3_iw_state,
  input         io_enq_6_dec_uops_3_iw_p1_poisoned,
  input         io_enq_6_dec_uops_3_iw_p2_poisoned,
  input         io_enq_6_dec_uops_3_is_br,
  input         io_enq_6_dec_uops_3_is_jalr,
  input         io_enq_6_dec_uops_3_is_jal,
  input         io_enq_6_dec_uops_3_is_sfb,
  input  [11:0] io_enq_6_dec_uops_3_br_mask,
  input  [3:0]  io_enq_6_dec_uops_3_br_tag,
  input  [4:0]  io_enq_6_dec_uops_3_ftq_idx,
  input         io_enq_6_dec_uops_3_edge_inst,
  input  [5:0]  io_enq_6_dec_uops_3_pc_lob,
  input         io_enq_6_dec_uops_3_taken,
  input  [19:0] io_enq_6_dec_uops_3_imm_packed,
  input  [11:0] io_enq_6_dec_uops_3_csr_addr,
  input  [5:0]  io_enq_6_dec_uops_3_rob_idx,
  input  [4:0]  io_enq_6_dec_uops_3_ldq_idx,
  input  [4:0]  io_enq_6_dec_uops_3_stq_idx,
  input  [1:0]  io_enq_6_dec_uops_3_rxq_idx,
  input  [6:0]  io_enq_6_dec_uops_3_pdst,
  input  [6:0]  io_enq_6_dec_uops_3_prs1,
  input  [6:0]  io_enq_6_dec_uops_3_prs2,
  input  [6:0]  io_enq_6_dec_uops_3_prs3,
  input  [4:0]  io_enq_6_dec_uops_3_ppred,
  input         io_enq_6_dec_uops_3_prs1_busy,
  input         io_enq_6_dec_uops_3_prs2_busy,
  input         io_enq_6_dec_uops_3_prs3_busy,
  input         io_enq_6_dec_uops_3_ppred_busy,
  input  [6:0]  io_enq_6_dec_uops_3_stale_pdst,
  input         io_enq_6_dec_uops_3_exception,
  input  [63:0] io_enq_6_dec_uops_3_exc_cause,
  input         io_enq_6_dec_uops_3_bypassable,
  input  [4:0]  io_enq_6_dec_uops_3_mem_cmd,
  input  [1:0]  io_enq_6_dec_uops_3_mem_size,
  input         io_enq_6_dec_uops_3_mem_signed,
  input         io_enq_6_dec_uops_3_is_fence,
  input         io_enq_6_dec_uops_3_is_fencei,
  input         io_enq_6_dec_uops_3_is_amo,
  input         io_enq_6_dec_uops_3_uses_ldq,
  input         io_enq_6_dec_uops_3_uses_stq,
  input         io_enq_6_dec_uops_3_is_sys_pc2epc,
  input         io_enq_6_dec_uops_3_is_unique,
  input         io_enq_6_dec_uops_3_flush_on_commit,
  input         io_enq_6_dec_uops_3_ldst_is_rs1,
  input  [5:0]  io_enq_6_dec_uops_3_ldst,
  input  [5:0]  io_enq_6_dec_uops_3_lrs1,
  input  [5:0]  io_enq_6_dec_uops_3_lrs2,
  input  [5:0]  io_enq_6_dec_uops_3_lrs3,
  input         io_enq_6_dec_uops_3_ldst_val,
  input  [1:0]  io_enq_6_dec_uops_3_dst_rtype,
  input  [1:0]  io_enq_6_dec_uops_3_lrs1_rtype,
  input  [1:0]  io_enq_6_dec_uops_3_lrs2_rtype,
  input         io_enq_6_dec_uops_3_frs3_en,
  input         io_enq_6_dec_uops_3_fp_val,
  input         io_enq_6_dec_uops_3_fp_single,
  input         io_enq_6_dec_uops_3_xcpt_pf_if,
  input         io_enq_6_dec_uops_3_xcpt_ae_if,
  input         io_enq_6_dec_uops_3_xcpt_ma_if,
  input         io_enq_6_dec_uops_3_bp_debug_if,
  input         io_enq_6_dec_uops_3_bp_xcpt_if,
  input  [1:0]  io_enq_6_dec_uops_3_debug_fsrc,
  input  [1:0]  io_enq_6_dec_uops_3_debug_tsrc,
  input         io_enq_6_val_mask_0,
  input         io_enq_6_val_mask_1,
  input         io_enq_6_val_mask_2,
  input         io_enq_6_val_mask_3,
  input         io_enq_7_dec_uops_0_switch,
  input         io_enq_7_dec_uops_0_switch_off,
  input         io_enq_7_dec_uops_0_is_unicore,
  input  [2:0]  io_enq_7_dec_uops_0_shift,
  input  [1:0]  io_enq_7_dec_uops_0_lrs3_rtype,
  input         io_enq_7_dec_uops_0_rflag,
  input         io_enq_7_dec_uops_0_wflag,
  input  [3:0]  io_enq_7_dec_uops_0_prflag,
  input  [3:0]  io_enq_7_dec_uops_0_pwflag,
  input         io_enq_7_dec_uops_0_pflag_busy,
  input  [3:0]  io_enq_7_dec_uops_0_stale_pflag,
  input  [3:0]  io_enq_7_dec_uops_0_op1_sel,
  input  [3:0]  io_enq_7_dec_uops_0_op2_sel,
  input  [5:0]  io_enq_7_dec_uops_0_split_num,
  input  [5:0]  io_enq_7_dec_uops_0_self_index,
  input  [5:0]  io_enq_7_dec_uops_0_rob_inst_idx,
  input  [5:0]  io_enq_7_dec_uops_0_address_num,
  input  [6:0]  io_enq_7_dec_uops_0_uopc,
  input  [31:0] io_enq_7_dec_uops_0_inst,
  input  [31:0] io_enq_7_dec_uops_0_debug_inst,
  input         io_enq_7_dec_uops_0_is_rvc,
  input  [39:0] io_enq_7_dec_uops_0_debug_pc,
  input  [2:0]  io_enq_7_dec_uops_0_iq_type,
  input  [9:0]  io_enq_7_dec_uops_0_fu_code,
  input  [3:0]  io_enq_7_dec_uops_0_ctrl_br_type,
  input  [1:0]  io_enq_7_dec_uops_0_ctrl_op1_sel,
  input  [2:0]  io_enq_7_dec_uops_0_ctrl_op2_sel,
  input  [2:0]  io_enq_7_dec_uops_0_ctrl_imm_sel,
  input  [3:0]  io_enq_7_dec_uops_0_ctrl_op_fcn,
  input         io_enq_7_dec_uops_0_ctrl_fcn_dw,
  input  [2:0]  io_enq_7_dec_uops_0_ctrl_csr_cmd,
  input         io_enq_7_dec_uops_0_ctrl_is_load,
  input         io_enq_7_dec_uops_0_ctrl_is_sta,
  input         io_enq_7_dec_uops_0_ctrl_is_std,
  input  [1:0]  io_enq_7_dec_uops_0_ctrl_op3_sel,
  input  [1:0]  io_enq_7_dec_uops_0_iw_state,
  input         io_enq_7_dec_uops_0_iw_p1_poisoned,
  input         io_enq_7_dec_uops_0_iw_p2_poisoned,
  input         io_enq_7_dec_uops_0_is_br,
  input         io_enq_7_dec_uops_0_is_jalr,
  input         io_enq_7_dec_uops_0_is_jal,
  input         io_enq_7_dec_uops_0_is_sfb,
  input  [11:0] io_enq_7_dec_uops_0_br_mask,
  input  [3:0]  io_enq_7_dec_uops_0_br_tag,
  input  [4:0]  io_enq_7_dec_uops_0_ftq_idx,
  input         io_enq_7_dec_uops_0_edge_inst,
  input  [5:0]  io_enq_7_dec_uops_0_pc_lob,
  input         io_enq_7_dec_uops_0_taken,
  input  [19:0] io_enq_7_dec_uops_0_imm_packed,
  input  [11:0] io_enq_7_dec_uops_0_csr_addr,
  input  [5:0]  io_enq_7_dec_uops_0_rob_idx,
  input  [4:0]  io_enq_7_dec_uops_0_ldq_idx,
  input  [4:0]  io_enq_7_dec_uops_0_stq_idx,
  input  [1:0]  io_enq_7_dec_uops_0_rxq_idx,
  input  [6:0]  io_enq_7_dec_uops_0_pdst,
  input  [6:0]  io_enq_7_dec_uops_0_prs1,
  input  [6:0]  io_enq_7_dec_uops_0_prs2,
  input  [6:0]  io_enq_7_dec_uops_0_prs3,
  input  [4:0]  io_enq_7_dec_uops_0_ppred,
  input         io_enq_7_dec_uops_0_prs1_busy,
  input         io_enq_7_dec_uops_0_prs2_busy,
  input         io_enq_7_dec_uops_0_prs3_busy,
  input         io_enq_7_dec_uops_0_ppred_busy,
  input  [6:0]  io_enq_7_dec_uops_0_stale_pdst,
  input         io_enq_7_dec_uops_0_exception,
  input  [63:0] io_enq_7_dec_uops_0_exc_cause,
  input         io_enq_7_dec_uops_0_bypassable,
  input  [4:0]  io_enq_7_dec_uops_0_mem_cmd,
  input  [1:0]  io_enq_7_dec_uops_0_mem_size,
  input         io_enq_7_dec_uops_0_mem_signed,
  input         io_enq_7_dec_uops_0_is_fence,
  input         io_enq_7_dec_uops_0_is_fencei,
  input         io_enq_7_dec_uops_0_is_amo,
  input         io_enq_7_dec_uops_0_uses_ldq,
  input         io_enq_7_dec_uops_0_uses_stq,
  input         io_enq_7_dec_uops_0_is_sys_pc2epc,
  input         io_enq_7_dec_uops_0_is_unique,
  input         io_enq_7_dec_uops_0_flush_on_commit,
  input         io_enq_7_dec_uops_0_ldst_is_rs1,
  input  [5:0]  io_enq_7_dec_uops_0_ldst,
  input  [5:0]  io_enq_7_dec_uops_0_lrs1,
  input  [5:0]  io_enq_7_dec_uops_0_lrs2,
  input  [5:0]  io_enq_7_dec_uops_0_lrs3,
  input         io_enq_7_dec_uops_0_ldst_val,
  input  [1:0]  io_enq_7_dec_uops_0_dst_rtype,
  input  [1:0]  io_enq_7_dec_uops_0_lrs1_rtype,
  input  [1:0]  io_enq_7_dec_uops_0_lrs2_rtype,
  input         io_enq_7_dec_uops_0_frs3_en,
  input         io_enq_7_dec_uops_0_fp_val,
  input         io_enq_7_dec_uops_0_fp_single,
  input         io_enq_7_dec_uops_0_xcpt_pf_if,
  input         io_enq_7_dec_uops_0_xcpt_ae_if,
  input         io_enq_7_dec_uops_0_xcpt_ma_if,
  input         io_enq_7_dec_uops_0_bp_debug_if,
  input         io_enq_7_dec_uops_0_bp_xcpt_if,
  input  [1:0]  io_enq_7_dec_uops_0_debug_fsrc,
  input  [1:0]  io_enq_7_dec_uops_0_debug_tsrc,
  input         io_enq_7_dec_uops_1_switch,
  input         io_enq_7_dec_uops_1_switch_off,
  input         io_enq_7_dec_uops_1_is_unicore,
  input  [2:0]  io_enq_7_dec_uops_1_shift,
  input  [1:0]  io_enq_7_dec_uops_1_lrs3_rtype,
  input         io_enq_7_dec_uops_1_rflag,
  input         io_enq_7_dec_uops_1_wflag,
  input  [3:0]  io_enq_7_dec_uops_1_prflag,
  input  [3:0]  io_enq_7_dec_uops_1_pwflag,
  input         io_enq_7_dec_uops_1_pflag_busy,
  input  [3:0]  io_enq_7_dec_uops_1_stale_pflag,
  input  [3:0]  io_enq_7_dec_uops_1_op1_sel,
  input  [3:0]  io_enq_7_dec_uops_1_op2_sel,
  input  [5:0]  io_enq_7_dec_uops_1_split_num,
  input  [5:0]  io_enq_7_dec_uops_1_self_index,
  input  [5:0]  io_enq_7_dec_uops_1_rob_inst_idx,
  input  [5:0]  io_enq_7_dec_uops_1_address_num,
  input  [6:0]  io_enq_7_dec_uops_1_uopc,
  input  [31:0] io_enq_7_dec_uops_1_inst,
  input  [31:0] io_enq_7_dec_uops_1_debug_inst,
  input         io_enq_7_dec_uops_1_is_rvc,
  input  [39:0] io_enq_7_dec_uops_1_debug_pc,
  input  [2:0]  io_enq_7_dec_uops_1_iq_type,
  input  [9:0]  io_enq_7_dec_uops_1_fu_code,
  input  [3:0]  io_enq_7_dec_uops_1_ctrl_br_type,
  input  [1:0]  io_enq_7_dec_uops_1_ctrl_op1_sel,
  input  [2:0]  io_enq_7_dec_uops_1_ctrl_op2_sel,
  input  [2:0]  io_enq_7_dec_uops_1_ctrl_imm_sel,
  input  [3:0]  io_enq_7_dec_uops_1_ctrl_op_fcn,
  input         io_enq_7_dec_uops_1_ctrl_fcn_dw,
  input  [2:0]  io_enq_7_dec_uops_1_ctrl_csr_cmd,
  input         io_enq_7_dec_uops_1_ctrl_is_load,
  input         io_enq_7_dec_uops_1_ctrl_is_sta,
  input         io_enq_7_dec_uops_1_ctrl_is_std,
  input  [1:0]  io_enq_7_dec_uops_1_ctrl_op3_sel,
  input  [1:0]  io_enq_7_dec_uops_1_iw_state,
  input         io_enq_7_dec_uops_1_iw_p1_poisoned,
  input         io_enq_7_dec_uops_1_iw_p2_poisoned,
  input         io_enq_7_dec_uops_1_is_br,
  input         io_enq_7_dec_uops_1_is_jalr,
  input         io_enq_7_dec_uops_1_is_jal,
  input         io_enq_7_dec_uops_1_is_sfb,
  input  [11:0] io_enq_7_dec_uops_1_br_mask,
  input  [3:0]  io_enq_7_dec_uops_1_br_tag,
  input  [4:0]  io_enq_7_dec_uops_1_ftq_idx,
  input         io_enq_7_dec_uops_1_edge_inst,
  input  [5:0]  io_enq_7_dec_uops_1_pc_lob,
  input         io_enq_7_dec_uops_1_taken,
  input  [19:0] io_enq_7_dec_uops_1_imm_packed,
  input  [11:0] io_enq_7_dec_uops_1_csr_addr,
  input  [5:0]  io_enq_7_dec_uops_1_rob_idx,
  input  [4:0]  io_enq_7_dec_uops_1_ldq_idx,
  input  [4:0]  io_enq_7_dec_uops_1_stq_idx,
  input  [1:0]  io_enq_7_dec_uops_1_rxq_idx,
  input  [6:0]  io_enq_7_dec_uops_1_pdst,
  input  [6:0]  io_enq_7_dec_uops_1_prs1,
  input  [6:0]  io_enq_7_dec_uops_1_prs2,
  input  [6:0]  io_enq_7_dec_uops_1_prs3,
  input  [4:0]  io_enq_7_dec_uops_1_ppred,
  input         io_enq_7_dec_uops_1_prs1_busy,
  input         io_enq_7_dec_uops_1_prs2_busy,
  input         io_enq_7_dec_uops_1_prs3_busy,
  input         io_enq_7_dec_uops_1_ppred_busy,
  input  [6:0]  io_enq_7_dec_uops_1_stale_pdst,
  input         io_enq_7_dec_uops_1_exception,
  input  [63:0] io_enq_7_dec_uops_1_exc_cause,
  input         io_enq_7_dec_uops_1_bypassable,
  input  [4:0]  io_enq_7_dec_uops_1_mem_cmd,
  input  [1:0]  io_enq_7_dec_uops_1_mem_size,
  input         io_enq_7_dec_uops_1_mem_signed,
  input         io_enq_7_dec_uops_1_is_fence,
  input         io_enq_7_dec_uops_1_is_fencei,
  input         io_enq_7_dec_uops_1_is_amo,
  input         io_enq_7_dec_uops_1_uses_ldq,
  input         io_enq_7_dec_uops_1_uses_stq,
  input         io_enq_7_dec_uops_1_is_sys_pc2epc,
  input         io_enq_7_dec_uops_1_is_unique,
  input         io_enq_7_dec_uops_1_flush_on_commit,
  input         io_enq_7_dec_uops_1_ldst_is_rs1,
  input  [5:0]  io_enq_7_dec_uops_1_ldst,
  input  [5:0]  io_enq_7_dec_uops_1_lrs1,
  input  [5:0]  io_enq_7_dec_uops_1_lrs2,
  input  [5:0]  io_enq_7_dec_uops_1_lrs3,
  input         io_enq_7_dec_uops_1_ldst_val,
  input  [1:0]  io_enq_7_dec_uops_1_dst_rtype,
  input  [1:0]  io_enq_7_dec_uops_1_lrs1_rtype,
  input  [1:0]  io_enq_7_dec_uops_1_lrs2_rtype,
  input         io_enq_7_dec_uops_1_frs3_en,
  input         io_enq_7_dec_uops_1_fp_val,
  input         io_enq_7_dec_uops_1_fp_single,
  input         io_enq_7_dec_uops_1_xcpt_pf_if,
  input         io_enq_7_dec_uops_1_xcpt_ae_if,
  input         io_enq_7_dec_uops_1_xcpt_ma_if,
  input         io_enq_7_dec_uops_1_bp_debug_if,
  input         io_enq_7_dec_uops_1_bp_xcpt_if,
  input  [1:0]  io_enq_7_dec_uops_1_debug_fsrc,
  input  [1:0]  io_enq_7_dec_uops_1_debug_tsrc,
  input         io_enq_7_dec_uops_2_switch,
  input         io_enq_7_dec_uops_2_switch_off,
  input         io_enq_7_dec_uops_2_is_unicore,
  input  [2:0]  io_enq_7_dec_uops_2_shift,
  input  [1:0]  io_enq_7_dec_uops_2_lrs3_rtype,
  input         io_enq_7_dec_uops_2_rflag,
  input         io_enq_7_dec_uops_2_wflag,
  input  [3:0]  io_enq_7_dec_uops_2_prflag,
  input  [3:0]  io_enq_7_dec_uops_2_pwflag,
  input         io_enq_7_dec_uops_2_pflag_busy,
  input  [3:0]  io_enq_7_dec_uops_2_stale_pflag,
  input  [3:0]  io_enq_7_dec_uops_2_op1_sel,
  input  [3:0]  io_enq_7_dec_uops_2_op2_sel,
  input  [5:0]  io_enq_7_dec_uops_2_split_num,
  input  [5:0]  io_enq_7_dec_uops_2_self_index,
  input  [5:0]  io_enq_7_dec_uops_2_rob_inst_idx,
  input  [5:0]  io_enq_7_dec_uops_2_address_num,
  input  [6:0]  io_enq_7_dec_uops_2_uopc,
  input  [31:0] io_enq_7_dec_uops_2_inst,
  input  [31:0] io_enq_7_dec_uops_2_debug_inst,
  input         io_enq_7_dec_uops_2_is_rvc,
  input  [39:0] io_enq_7_dec_uops_2_debug_pc,
  input  [2:0]  io_enq_7_dec_uops_2_iq_type,
  input  [9:0]  io_enq_7_dec_uops_2_fu_code,
  input  [3:0]  io_enq_7_dec_uops_2_ctrl_br_type,
  input  [1:0]  io_enq_7_dec_uops_2_ctrl_op1_sel,
  input  [2:0]  io_enq_7_dec_uops_2_ctrl_op2_sel,
  input  [2:0]  io_enq_7_dec_uops_2_ctrl_imm_sel,
  input  [3:0]  io_enq_7_dec_uops_2_ctrl_op_fcn,
  input         io_enq_7_dec_uops_2_ctrl_fcn_dw,
  input  [2:0]  io_enq_7_dec_uops_2_ctrl_csr_cmd,
  input         io_enq_7_dec_uops_2_ctrl_is_load,
  input         io_enq_7_dec_uops_2_ctrl_is_sta,
  input         io_enq_7_dec_uops_2_ctrl_is_std,
  input  [1:0]  io_enq_7_dec_uops_2_ctrl_op3_sel,
  input  [1:0]  io_enq_7_dec_uops_2_iw_state,
  input         io_enq_7_dec_uops_2_iw_p1_poisoned,
  input         io_enq_7_dec_uops_2_iw_p2_poisoned,
  input         io_enq_7_dec_uops_2_is_br,
  input         io_enq_7_dec_uops_2_is_jalr,
  input         io_enq_7_dec_uops_2_is_jal,
  input         io_enq_7_dec_uops_2_is_sfb,
  input  [11:0] io_enq_7_dec_uops_2_br_mask,
  input  [3:0]  io_enq_7_dec_uops_2_br_tag,
  input  [4:0]  io_enq_7_dec_uops_2_ftq_idx,
  input         io_enq_7_dec_uops_2_edge_inst,
  input  [5:0]  io_enq_7_dec_uops_2_pc_lob,
  input         io_enq_7_dec_uops_2_taken,
  input  [19:0] io_enq_7_dec_uops_2_imm_packed,
  input  [11:0] io_enq_7_dec_uops_2_csr_addr,
  input  [5:0]  io_enq_7_dec_uops_2_rob_idx,
  input  [4:0]  io_enq_7_dec_uops_2_ldq_idx,
  input  [4:0]  io_enq_7_dec_uops_2_stq_idx,
  input  [1:0]  io_enq_7_dec_uops_2_rxq_idx,
  input  [6:0]  io_enq_7_dec_uops_2_pdst,
  input  [6:0]  io_enq_7_dec_uops_2_prs1,
  input  [6:0]  io_enq_7_dec_uops_2_prs2,
  input  [6:0]  io_enq_7_dec_uops_2_prs3,
  input  [4:0]  io_enq_7_dec_uops_2_ppred,
  input         io_enq_7_dec_uops_2_prs1_busy,
  input         io_enq_7_dec_uops_2_prs2_busy,
  input         io_enq_7_dec_uops_2_prs3_busy,
  input         io_enq_7_dec_uops_2_ppred_busy,
  input  [6:0]  io_enq_7_dec_uops_2_stale_pdst,
  input         io_enq_7_dec_uops_2_exception,
  input  [63:0] io_enq_7_dec_uops_2_exc_cause,
  input         io_enq_7_dec_uops_2_bypassable,
  input  [4:0]  io_enq_7_dec_uops_2_mem_cmd,
  input  [1:0]  io_enq_7_dec_uops_2_mem_size,
  input         io_enq_7_dec_uops_2_mem_signed,
  input         io_enq_7_dec_uops_2_is_fence,
  input         io_enq_7_dec_uops_2_is_fencei,
  input         io_enq_7_dec_uops_2_is_amo,
  input         io_enq_7_dec_uops_2_uses_ldq,
  input         io_enq_7_dec_uops_2_uses_stq,
  input         io_enq_7_dec_uops_2_is_sys_pc2epc,
  input         io_enq_7_dec_uops_2_is_unique,
  input         io_enq_7_dec_uops_2_flush_on_commit,
  input         io_enq_7_dec_uops_2_ldst_is_rs1,
  input  [5:0]  io_enq_7_dec_uops_2_ldst,
  input  [5:0]  io_enq_7_dec_uops_2_lrs1,
  input  [5:0]  io_enq_7_dec_uops_2_lrs2,
  input  [5:0]  io_enq_7_dec_uops_2_lrs3,
  input         io_enq_7_dec_uops_2_ldst_val,
  input  [1:0]  io_enq_7_dec_uops_2_dst_rtype,
  input  [1:0]  io_enq_7_dec_uops_2_lrs1_rtype,
  input  [1:0]  io_enq_7_dec_uops_2_lrs2_rtype,
  input         io_enq_7_dec_uops_2_frs3_en,
  input         io_enq_7_dec_uops_2_fp_val,
  input         io_enq_7_dec_uops_2_fp_single,
  input         io_enq_7_dec_uops_2_xcpt_pf_if,
  input         io_enq_7_dec_uops_2_xcpt_ae_if,
  input         io_enq_7_dec_uops_2_xcpt_ma_if,
  input         io_enq_7_dec_uops_2_bp_debug_if,
  input         io_enq_7_dec_uops_2_bp_xcpt_if,
  input  [1:0]  io_enq_7_dec_uops_2_debug_fsrc,
  input  [1:0]  io_enq_7_dec_uops_2_debug_tsrc,
  input         io_enq_7_dec_uops_3_switch,
  input         io_enq_7_dec_uops_3_switch_off,
  input         io_enq_7_dec_uops_3_is_unicore,
  input  [2:0]  io_enq_7_dec_uops_3_shift,
  input  [1:0]  io_enq_7_dec_uops_3_lrs3_rtype,
  input         io_enq_7_dec_uops_3_rflag,
  input         io_enq_7_dec_uops_3_wflag,
  input  [3:0]  io_enq_7_dec_uops_3_prflag,
  input  [3:0]  io_enq_7_dec_uops_3_pwflag,
  input         io_enq_7_dec_uops_3_pflag_busy,
  input  [3:0]  io_enq_7_dec_uops_3_stale_pflag,
  input  [3:0]  io_enq_7_dec_uops_3_op1_sel,
  input  [3:0]  io_enq_7_dec_uops_3_op2_sel,
  input  [5:0]  io_enq_7_dec_uops_3_split_num,
  input  [5:0]  io_enq_7_dec_uops_3_self_index,
  input  [5:0]  io_enq_7_dec_uops_3_rob_inst_idx,
  input  [5:0]  io_enq_7_dec_uops_3_address_num,
  input  [6:0]  io_enq_7_dec_uops_3_uopc,
  input  [31:0] io_enq_7_dec_uops_3_inst,
  input  [31:0] io_enq_7_dec_uops_3_debug_inst,
  input         io_enq_7_dec_uops_3_is_rvc,
  input  [39:0] io_enq_7_dec_uops_3_debug_pc,
  input  [2:0]  io_enq_7_dec_uops_3_iq_type,
  input  [9:0]  io_enq_7_dec_uops_3_fu_code,
  input  [3:0]  io_enq_7_dec_uops_3_ctrl_br_type,
  input  [1:0]  io_enq_7_dec_uops_3_ctrl_op1_sel,
  input  [2:0]  io_enq_7_dec_uops_3_ctrl_op2_sel,
  input  [2:0]  io_enq_7_dec_uops_3_ctrl_imm_sel,
  input  [3:0]  io_enq_7_dec_uops_3_ctrl_op_fcn,
  input         io_enq_7_dec_uops_3_ctrl_fcn_dw,
  input  [2:0]  io_enq_7_dec_uops_3_ctrl_csr_cmd,
  input         io_enq_7_dec_uops_3_ctrl_is_load,
  input         io_enq_7_dec_uops_3_ctrl_is_sta,
  input         io_enq_7_dec_uops_3_ctrl_is_std,
  input  [1:0]  io_enq_7_dec_uops_3_ctrl_op3_sel,
  input  [1:0]  io_enq_7_dec_uops_3_iw_state,
  input         io_enq_7_dec_uops_3_iw_p1_poisoned,
  input         io_enq_7_dec_uops_3_iw_p2_poisoned,
  input         io_enq_7_dec_uops_3_is_br,
  input         io_enq_7_dec_uops_3_is_jalr,
  input         io_enq_7_dec_uops_3_is_jal,
  input         io_enq_7_dec_uops_3_is_sfb,
  input  [11:0] io_enq_7_dec_uops_3_br_mask,
  input  [3:0]  io_enq_7_dec_uops_3_br_tag,
  input  [4:0]  io_enq_7_dec_uops_3_ftq_idx,
  input         io_enq_7_dec_uops_3_edge_inst,
  input  [5:0]  io_enq_7_dec_uops_3_pc_lob,
  input         io_enq_7_dec_uops_3_taken,
  input  [19:0] io_enq_7_dec_uops_3_imm_packed,
  input  [11:0] io_enq_7_dec_uops_3_csr_addr,
  input  [5:0]  io_enq_7_dec_uops_3_rob_idx,
  input  [4:0]  io_enq_7_dec_uops_3_ldq_idx,
  input  [4:0]  io_enq_7_dec_uops_3_stq_idx,
  input  [1:0]  io_enq_7_dec_uops_3_rxq_idx,
  input  [6:0]  io_enq_7_dec_uops_3_pdst,
  input  [6:0]  io_enq_7_dec_uops_3_prs1,
  input  [6:0]  io_enq_7_dec_uops_3_prs2,
  input  [6:0]  io_enq_7_dec_uops_3_prs3,
  input  [4:0]  io_enq_7_dec_uops_3_ppred,
  input         io_enq_7_dec_uops_3_prs1_busy,
  input         io_enq_7_dec_uops_3_prs2_busy,
  input         io_enq_7_dec_uops_3_prs3_busy,
  input         io_enq_7_dec_uops_3_ppred_busy,
  input  [6:0]  io_enq_7_dec_uops_3_stale_pdst,
  input         io_enq_7_dec_uops_3_exception,
  input  [63:0] io_enq_7_dec_uops_3_exc_cause,
  input         io_enq_7_dec_uops_3_bypassable,
  input  [4:0]  io_enq_7_dec_uops_3_mem_cmd,
  input  [1:0]  io_enq_7_dec_uops_3_mem_size,
  input         io_enq_7_dec_uops_3_mem_signed,
  input         io_enq_7_dec_uops_3_is_fence,
  input         io_enq_7_dec_uops_3_is_fencei,
  input         io_enq_7_dec_uops_3_is_amo,
  input         io_enq_7_dec_uops_3_uses_ldq,
  input         io_enq_7_dec_uops_3_uses_stq,
  input         io_enq_7_dec_uops_3_is_sys_pc2epc,
  input         io_enq_7_dec_uops_3_is_unique,
  input         io_enq_7_dec_uops_3_flush_on_commit,
  input         io_enq_7_dec_uops_3_ldst_is_rs1,
  input  [5:0]  io_enq_7_dec_uops_3_ldst,
  input  [5:0]  io_enq_7_dec_uops_3_lrs1,
  input  [5:0]  io_enq_7_dec_uops_3_lrs2,
  input  [5:0]  io_enq_7_dec_uops_3_lrs3,
  input         io_enq_7_dec_uops_3_ldst_val,
  input  [1:0]  io_enq_7_dec_uops_3_dst_rtype,
  input  [1:0]  io_enq_7_dec_uops_3_lrs1_rtype,
  input  [1:0]  io_enq_7_dec_uops_3_lrs2_rtype,
  input         io_enq_7_dec_uops_3_frs3_en,
  input         io_enq_7_dec_uops_3_fp_val,
  input         io_enq_7_dec_uops_3_fp_single,
  input         io_enq_7_dec_uops_3_xcpt_pf_if,
  input         io_enq_7_dec_uops_3_xcpt_ae_if,
  input         io_enq_7_dec_uops_3_xcpt_ma_if,
  input         io_enq_7_dec_uops_3_bp_debug_if,
  input         io_enq_7_dec_uops_3_bp_xcpt_if,
  input  [1:0]  io_enq_7_dec_uops_3_debug_fsrc,
  input  [1:0]  io_enq_7_dec_uops_3_debug_tsrc,
  input         io_enq_7_val_mask_0,
  input         io_enq_7_val_mask_1,
  input         io_enq_7_val_mask_2,
  input         io_enq_7_val_mask_3,
  input  [4:0]  io_set_num,
  input         io_enq_valid,
  output        io_enq_ready,
  output        io_deq_tran_uops_0_switch,
  output        io_deq_tran_uops_0_switch_off,
  output        io_deq_tran_uops_0_is_unicore,
  output [2:0]  io_deq_tran_uops_0_shift,
  output [1:0]  io_deq_tran_uops_0_lrs3_rtype,
  output        io_deq_tran_uops_0_rflag,
  output        io_deq_tran_uops_0_wflag,
  output [3:0]  io_deq_tran_uops_0_prflag,
  output [3:0]  io_deq_tran_uops_0_pwflag,
  output        io_deq_tran_uops_0_pflag_busy,
  output [3:0]  io_deq_tran_uops_0_stale_pflag,
  output [3:0]  io_deq_tran_uops_0_op1_sel,
  output [3:0]  io_deq_tran_uops_0_op2_sel,
  output [5:0]  io_deq_tran_uops_0_split_num,
  output [5:0]  io_deq_tran_uops_0_self_index,
  output [5:0]  io_deq_tran_uops_0_rob_inst_idx,
  output [5:0]  io_deq_tran_uops_0_address_num,
  output [6:0]  io_deq_tran_uops_0_uopc,
  output [31:0] io_deq_tran_uops_0_inst,
  output [31:0] io_deq_tran_uops_0_debug_inst,
  output        io_deq_tran_uops_0_is_rvc,
  output [39:0] io_deq_tran_uops_0_debug_pc,
  output [2:0]  io_deq_tran_uops_0_iq_type,
  output [9:0]  io_deq_tran_uops_0_fu_code,
  output [3:0]  io_deq_tran_uops_0_ctrl_br_type,
  output [1:0]  io_deq_tran_uops_0_ctrl_op1_sel,
  output [2:0]  io_deq_tran_uops_0_ctrl_op2_sel,
  output [2:0]  io_deq_tran_uops_0_ctrl_imm_sel,
  output [3:0]  io_deq_tran_uops_0_ctrl_op_fcn,
  output        io_deq_tran_uops_0_ctrl_fcn_dw,
  output [2:0]  io_deq_tran_uops_0_ctrl_csr_cmd,
  output        io_deq_tran_uops_0_ctrl_is_load,
  output        io_deq_tran_uops_0_ctrl_is_sta,
  output        io_deq_tran_uops_0_ctrl_is_std,
  output [1:0]  io_deq_tran_uops_0_ctrl_op3_sel,
  output [1:0]  io_deq_tran_uops_0_iw_state,
  output        io_deq_tran_uops_0_iw_p1_poisoned,
  output        io_deq_tran_uops_0_iw_p2_poisoned,
  output        io_deq_tran_uops_0_is_br,
  output        io_deq_tran_uops_0_is_jalr,
  output        io_deq_tran_uops_0_is_jal,
  output        io_deq_tran_uops_0_is_sfb,
  output [11:0] io_deq_tran_uops_0_br_mask,
  output [3:0]  io_deq_tran_uops_0_br_tag,
  output [4:0]  io_deq_tran_uops_0_ftq_idx,
  output        io_deq_tran_uops_0_edge_inst,
  output [5:0]  io_deq_tran_uops_0_pc_lob,
  output        io_deq_tran_uops_0_taken,
  output [19:0] io_deq_tran_uops_0_imm_packed,
  output [11:0] io_deq_tran_uops_0_csr_addr,
  output [5:0]  io_deq_tran_uops_0_rob_idx,
  output [4:0]  io_deq_tran_uops_0_ldq_idx,
  output [4:0]  io_deq_tran_uops_0_stq_idx,
  output [1:0]  io_deq_tran_uops_0_rxq_idx,
  output [6:0]  io_deq_tran_uops_0_pdst,
  output [6:0]  io_deq_tran_uops_0_prs1,
  output [6:0]  io_deq_tran_uops_0_prs2,
  output [6:0]  io_deq_tran_uops_0_prs3,
  output [4:0]  io_deq_tran_uops_0_ppred,
  output        io_deq_tran_uops_0_prs1_busy,
  output        io_deq_tran_uops_0_prs2_busy,
  output        io_deq_tran_uops_0_prs3_busy,
  output        io_deq_tran_uops_0_ppred_busy,
  output [6:0]  io_deq_tran_uops_0_stale_pdst,
  output        io_deq_tran_uops_0_exception,
  output [63:0] io_deq_tran_uops_0_exc_cause,
  output        io_deq_tran_uops_0_bypassable,
  output [4:0]  io_deq_tran_uops_0_mem_cmd,
  output [1:0]  io_deq_tran_uops_0_mem_size,
  output        io_deq_tran_uops_0_mem_signed,
  output        io_deq_tran_uops_0_is_fence,
  output        io_deq_tran_uops_0_is_fencei,
  output        io_deq_tran_uops_0_is_amo,
  output        io_deq_tran_uops_0_uses_ldq,
  output        io_deq_tran_uops_0_uses_stq,
  output        io_deq_tran_uops_0_is_sys_pc2epc,
  output        io_deq_tran_uops_0_is_unique,
  output        io_deq_tran_uops_0_flush_on_commit,
  output        io_deq_tran_uops_0_ldst_is_rs1,
  output [5:0]  io_deq_tran_uops_0_ldst,
  output [5:0]  io_deq_tran_uops_0_lrs1,
  output [5:0]  io_deq_tran_uops_0_lrs2,
  output [5:0]  io_deq_tran_uops_0_lrs3,
  output        io_deq_tran_uops_0_ldst_val,
  output [1:0]  io_deq_tran_uops_0_dst_rtype,
  output [1:0]  io_deq_tran_uops_0_lrs1_rtype,
  output [1:0]  io_deq_tran_uops_0_lrs2_rtype,
  output        io_deq_tran_uops_0_frs3_en,
  output        io_deq_tran_uops_0_fp_val,
  output        io_deq_tran_uops_0_fp_single,
  output        io_deq_tran_uops_0_xcpt_pf_if,
  output        io_deq_tran_uops_0_xcpt_ae_if,
  output        io_deq_tran_uops_0_xcpt_ma_if,
  output        io_deq_tran_uops_0_bp_debug_if,
  output        io_deq_tran_uops_0_bp_xcpt_if,
  output [1:0]  io_deq_tran_uops_0_debug_fsrc,
  output [1:0]  io_deq_tran_uops_0_debug_tsrc,
  output        io_deq_tran_uops_1_switch,
  output        io_deq_tran_uops_1_switch_off,
  output        io_deq_tran_uops_1_is_unicore,
  output [2:0]  io_deq_tran_uops_1_shift,
  output [1:0]  io_deq_tran_uops_1_lrs3_rtype,
  output        io_deq_tran_uops_1_rflag,
  output        io_deq_tran_uops_1_wflag,
  output [3:0]  io_deq_tran_uops_1_prflag,
  output [3:0]  io_deq_tran_uops_1_pwflag,
  output        io_deq_tran_uops_1_pflag_busy,
  output [3:0]  io_deq_tran_uops_1_stale_pflag,
  output [3:0]  io_deq_tran_uops_1_op1_sel,
  output [3:0]  io_deq_tran_uops_1_op2_sel,
  output [5:0]  io_deq_tran_uops_1_split_num,
  output [5:0]  io_deq_tran_uops_1_self_index,
  output [5:0]  io_deq_tran_uops_1_rob_inst_idx,
  output [5:0]  io_deq_tran_uops_1_address_num,
  output [6:0]  io_deq_tran_uops_1_uopc,
  output [31:0] io_deq_tran_uops_1_inst,
  output [31:0] io_deq_tran_uops_1_debug_inst,
  output        io_deq_tran_uops_1_is_rvc,
  output [39:0] io_deq_tran_uops_1_debug_pc,
  output [2:0]  io_deq_tran_uops_1_iq_type,
  output [9:0]  io_deq_tran_uops_1_fu_code,
  output [3:0]  io_deq_tran_uops_1_ctrl_br_type,
  output [1:0]  io_deq_tran_uops_1_ctrl_op1_sel,
  output [2:0]  io_deq_tran_uops_1_ctrl_op2_sel,
  output [2:0]  io_deq_tran_uops_1_ctrl_imm_sel,
  output [3:0]  io_deq_tran_uops_1_ctrl_op_fcn,
  output        io_deq_tran_uops_1_ctrl_fcn_dw,
  output [2:0]  io_deq_tran_uops_1_ctrl_csr_cmd,
  output        io_deq_tran_uops_1_ctrl_is_load,
  output        io_deq_tran_uops_1_ctrl_is_sta,
  output        io_deq_tran_uops_1_ctrl_is_std,
  output [1:0]  io_deq_tran_uops_1_ctrl_op3_sel,
  output [1:0]  io_deq_tran_uops_1_iw_state,
  output        io_deq_tran_uops_1_iw_p1_poisoned,
  output        io_deq_tran_uops_1_iw_p2_poisoned,
  output        io_deq_tran_uops_1_is_br,
  output        io_deq_tran_uops_1_is_jalr,
  output        io_deq_tran_uops_1_is_jal,
  output        io_deq_tran_uops_1_is_sfb,
  output [11:0] io_deq_tran_uops_1_br_mask,
  output [3:0]  io_deq_tran_uops_1_br_tag,
  output [4:0]  io_deq_tran_uops_1_ftq_idx,
  output        io_deq_tran_uops_1_edge_inst,
  output [5:0]  io_deq_tran_uops_1_pc_lob,
  output        io_deq_tran_uops_1_taken,
  output [19:0] io_deq_tran_uops_1_imm_packed,
  output [11:0] io_deq_tran_uops_1_csr_addr,
  output [5:0]  io_deq_tran_uops_1_rob_idx,
  output [4:0]  io_deq_tran_uops_1_ldq_idx,
  output [4:0]  io_deq_tran_uops_1_stq_idx,
  output [1:0]  io_deq_tran_uops_1_rxq_idx,
  output [6:0]  io_deq_tran_uops_1_pdst,
  output [6:0]  io_deq_tran_uops_1_prs1,
  output [6:0]  io_deq_tran_uops_1_prs2,
  output [6:0]  io_deq_tran_uops_1_prs3,
  output [4:0]  io_deq_tran_uops_1_ppred,
  output        io_deq_tran_uops_1_prs1_busy,
  output        io_deq_tran_uops_1_prs2_busy,
  output        io_deq_tran_uops_1_prs3_busy,
  output        io_deq_tran_uops_1_ppred_busy,
  output [6:0]  io_deq_tran_uops_1_stale_pdst,
  output        io_deq_tran_uops_1_exception,
  output [63:0] io_deq_tran_uops_1_exc_cause,
  output        io_deq_tran_uops_1_bypassable,
  output [4:0]  io_deq_tran_uops_1_mem_cmd,
  output [1:0]  io_deq_tran_uops_1_mem_size,
  output        io_deq_tran_uops_1_mem_signed,
  output        io_deq_tran_uops_1_is_fence,
  output        io_deq_tran_uops_1_is_fencei,
  output        io_deq_tran_uops_1_is_amo,
  output        io_deq_tran_uops_1_uses_ldq,
  output        io_deq_tran_uops_1_uses_stq,
  output        io_deq_tran_uops_1_is_sys_pc2epc,
  output        io_deq_tran_uops_1_is_unique,
  output        io_deq_tran_uops_1_flush_on_commit,
  output        io_deq_tran_uops_1_ldst_is_rs1,
  output [5:0]  io_deq_tran_uops_1_ldst,
  output [5:0]  io_deq_tran_uops_1_lrs1,
  output [5:0]  io_deq_tran_uops_1_lrs2,
  output [5:0]  io_deq_tran_uops_1_lrs3,
  output        io_deq_tran_uops_1_ldst_val,
  output [1:0]  io_deq_tran_uops_1_dst_rtype,
  output [1:0]  io_deq_tran_uops_1_lrs1_rtype,
  output [1:0]  io_deq_tran_uops_1_lrs2_rtype,
  output        io_deq_tran_uops_1_frs3_en,
  output        io_deq_tran_uops_1_fp_val,
  output        io_deq_tran_uops_1_fp_single,
  output        io_deq_tran_uops_1_xcpt_pf_if,
  output        io_deq_tran_uops_1_xcpt_ae_if,
  output        io_deq_tran_uops_1_xcpt_ma_if,
  output        io_deq_tran_uops_1_bp_debug_if,
  output        io_deq_tran_uops_1_bp_xcpt_if,
  output [1:0]  io_deq_tran_uops_1_debug_fsrc,
  output [1:0]  io_deq_tran_uops_1_debug_tsrc,
  output        io_deq_tran_valids_0,
  output        io_deq_tran_valids_1,
  output        io_deq_valid,
  input         io_deq_ready,
  input         io_clear,
  input         io_isUnicoreMode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [63:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [63:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [63:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [63:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [63:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [63:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [63:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [63:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [63:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [63:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [63:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [63:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [63:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [63:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [63:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [63:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [63:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [63:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [63:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [63:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [63:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [63:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [63:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [63:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [63:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [63:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [63:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [63:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [63:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1549;
  reg [31:0] _RAND_1550;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [31:0] _RAND_1554;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1557;
  reg [31:0] _RAND_1558;
  reg [31:0] _RAND_1559;
  reg [31:0] _RAND_1560;
  reg [31:0] _RAND_1561;
  reg [31:0] _RAND_1562;
  reg [31:0] _RAND_1563;
  reg [31:0] _RAND_1564;
  reg [31:0] _RAND_1565;
  reg [31:0] _RAND_1566;
  reg [31:0] _RAND_1567;
  reg [31:0] _RAND_1568;
  reg [31:0] _RAND_1569;
  reg [31:0] _RAND_1570;
  reg [31:0] _RAND_1571;
  reg [31:0] _RAND_1572;
  reg [31:0] _RAND_1573;
  reg [31:0] _RAND_1574;
  reg [31:0] _RAND_1575;
  reg [31:0] _RAND_1576;
  reg [31:0] _RAND_1577;
  reg [31:0] _RAND_1578;
  reg [31:0] _RAND_1579;
  reg [31:0] _RAND_1580;
  reg [31:0] _RAND_1581;
  reg [31:0] _RAND_1582;
  reg [31:0] _RAND_1583;
  reg [31:0] _RAND_1584;
  reg [31:0] _RAND_1585;
  reg [31:0] _RAND_1586;
  reg [31:0] _RAND_1587;
  reg [31:0] _RAND_1588;
  reg [63:0] _RAND_1589;
  reg [31:0] _RAND_1590;
  reg [31:0] _RAND_1591;
  reg [31:0] _RAND_1592;
  reg [31:0] _RAND_1593;
  reg [31:0] _RAND_1594;
  reg [31:0] _RAND_1595;
  reg [31:0] _RAND_1596;
  reg [31:0] _RAND_1597;
  reg [31:0] _RAND_1598;
  reg [31:0] _RAND_1599;
  reg [31:0] _RAND_1600;
  reg [31:0] _RAND_1601;
  reg [31:0] _RAND_1602;
  reg [31:0] _RAND_1603;
  reg [31:0] _RAND_1604;
  reg [31:0] _RAND_1605;
  reg [31:0] _RAND_1606;
  reg [31:0] _RAND_1607;
  reg [31:0] _RAND_1608;
  reg [31:0] _RAND_1609;
  reg [31:0] _RAND_1610;
  reg [31:0] _RAND_1611;
  reg [31:0] _RAND_1612;
  reg [31:0] _RAND_1613;
  reg [31:0] _RAND_1614;
  reg [31:0] _RAND_1615;
  reg [31:0] _RAND_1616;
  reg [31:0] _RAND_1617;
  reg [31:0] _RAND_1618;
  reg [31:0] _RAND_1619;
  reg [31:0] _RAND_1620;
  reg [31:0] _RAND_1621;
  reg [31:0] _RAND_1622;
  reg [31:0] _RAND_1623;
  reg [31:0] _RAND_1624;
  reg [31:0] _RAND_1625;
  reg [31:0] _RAND_1626;
  reg [31:0] _RAND_1627;
  reg [31:0] _RAND_1628;
  reg [31:0] _RAND_1629;
  reg [31:0] _RAND_1630;
  reg [31:0] _RAND_1631;
  reg [31:0] _RAND_1632;
  reg [63:0] _RAND_1633;
  reg [31:0] _RAND_1634;
  reg [31:0] _RAND_1635;
  reg [31:0] _RAND_1636;
  reg [31:0] _RAND_1637;
  reg [31:0] _RAND_1638;
  reg [31:0] _RAND_1639;
  reg [31:0] _RAND_1640;
  reg [31:0] _RAND_1641;
  reg [31:0] _RAND_1642;
  reg [31:0] _RAND_1643;
  reg [31:0] _RAND_1644;
  reg [31:0] _RAND_1645;
  reg [31:0] _RAND_1646;
  reg [31:0] _RAND_1647;
  reg [31:0] _RAND_1648;
  reg [31:0] _RAND_1649;
  reg [31:0] _RAND_1650;
  reg [31:0] _RAND_1651;
  reg [31:0] _RAND_1652;
  reg [31:0] _RAND_1653;
  reg [31:0] _RAND_1654;
  reg [31:0] _RAND_1655;
  reg [31:0] _RAND_1656;
  reg [31:0] _RAND_1657;
  reg [31:0] _RAND_1658;
  reg [31:0] _RAND_1659;
  reg [31:0] _RAND_1660;
  reg [31:0] _RAND_1661;
  reg [31:0] _RAND_1662;
  reg [31:0] _RAND_1663;
  reg [31:0] _RAND_1664;
  reg [31:0] _RAND_1665;
  reg [31:0] _RAND_1666;
  reg [31:0] _RAND_1667;
  reg [31:0] _RAND_1668;
  reg [31:0] _RAND_1669;
  reg [31:0] _RAND_1670;
  reg [31:0] _RAND_1671;
  reg [31:0] _RAND_1672;
  reg [31:0] _RAND_1673;
  reg [31:0] _RAND_1674;
  reg [31:0] _RAND_1675;
  reg [31:0] _RAND_1676;
  reg [31:0] _RAND_1677;
  reg [31:0] _RAND_1678;
  reg [31:0] _RAND_1679;
  reg [31:0] _RAND_1680;
  reg [31:0] _RAND_1681;
  reg [31:0] _RAND_1682;
  reg [31:0] _RAND_1683;
  reg [31:0] _RAND_1684;
  reg [31:0] _RAND_1685;
  reg [63:0] _RAND_1686;
  reg [31:0] _RAND_1687;
  reg [31:0] _RAND_1688;
  reg [31:0] _RAND_1689;
  reg [31:0] _RAND_1690;
  reg [31:0] _RAND_1691;
  reg [31:0] _RAND_1692;
  reg [31:0] _RAND_1693;
  reg [31:0] _RAND_1694;
  reg [31:0] _RAND_1695;
  reg [31:0] _RAND_1696;
  reg [31:0] _RAND_1697;
  reg [31:0] _RAND_1698;
  reg [31:0] _RAND_1699;
  reg [31:0] _RAND_1700;
  reg [31:0] _RAND_1701;
  reg [31:0] _RAND_1702;
  reg [31:0] _RAND_1703;
  reg [31:0] _RAND_1704;
  reg [31:0] _RAND_1705;
  reg [31:0] _RAND_1706;
  reg [31:0] _RAND_1707;
  reg [31:0] _RAND_1708;
  reg [31:0] _RAND_1709;
  reg [31:0] _RAND_1710;
  reg [31:0] _RAND_1711;
  reg [31:0] _RAND_1712;
  reg [31:0] _RAND_1713;
  reg [31:0] _RAND_1714;
  reg [31:0] _RAND_1715;
  reg [31:0] _RAND_1716;
  reg [31:0] _RAND_1717;
  reg [31:0] _RAND_1718;
  reg [31:0] _RAND_1719;
  reg [31:0] _RAND_1720;
  reg [31:0] _RAND_1721;
  reg [31:0] _RAND_1722;
  reg [31:0] _RAND_1723;
  reg [31:0] _RAND_1724;
  reg [31:0] _RAND_1725;
  reg [31:0] _RAND_1726;
  reg [31:0] _RAND_1727;
  reg [31:0] _RAND_1728;
  reg [31:0] _RAND_1729;
  reg [63:0] _RAND_1730;
  reg [31:0] _RAND_1731;
  reg [31:0] _RAND_1732;
  reg [31:0] _RAND_1733;
  reg [31:0] _RAND_1734;
  reg [31:0] _RAND_1735;
  reg [31:0] _RAND_1736;
  reg [31:0] _RAND_1737;
  reg [31:0] _RAND_1738;
  reg [31:0] _RAND_1739;
  reg [31:0] _RAND_1740;
  reg [31:0] _RAND_1741;
  reg [31:0] _RAND_1742;
  reg [31:0] _RAND_1743;
  reg [31:0] _RAND_1744;
  reg [31:0] _RAND_1745;
  reg [31:0] _RAND_1746;
  reg [31:0] _RAND_1747;
  reg [31:0] _RAND_1748;
  reg [31:0] _RAND_1749;
  reg [31:0] _RAND_1750;
  reg [31:0] _RAND_1751;
  reg [31:0] _RAND_1752;
  reg [31:0] _RAND_1753;
  reg [31:0] _RAND_1754;
  reg [31:0] _RAND_1755;
  reg [31:0] _RAND_1756;
  reg [31:0] _RAND_1757;
  reg [31:0] _RAND_1758;
  reg [31:0] _RAND_1759;
  reg [31:0] _RAND_1760;
  reg [31:0] _RAND_1761;
  reg [31:0] _RAND_1762;
  reg [31:0] _RAND_1763;
  reg [31:0] _RAND_1764;
  reg [31:0] _RAND_1765;
  reg [31:0] _RAND_1766;
  reg [31:0] _RAND_1767;
  reg [31:0] _RAND_1768;
  reg [31:0] _RAND_1769;
  reg [31:0] _RAND_1770;
  reg [31:0] _RAND_1771;
  reg [31:0] _RAND_1772;
  reg [31:0] _RAND_1773;
  reg [31:0] _RAND_1774;
  reg [31:0] _RAND_1775;
  reg [31:0] _RAND_1776;
  reg [31:0] _RAND_1777;
  reg [31:0] _RAND_1778;
  reg [31:0] _RAND_1779;
  reg [31:0] _RAND_1780;
  reg [31:0] _RAND_1781;
  reg [31:0] _RAND_1782;
  reg [63:0] _RAND_1783;
  reg [31:0] _RAND_1784;
  reg [31:0] _RAND_1785;
  reg [31:0] _RAND_1786;
  reg [31:0] _RAND_1787;
  reg [31:0] _RAND_1788;
  reg [31:0] _RAND_1789;
  reg [31:0] _RAND_1790;
  reg [31:0] _RAND_1791;
  reg [31:0] _RAND_1792;
  reg [31:0] _RAND_1793;
  reg [31:0] _RAND_1794;
  reg [31:0] _RAND_1795;
  reg [31:0] _RAND_1796;
  reg [31:0] _RAND_1797;
  reg [31:0] _RAND_1798;
  reg [31:0] _RAND_1799;
  reg [31:0] _RAND_1800;
  reg [31:0] _RAND_1801;
  reg [31:0] _RAND_1802;
  reg [31:0] _RAND_1803;
  reg [31:0] _RAND_1804;
  reg [31:0] _RAND_1805;
  reg [31:0] _RAND_1806;
  reg [31:0] _RAND_1807;
  reg [31:0] _RAND_1808;
  reg [31:0] _RAND_1809;
  reg [31:0] _RAND_1810;
  reg [31:0] _RAND_1811;
  reg [31:0] _RAND_1812;
  reg [31:0] _RAND_1813;
  reg [31:0] _RAND_1814;
  reg [31:0] _RAND_1815;
  reg [31:0] _RAND_1816;
  reg [31:0] _RAND_1817;
  reg [31:0] _RAND_1818;
  reg [31:0] _RAND_1819;
  reg [31:0] _RAND_1820;
  reg [31:0] _RAND_1821;
  reg [31:0] _RAND_1822;
  reg [31:0] _RAND_1823;
  reg [31:0] _RAND_1824;
  reg [31:0] _RAND_1825;
  reg [31:0] _RAND_1826;
  reg [63:0] _RAND_1827;
  reg [31:0] _RAND_1828;
  reg [31:0] _RAND_1829;
  reg [31:0] _RAND_1830;
  reg [31:0] _RAND_1831;
  reg [31:0] _RAND_1832;
  reg [31:0] _RAND_1833;
  reg [31:0] _RAND_1834;
  reg [31:0] _RAND_1835;
  reg [31:0] _RAND_1836;
  reg [31:0] _RAND_1837;
  reg [31:0] _RAND_1838;
  reg [31:0] _RAND_1839;
  reg [31:0] _RAND_1840;
  reg [31:0] _RAND_1841;
  reg [31:0] _RAND_1842;
  reg [31:0] _RAND_1843;
  reg [31:0] _RAND_1844;
  reg [31:0] _RAND_1845;
  reg [31:0] _RAND_1846;
  reg [31:0] _RAND_1847;
  reg [31:0] _RAND_1848;
  reg [31:0] _RAND_1849;
  reg [31:0] _RAND_1850;
  reg [31:0] _RAND_1851;
  reg [31:0] _RAND_1852;
  reg [31:0] _RAND_1853;
  reg [31:0] _RAND_1854;
  reg [31:0] _RAND_1855;
  reg [31:0] _RAND_1856;
  reg [31:0] _RAND_1857;
  reg [31:0] _RAND_1858;
  reg [31:0] _RAND_1859;
  reg [31:0] _RAND_1860;
  reg [31:0] _RAND_1861;
  reg [31:0] _RAND_1862;
  reg [31:0] _RAND_1863;
  reg [31:0] _RAND_1864;
  reg [31:0] _RAND_1865;
  reg [31:0] _RAND_1866;
  reg [31:0] _RAND_1867;
  reg [31:0] _RAND_1868;
  reg [31:0] _RAND_1869;
  reg [31:0] _RAND_1870;
  reg [31:0] _RAND_1871;
  reg [31:0] _RAND_1872;
  reg [31:0] _RAND_1873;
  reg [31:0] _RAND_1874;
  reg [31:0] _RAND_1875;
  reg [31:0] _RAND_1876;
  reg [31:0] _RAND_1877;
  reg [31:0] _RAND_1878;
  reg [31:0] _RAND_1879;
  reg [63:0] _RAND_1880;
  reg [31:0] _RAND_1881;
  reg [31:0] _RAND_1882;
  reg [31:0] _RAND_1883;
  reg [31:0] _RAND_1884;
  reg [31:0] _RAND_1885;
  reg [31:0] _RAND_1886;
  reg [31:0] _RAND_1887;
  reg [31:0] _RAND_1888;
  reg [31:0] _RAND_1889;
  reg [31:0] _RAND_1890;
  reg [31:0] _RAND_1891;
  reg [31:0] _RAND_1892;
  reg [31:0] _RAND_1893;
  reg [31:0] _RAND_1894;
  reg [31:0] _RAND_1895;
  reg [31:0] _RAND_1896;
  reg [31:0] _RAND_1897;
  reg [31:0] _RAND_1898;
  reg [31:0] _RAND_1899;
  reg [31:0] _RAND_1900;
  reg [31:0] _RAND_1901;
  reg [31:0] _RAND_1902;
  reg [31:0] _RAND_1903;
  reg [31:0] _RAND_1904;
  reg [31:0] _RAND_1905;
  reg [31:0] _RAND_1906;
  reg [31:0] _RAND_1907;
  reg [31:0] _RAND_1908;
  reg [31:0] _RAND_1909;
  reg [31:0] _RAND_1910;
  reg [31:0] _RAND_1911;
  reg [31:0] _RAND_1912;
  reg [31:0] _RAND_1913;
  reg [31:0] _RAND_1914;
  reg [31:0] _RAND_1915;
  reg [31:0] _RAND_1916;
  reg [31:0] _RAND_1917;
  reg [31:0] _RAND_1918;
  reg [31:0] _RAND_1919;
  reg [31:0] _RAND_1920;
  reg [31:0] _RAND_1921;
  reg [31:0] _RAND_1922;
  reg [31:0] _RAND_1923;
  reg [63:0] _RAND_1924;
  reg [31:0] _RAND_1925;
  reg [31:0] _RAND_1926;
  reg [31:0] _RAND_1927;
  reg [31:0] _RAND_1928;
  reg [31:0] _RAND_1929;
  reg [31:0] _RAND_1930;
  reg [31:0] _RAND_1931;
  reg [31:0] _RAND_1932;
  reg [31:0] _RAND_1933;
  reg [31:0] _RAND_1934;
  reg [31:0] _RAND_1935;
  reg [31:0] _RAND_1936;
  reg [31:0] _RAND_1937;
  reg [31:0] _RAND_1938;
  reg [31:0] _RAND_1939;
  reg [31:0] _RAND_1940;
  reg [31:0] _RAND_1941;
  reg [31:0] _RAND_1942;
  reg [31:0] _RAND_1943;
  reg [31:0] _RAND_1944;
  reg [31:0] _RAND_1945;
  reg [31:0] _RAND_1946;
  reg [31:0] _RAND_1947;
  reg [31:0] _RAND_1948;
  reg [31:0] _RAND_1949;
  reg [31:0] _RAND_1950;
  reg [31:0] _RAND_1951;
  reg [31:0] _RAND_1952;
  reg [31:0] _RAND_1953;
  reg [31:0] _RAND_1954;
  reg [31:0] _RAND_1955;
  reg [31:0] _RAND_1956;
  reg [31:0] _RAND_1957;
  reg [31:0] _RAND_1958;
  reg [31:0] _RAND_1959;
  reg [31:0] _RAND_1960;
  reg [31:0] _RAND_1961;
  reg [31:0] _RAND_1962;
  reg [31:0] _RAND_1963;
  reg [31:0] _RAND_1964;
  reg [31:0] _RAND_1965;
  reg [31:0] _RAND_1966;
  reg [31:0] _RAND_1967;
  reg [31:0] _RAND_1968;
  reg [31:0] _RAND_1969;
  reg [31:0] _RAND_1970;
  reg [31:0] _RAND_1971;
  reg [31:0] _RAND_1972;
  reg [31:0] _RAND_1973;
  reg [31:0] _RAND_1974;
  reg [31:0] _RAND_1975;
  reg [31:0] _RAND_1976;
  reg [31:0] _RAND_1977;
  reg [31:0] _RAND_1978;
  reg [31:0] _RAND_1979;
  reg [31:0] _RAND_1980;
  reg [63:0] _RAND_1981;
  reg [31:0] _RAND_1982;
  reg [31:0] _RAND_1983;
  reg [31:0] _RAND_1984;
  reg [31:0] _RAND_1985;
  reg [31:0] _RAND_1986;
  reg [31:0] _RAND_1987;
  reg [31:0] _RAND_1988;
  reg [31:0] _RAND_1989;
  reg [31:0] _RAND_1990;
  reg [31:0] _RAND_1991;
  reg [31:0] _RAND_1992;
  reg [31:0] _RAND_1993;
  reg [31:0] _RAND_1994;
  reg [31:0] _RAND_1995;
  reg [31:0] _RAND_1996;
  reg [31:0] _RAND_1997;
  reg [31:0] _RAND_1998;
  reg [31:0] _RAND_1999;
  reg [31:0] _RAND_2000;
  reg [31:0] _RAND_2001;
  reg [31:0] _RAND_2002;
  reg [31:0] _RAND_2003;
  reg [31:0] _RAND_2004;
  reg [31:0] _RAND_2005;
  reg [31:0] _RAND_2006;
  reg [31:0] _RAND_2007;
  reg [31:0] _RAND_2008;
  reg [31:0] _RAND_2009;
  reg [31:0] _RAND_2010;
  reg [31:0] _RAND_2011;
  reg [31:0] _RAND_2012;
  reg [31:0] _RAND_2013;
  reg [31:0] _RAND_2014;
  reg [31:0] _RAND_2015;
  reg [31:0] _RAND_2016;
  reg [31:0] _RAND_2017;
  reg [31:0] _RAND_2018;
  reg [31:0] _RAND_2019;
  reg [31:0] _RAND_2020;
  reg [31:0] _RAND_2021;
  reg [31:0] _RAND_2022;
  reg [31:0] _RAND_2023;
  reg [31:0] _RAND_2024;
  reg [63:0] _RAND_2025;
  reg [31:0] _RAND_2026;
  reg [31:0] _RAND_2027;
  reg [31:0] _RAND_2028;
  reg [31:0] _RAND_2029;
  reg [31:0] _RAND_2030;
  reg [31:0] _RAND_2031;
  reg [31:0] _RAND_2032;
  reg [31:0] _RAND_2033;
  reg [31:0] _RAND_2034;
  reg [31:0] _RAND_2035;
  reg [31:0] _RAND_2036;
  reg [31:0] _RAND_2037;
  reg [31:0] _RAND_2038;
  reg [31:0] _RAND_2039;
  reg [31:0] _RAND_2040;
  reg [31:0] _RAND_2041;
  reg [31:0] _RAND_2042;
  reg [31:0] _RAND_2043;
  reg [31:0] _RAND_2044;
  reg [31:0] _RAND_2045;
  reg [31:0] _RAND_2046;
  reg [31:0] _RAND_2047;
  reg [31:0] _RAND_2048;
  reg [31:0] _RAND_2049;
  reg [31:0] _RAND_2050;
  reg [31:0] _RAND_2051;
  reg [31:0] _RAND_2052;
  reg [31:0] _RAND_2053;
  reg [31:0] _RAND_2054;
  reg [31:0] _RAND_2055;
  reg [31:0] _RAND_2056;
  reg [31:0] _RAND_2057;
  reg [31:0] _RAND_2058;
  reg [31:0] _RAND_2059;
  reg [31:0] _RAND_2060;
  reg [31:0] _RAND_2061;
  reg [31:0] _RAND_2062;
  reg [31:0] _RAND_2063;
  reg [31:0] _RAND_2064;
  reg [31:0] _RAND_2065;
  reg [31:0] _RAND_2066;
  reg [31:0] _RAND_2067;
  reg [31:0] _RAND_2068;
  reg [31:0] _RAND_2069;
  reg [31:0] _RAND_2070;
  reg [31:0] _RAND_2071;
  reg [31:0] _RAND_2072;
  reg [31:0] _RAND_2073;
  reg [31:0] _RAND_2074;
  reg [31:0] _RAND_2075;
  reg [31:0] _RAND_2076;
  reg [31:0] _RAND_2077;
  reg [63:0] _RAND_2078;
  reg [31:0] _RAND_2079;
  reg [31:0] _RAND_2080;
  reg [31:0] _RAND_2081;
  reg [31:0] _RAND_2082;
  reg [31:0] _RAND_2083;
  reg [31:0] _RAND_2084;
  reg [31:0] _RAND_2085;
  reg [31:0] _RAND_2086;
  reg [31:0] _RAND_2087;
  reg [31:0] _RAND_2088;
  reg [31:0] _RAND_2089;
  reg [31:0] _RAND_2090;
  reg [31:0] _RAND_2091;
  reg [31:0] _RAND_2092;
  reg [31:0] _RAND_2093;
  reg [31:0] _RAND_2094;
  reg [31:0] _RAND_2095;
  reg [31:0] _RAND_2096;
  reg [31:0] _RAND_2097;
  reg [31:0] _RAND_2098;
  reg [31:0] _RAND_2099;
  reg [31:0] _RAND_2100;
  reg [31:0] _RAND_2101;
  reg [31:0] _RAND_2102;
  reg [31:0] _RAND_2103;
  reg [31:0] _RAND_2104;
  reg [31:0] _RAND_2105;
  reg [31:0] _RAND_2106;
  reg [31:0] _RAND_2107;
  reg [31:0] _RAND_2108;
  reg [31:0] _RAND_2109;
  reg [31:0] _RAND_2110;
  reg [31:0] _RAND_2111;
  reg [31:0] _RAND_2112;
  reg [31:0] _RAND_2113;
  reg [31:0] _RAND_2114;
  reg [31:0] _RAND_2115;
  reg [31:0] _RAND_2116;
  reg [31:0] _RAND_2117;
  reg [31:0] _RAND_2118;
  reg [31:0] _RAND_2119;
  reg [31:0] _RAND_2120;
  reg [31:0] _RAND_2121;
  reg [63:0] _RAND_2122;
  reg [31:0] _RAND_2123;
  reg [31:0] _RAND_2124;
  reg [31:0] _RAND_2125;
  reg [31:0] _RAND_2126;
  reg [31:0] _RAND_2127;
  reg [31:0] _RAND_2128;
  reg [31:0] _RAND_2129;
  reg [31:0] _RAND_2130;
  reg [31:0] _RAND_2131;
  reg [31:0] _RAND_2132;
  reg [31:0] _RAND_2133;
  reg [31:0] _RAND_2134;
  reg [31:0] _RAND_2135;
  reg [31:0] _RAND_2136;
  reg [31:0] _RAND_2137;
  reg [31:0] _RAND_2138;
  reg [31:0] _RAND_2139;
  reg [31:0] _RAND_2140;
  reg [31:0] _RAND_2141;
  reg [31:0] _RAND_2142;
  reg [31:0] _RAND_2143;
  reg [31:0] _RAND_2144;
  reg [31:0] _RAND_2145;
  reg [31:0] _RAND_2146;
  reg [31:0] _RAND_2147;
  reg [31:0] _RAND_2148;
  reg [31:0] _RAND_2149;
  reg [31:0] _RAND_2150;
  reg [31:0] _RAND_2151;
  reg [31:0] _RAND_2152;
  reg [31:0] _RAND_2153;
  reg [31:0] _RAND_2154;
  reg [31:0] _RAND_2155;
  reg [31:0] _RAND_2156;
  reg [31:0] _RAND_2157;
  reg [31:0] _RAND_2158;
  reg [31:0] _RAND_2159;
  reg [31:0] _RAND_2160;
  reg [31:0] _RAND_2161;
  reg [31:0] _RAND_2162;
  reg [31:0] _RAND_2163;
  reg [31:0] _RAND_2164;
  reg [31:0] _RAND_2165;
  reg [31:0] _RAND_2166;
  reg [31:0] _RAND_2167;
  reg [31:0] _RAND_2168;
  reg [31:0] _RAND_2169;
  reg [31:0] _RAND_2170;
  reg [31:0] _RAND_2171;
  reg [31:0] _RAND_2172;
  reg [31:0] _RAND_2173;
  reg [31:0] _RAND_2174;
  reg [63:0] _RAND_2175;
  reg [31:0] _RAND_2176;
  reg [31:0] _RAND_2177;
  reg [31:0] _RAND_2178;
  reg [31:0] _RAND_2179;
  reg [31:0] _RAND_2180;
  reg [31:0] _RAND_2181;
  reg [31:0] _RAND_2182;
  reg [31:0] _RAND_2183;
  reg [31:0] _RAND_2184;
  reg [31:0] _RAND_2185;
  reg [31:0] _RAND_2186;
  reg [31:0] _RAND_2187;
  reg [31:0] _RAND_2188;
  reg [31:0] _RAND_2189;
  reg [31:0] _RAND_2190;
  reg [31:0] _RAND_2191;
  reg [31:0] _RAND_2192;
  reg [31:0] _RAND_2193;
  reg [31:0] _RAND_2194;
  reg [31:0] _RAND_2195;
  reg [31:0] _RAND_2196;
  reg [31:0] _RAND_2197;
  reg [31:0] _RAND_2198;
  reg [31:0] _RAND_2199;
  reg [31:0] _RAND_2200;
  reg [31:0] _RAND_2201;
  reg [31:0] _RAND_2202;
  reg [31:0] _RAND_2203;
  reg [31:0] _RAND_2204;
  reg [31:0] _RAND_2205;
  reg [31:0] _RAND_2206;
  reg [31:0] _RAND_2207;
  reg [31:0] _RAND_2208;
  reg [31:0] _RAND_2209;
  reg [31:0] _RAND_2210;
  reg [31:0] _RAND_2211;
  reg [31:0] _RAND_2212;
  reg [31:0] _RAND_2213;
  reg [31:0] _RAND_2214;
  reg [31:0] _RAND_2215;
  reg [31:0] _RAND_2216;
  reg [31:0] _RAND_2217;
  reg [31:0] _RAND_2218;
  reg [63:0] _RAND_2219;
  reg [31:0] _RAND_2220;
  reg [31:0] _RAND_2221;
  reg [31:0] _RAND_2222;
  reg [31:0] _RAND_2223;
  reg [31:0] _RAND_2224;
  reg [31:0] _RAND_2225;
  reg [31:0] _RAND_2226;
  reg [31:0] _RAND_2227;
  reg [31:0] _RAND_2228;
  reg [31:0] _RAND_2229;
  reg [31:0] _RAND_2230;
  reg [31:0] _RAND_2231;
  reg [31:0] _RAND_2232;
  reg [31:0] _RAND_2233;
  reg [31:0] _RAND_2234;
  reg [31:0] _RAND_2235;
  reg [31:0] _RAND_2236;
  reg [31:0] _RAND_2237;
  reg [31:0] _RAND_2238;
  reg [31:0] _RAND_2239;
  reg [31:0] _RAND_2240;
  reg [31:0] _RAND_2241;
  reg [31:0] _RAND_2242;
  reg [31:0] _RAND_2243;
  reg [31:0] _RAND_2244;
  reg [31:0] _RAND_2245;
  reg [31:0] _RAND_2246;
  reg [31:0] _RAND_2247;
  reg [31:0] _RAND_2248;
  reg [31:0] _RAND_2249;
  reg [31:0] _RAND_2250;
  reg [31:0] _RAND_2251;
  reg [31:0] _RAND_2252;
  reg [31:0] _RAND_2253;
  reg [31:0] _RAND_2254;
  reg [31:0] _RAND_2255;
  reg [31:0] _RAND_2256;
  reg [31:0] _RAND_2257;
  reg [31:0] _RAND_2258;
  reg [31:0] _RAND_2259;
  reg [31:0] _RAND_2260;
  reg [31:0] _RAND_2261;
  reg [31:0] _RAND_2262;
  reg [31:0] _RAND_2263;
  reg [31:0] _RAND_2264;
  reg [31:0] _RAND_2265;
  reg [31:0] _RAND_2266;
  reg [31:0] _RAND_2267;
  reg [31:0] _RAND_2268;
  reg [31:0] _RAND_2269;
  reg [31:0] _RAND_2270;
  reg [31:0] _RAND_2271;
  reg [63:0] _RAND_2272;
  reg [31:0] _RAND_2273;
  reg [31:0] _RAND_2274;
  reg [31:0] _RAND_2275;
  reg [31:0] _RAND_2276;
  reg [31:0] _RAND_2277;
  reg [31:0] _RAND_2278;
  reg [31:0] _RAND_2279;
  reg [31:0] _RAND_2280;
  reg [31:0] _RAND_2281;
  reg [31:0] _RAND_2282;
  reg [31:0] _RAND_2283;
  reg [31:0] _RAND_2284;
  reg [31:0] _RAND_2285;
  reg [31:0] _RAND_2286;
  reg [31:0] _RAND_2287;
  reg [31:0] _RAND_2288;
  reg [31:0] _RAND_2289;
  reg [31:0] _RAND_2290;
  reg [31:0] _RAND_2291;
  reg [31:0] _RAND_2292;
  reg [31:0] _RAND_2293;
  reg [31:0] _RAND_2294;
  reg [31:0] _RAND_2295;
  reg [31:0] _RAND_2296;
  reg [31:0] _RAND_2297;
  reg [31:0] _RAND_2298;
  reg [31:0] _RAND_2299;
  reg [31:0] _RAND_2300;
  reg [31:0] _RAND_2301;
  reg [31:0] _RAND_2302;
  reg [31:0] _RAND_2303;
  reg [31:0] _RAND_2304;
  reg [31:0] _RAND_2305;
  reg [31:0] _RAND_2306;
  reg [31:0] _RAND_2307;
  reg [31:0] _RAND_2308;
  reg [31:0] _RAND_2309;
  reg [31:0] _RAND_2310;
  reg [31:0] _RAND_2311;
  reg [31:0] _RAND_2312;
  reg [31:0] _RAND_2313;
  reg [31:0] _RAND_2314;
  reg [31:0] _RAND_2315;
  reg [63:0] _RAND_2316;
  reg [31:0] _RAND_2317;
  reg [31:0] _RAND_2318;
  reg [31:0] _RAND_2319;
  reg [31:0] _RAND_2320;
  reg [31:0] _RAND_2321;
  reg [31:0] _RAND_2322;
  reg [31:0] _RAND_2323;
  reg [31:0] _RAND_2324;
  reg [31:0] _RAND_2325;
  reg [31:0] _RAND_2326;
  reg [31:0] _RAND_2327;
  reg [31:0] _RAND_2328;
  reg [31:0] _RAND_2329;
  reg [31:0] _RAND_2330;
  reg [31:0] _RAND_2331;
  reg [31:0] _RAND_2332;
  reg [31:0] _RAND_2333;
  reg [31:0] _RAND_2334;
  reg [31:0] _RAND_2335;
  reg [31:0] _RAND_2336;
  reg [31:0] _RAND_2337;
  reg [31:0] _RAND_2338;
  reg [31:0] _RAND_2339;
  reg [31:0] _RAND_2340;
  reg [31:0] _RAND_2341;
  reg [31:0] _RAND_2342;
  reg [31:0] _RAND_2343;
  reg [31:0] _RAND_2344;
  reg [31:0] _RAND_2345;
  reg [31:0] _RAND_2346;
  reg [31:0] _RAND_2347;
  reg [31:0] _RAND_2348;
  reg [31:0] _RAND_2349;
  reg [31:0] _RAND_2350;
  reg [31:0] _RAND_2351;
  reg [31:0] _RAND_2352;
  reg [31:0] _RAND_2353;
  reg [31:0] _RAND_2354;
  reg [31:0] _RAND_2355;
  reg [31:0] _RAND_2356;
  reg [31:0] _RAND_2357;
  reg [31:0] _RAND_2358;
  reg [31:0] _RAND_2359;
  reg [31:0] _RAND_2360;
  reg [31:0] _RAND_2361;
  reg [31:0] _RAND_2362;
  reg [31:0] _RAND_2363;
  reg [31:0] _RAND_2364;
  reg [31:0] _RAND_2365;
  reg [31:0] _RAND_2366;
  reg [31:0] _RAND_2367;
  reg [31:0] _RAND_2368;
  reg [31:0] _RAND_2369;
  reg [31:0] _RAND_2370;
  reg [31:0] _RAND_2371;
  reg [31:0] _RAND_2372;
  reg [63:0] _RAND_2373;
  reg [31:0] _RAND_2374;
  reg [31:0] _RAND_2375;
  reg [31:0] _RAND_2376;
  reg [31:0] _RAND_2377;
  reg [31:0] _RAND_2378;
  reg [31:0] _RAND_2379;
  reg [31:0] _RAND_2380;
  reg [31:0] _RAND_2381;
  reg [31:0] _RAND_2382;
  reg [31:0] _RAND_2383;
  reg [31:0] _RAND_2384;
  reg [31:0] _RAND_2385;
  reg [31:0] _RAND_2386;
  reg [31:0] _RAND_2387;
  reg [31:0] _RAND_2388;
  reg [31:0] _RAND_2389;
  reg [31:0] _RAND_2390;
  reg [31:0] _RAND_2391;
  reg [31:0] _RAND_2392;
  reg [31:0] _RAND_2393;
  reg [31:0] _RAND_2394;
  reg [31:0] _RAND_2395;
  reg [31:0] _RAND_2396;
  reg [31:0] _RAND_2397;
  reg [31:0] _RAND_2398;
  reg [31:0] _RAND_2399;
  reg [31:0] _RAND_2400;
  reg [31:0] _RAND_2401;
  reg [31:0] _RAND_2402;
  reg [31:0] _RAND_2403;
  reg [31:0] _RAND_2404;
  reg [31:0] _RAND_2405;
  reg [31:0] _RAND_2406;
  reg [31:0] _RAND_2407;
  reg [31:0] _RAND_2408;
  reg [31:0] _RAND_2409;
  reg [31:0] _RAND_2410;
  reg [31:0] _RAND_2411;
  reg [31:0] _RAND_2412;
  reg [31:0] _RAND_2413;
  reg [31:0] _RAND_2414;
  reg [31:0] _RAND_2415;
  reg [31:0] _RAND_2416;
  reg [63:0] _RAND_2417;
  reg [31:0] _RAND_2418;
  reg [31:0] _RAND_2419;
  reg [31:0] _RAND_2420;
  reg [31:0] _RAND_2421;
  reg [31:0] _RAND_2422;
  reg [31:0] _RAND_2423;
  reg [31:0] _RAND_2424;
  reg [31:0] _RAND_2425;
  reg [31:0] _RAND_2426;
  reg [31:0] _RAND_2427;
  reg [31:0] _RAND_2428;
  reg [31:0] _RAND_2429;
  reg [31:0] _RAND_2430;
  reg [31:0] _RAND_2431;
  reg [31:0] _RAND_2432;
  reg [31:0] _RAND_2433;
  reg [31:0] _RAND_2434;
  reg [31:0] _RAND_2435;
  reg [31:0] _RAND_2436;
  reg [31:0] _RAND_2437;
  reg [31:0] _RAND_2438;
  reg [31:0] _RAND_2439;
  reg [31:0] _RAND_2440;
  reg [31:0] _RAND_2441;
  reg [31:0] _RAND_2442;
  reg [31:0] _RAND_2443;
  reg [31:0] _RAND_2444;
  reg [31:0] _RAND_2445;
  reg [31:0] _RAND_2446;
  reg [31:0] _RAND_2447;
  reg [31:0] _RAND_2448;
  reg [31:0] _RAND_2449;
  reg [31:0] _RAND_2450;
  reg [31:0] _RAND_2451;
  reg [31:0] _RAND_2452;
  reg [31:0] _RAND_2453;
  reg [31:0] _RAND_2454;
  reg [31:0] _RAND_2455;
  reg [31:0] _RAND_2456;
  reg [31:0] _RAND_2457;
  reg [31:0] _RAND_2458;
  reg [31:0] _RAND_2459;
  reg [31:0] _RAND_2460;
  reg [31:0] _RAND_2461;
  reg [31:0] _RAND_2462;
  reg [31:0] _RAND_2463;
  reg [31:0] _RAND_2464;
  reg [31:0] _RAND_2465;
  reg [31:0] _RAND_2466;
  reg [31:0] _RAND_2467;
  reg [31:0] _RAND_2468;
  reg [31:0] _RAND_2469;
  reg [63:0] _RAND_2470;
  reg [31:0] _RAND_2471;
  reg [31:0] _RAND_2472;
  reg [31:0] _RAND_2473;
  reg [31:0] _RAND_2474;
  reg [31:0] _RAND_2475;
  reg [31:0] _RAND_2476;
  reg [31:0] _RAND_2477;
  reg [31:0] _RAND_2478;
  reg [31:0] _RAND_2479;
  reg [31:0] _RAND_2480;
  reg [31:0] _RAND_2481;
  reg [31:0] _RAND_2482;
  reg [31:0] _RAND_2483;
  reg [31:0] _RAND_2484;
  reg [31:0] _RAND_2485;
  reg [31:0] _RAND_2486;
  reg [31:0] _RAND_2487;
  reg [31:0] _RAND_2488;
  reg [31:0] _RAND_2489;
  reg [31:0] _RAND_2490;
  reg [31:0] _RAND_2491;
  reg [31:0] _RAND_2492;
  reg [31:0] _RAND_2493;
  reg [31:0] _RAND_2494;
  reg [31:0] _RAND_2495;
  reg [31:0] _RAND_2496;
  reg [31:0] _RAND_2497;
  reg [31:0] _RAND_2498;
  reg [31:0] _RAND_2499;
  reg [31:0] _RAND_2500;
  reg [31:0] _RAND_2501;
  reg [31:0] _RAND_2502;
  reg [31:0] _RAND_2503;
  reg [31:0] _RAND_2504;
  reg [31:0] _RAND_2505;
  reg [31:0] _RAND_2506;
  reg [31:0] _RAND_2507;
  reg [31:0] _RAND_2508;
  reg [31:0] _RAND_2509;
  reg [31:0] _RAND_2510;
  reg [31:0] _RAND_2511;
  reg [31:0] _RAND_2512;
  reg [31:0] _RAND_2513;
  reg [63:0] _RAND_2514;
  reg [31:0] _RAND_2515;
  reg [31:0] _RAND_2516;
  reg [31:0] _RAND_2517;
  reg [31:0] _RAND_2518;
  reg [31:0] _RAND_2519;
  reg [31:0] _RAND_2520;
  reg [31:0] _RAND_2521;
  reg [31:0] _RAND_2522;
  reg [31:0] _RAND_2523;
  reg [31:0] _RAND_2524;
  reg [31:0] _RAND_2525;
  reg [31:0] _RAND_2526;
  reg [31:0] _RAND_2527;
  reg [31:0] _RAND_2528;
  reg [31:0] _RAND_2529;
  reg [31:0] _RAND_2530;
  reg [31:0] _RAND_2531;
  reg [31:0] _RAND_2532;
  reg [31:0] _RAND_2533;
  reg [31:0] _RAND_2534;
  reg [31:0] _RAND_2535;
  reg [31:0] _RAND_2536;
  reg [31:0] _RAND_2537;
  reg [31:0] _RAND_2538;
  reg [31:0] _RAND_2539;
  reg [31:0] _RAND_2540;
  reg [31:0] _RAND_2541;
  reg [31:0] _RAND_2542;
  reg [31:0] _RAND_2543;
  reg [31:0] _RAND_2544;
  reg [31:0] _RAND_2545;
  reg [31:0] _RAND_2546;
  reg [31:0] _RAND_2547;
  reg [31:0] _RAND_2548;
  reg [31:0] _RAND_2549;
  reg [31:0] _RAND_2550;
  reg [31:0] _RAND_2551;
  reg [31:0] _RAND_2552;
  reg [31:0] _RAND_2553;
  reg [31:0] _RAND_2554;
  reg [31:0] _RAND_2555;
  reg [31:0] _RAND_2556;
  reg [31:0] _RAND_2557;
  reg [31:0] _RAND_2558;
  reg [31:0] _RAND_2559;
  reg [31:0] _RAND_2560;
  reg [31:0] _RAND_2561;
  reg [31:0] _RAND_2562;
  reg [31:0] _RAND_2563;
  reg [31:0] _RAND_2564;
  reg [31:0] _RAND_2565;
  reg [31:0] _RAND_2566;
  reg [63:0] _RAND_2567;
  reg [31:0] _RAND_2568;
  reg [31:0] _RAND_2569;
  reg [31:0] _RAND_2570;
  reg [31:0] _RAND_2571;
  reg [31:0] _RAND_2572;
  reg [31:0] _RAND_2573;
  reg [31:0] _RAND_2574;
  reg [31:0] _RAND_2575;
  reg [31:0] _RAND_2576;
  reg [31:0] _RAND_2577;
  reg [31:0] _RAND_2578;
  reg [31:0] _RAND_2579;
  reg [31:0] _RAND_2580;
  reg [31:0] _RAND_2581;
  reg [31:0] _RAND_2582;
  reg [31:0] _RAND_2583;
  reg [31:0] _RAND_2584;
  reg [31:0] _RAND_2585;
  reg [31:0] _RAND_2586;
  reg [31:0] _RAND_2587;
  reg [31:0] _RAND_2588;
  reg [31:0] _RAND_2589;
  reg [31:0] _RAND_2590;
  reg [31:0] _RAND_2591;
  reg [31:0] _RAND_2592;
  reg [31:0] _RAND_2593;
  reg [31:0] _RAND_2594;
  reg [31:0] _RAND_2595;
  reg [31:0] _RAND_2596;
  reg [31:0] _RAND_2597;
  reg [31:0] _RAND_2598;
  reg [31:0] _RAND_2599;
  reg [31:0] _RAND_2600;
  reg [31:0] _RAND_2601;
  reg [31:0] _RAND_2602;
  reg [31:0] _RAND_2603;
  reg [31:0] _RAND_2604;
  reg [31:0] _RAND_2605;
  reg [31:0] _RAND_2606;
  reg [31:0] _RAND_2607;
  reg [31:0] _RAND_2608;
  reg [31:0] _RAND_2609;
  reg [31:0] _RAND_2610;
  reg [63:0] _RAND_2611;
  reg [31:0] _RAND_2612;
  reg [31:0] _RAND_2613;
  reg [31:0] _RAND_2614;
  reg [31:0] _RAND_2615;
  reg [31:0] _RAND_2616;
  reg [31:0] _RAND_2617;
  reg [31:0] _RAND_2618;
  reg [31:0] _RAND_2619;
  reg [31:0] _RAND_2620;
  reg [31:0] _RAND_2621;
  reg [31:0] _RAND_2622;
  reg [31:0] _RAND_2623;
  reg [31:0] _RAND_2624;
  reg [31:0] _RAND_2625;
  reg [31:0] _RAND_2626;
  reg [31:0] _RAND_2627;
  reg [31:0] _RAND_2628;
  reg [31:0] _RAND_2629;
  reg [31:0] _RAND_2630;
  reg [31:0] _RAND_2631;
  reg [31:0] _RAND_2632;
  reg [31:0] _RAND_2633;
  reg [31:0] _RAND_2634;
  reg [31:0] _RAND_2635;
  reg [31:0] _RAND_2636;
  reg [31:0] _RAND_2637;
  reg [31:0] _RAND_2638;
  reg [31:0] _RAND_2639;
  reg [31:0] _RAND_2640;
  reg [31:0] _RAND_2641;
  reg [31:0] _RAND_2642;
  reg [31:0] _RAND_2643;
  reg [31:0] _RAND_2644;
  reg [31:0] _RAND_2645;
  reg [31:0] _RAND_2646;
  reg [31:0] _RAND_2647;
  reg [31:0] _RAND_2648;
  reg [31:0] _RAND_2649;
  reg [31:0] _RAND_2650;
  reg [31:0] _RAND_2651;
  reg [31:0] _RAND_2652;
  reg [31:0] _RAND_2653;
  reg [31:0] _RAND_2654;
  reg [31:0] _RAND_2655;
  reg [31:0] _RAND_2656;
  reg [31:0] _RAND_2657;
  reg [31:0] _RAND_2658;
  reg [31:0] _RAND_2659;
  reg [31:0] _RAND_2660;
  reg [31:0] _RAND_2661;
  reg [31:0] _RAND_2662;
  reg [31:0] _RAND_2663;
  reg [63:0] _RAND_2664;
  reg [31:0] _RAND_2665;
  reg [31:0] _RAND_2666;
  reg [31:0] _RAND_2667;
  reg [31:0] _RAND_2668;
  reg [31:0] _RAND_2669;
  reg [31:0] _RAND_2670;
  reg [31:0] _RAND_2671;
  reg [31:0] _RAND_2672;
  reg [31:0] _RAND_2673;
  reg [31:0] _RAND_2674;
  reg [31:0] _RAND_2675;
  reg [31:0] _RAND_2676;
  reg [31:0] _RAND_2677;
  reg [31:0] _RAND_2678;
  reg [31:0] _RAND_2679;
  reg [31:0] _RAND_2680;
  reg [31:0] _RAND_2681;
  reg [31:0] _RAND_2682;
  reg [31:0] _RAND_2683;
  reg [31:0] _RAND_2684;
  reg [31:0] _RAND_2685;
  reg [31:0] _RAND_2686;
  reg [31:0] _RAND_2687;
  reg [31:0] _RAND_2688;
  reg [31:0] _RAND_2689;
  reg [31:0] _RAND_2690;
  reg [31:0] _RAND_2691;
  reg [31:0] _RAND_2692;
  reg [31:0] _RAND_2693;
  reg [31:0] _RAND_2694;
  reg [31:0] _RAND_2695;
  reg [31:0] _RAND_2696;
  reg [31:0] _RAND_2697;
  reg [31:0] _RAND_2698;
  reg [31:0] _RAND_2699;
  reg [31:0] _RAND_2700;
  reg [31:0] _RAND_2701;
  reg [31:0] _RAND_2702;
  reg [31:0] _RAND_2703;
  reg [31:0] _RAND_2704;
  reg [31:0] _RAND_2705;
  reg [31:0] _RAND_2706;
  reg [31:0] _RAND_2707;
  reg [63:0] _RAND_2708;
  reg [31:0] _RAND_2709;
  reg [31:0] _RAND_2710;
  reg [31:0] _RAND_2711;
  reg [31:0] _RAND_2712;
  reg [31:0] _RAND_2713;
  reg [31:0] _RAND_2714;
  reg [31:0] _RAND_2715;
  reg [31:0] _RAND_2716;
  reg [31:0] _RAND_2717;
  reg [31:0] _RAND_2718;
  reg [31:0] _RAND_2719;
  reg [31:0] _RAND_2720;
  reg [31:0] _RAND_2721;
  reg [31:0] _RAND_2722;
  reg [31:0] _RAND_2723;
  reg [31:0] _RAND_2724;
  reg [31:0] _RAND_2725;
  reg [31:0] _RAND_2726;
  reg [31:0] _RAND_2727;
  reg [31:0] _RAND_2728;
  reg [31:0] _RAND_2729;
  reg [31:0] _RAND_2730;
  reg [31:0] _RAND_2731;
  reg [31:0] _RAND_2732;
  reg [31:0] _RAND_2733;
  reg [31:0] _RAND_2734;
  reg [31:0] _RAND_2735;
  reg [31:0] _RAND_2736;
  reg [31:0] _RAND_2737;
  reg [31:0] _RAND_2738;
  reg [31:0] _RAND_2739;
  reg [31:0] _RAND_2740;
  reg [31:0] _RAND_2741;
  reg [31:0] _RAND_2742;
  reg [31:0] _RAND_2743;
  reg [31:0] _RAND_2744;
  reg [31:0] _RAND_2745;
  reg [31:0] _RAND_2746;
  reg [31:0] _RAND_2747;
  reg [31:0] _RAND_2748;
  reg [31:0] _RAND_2749;
  reg [31:0] _RAND_2750;
  reg [31:0] _RAND_2751;
  reg [31:0] _RAND_2752;
  reg [31:0] _RAND_2753;
  reg [31:0] _RAND_2754;
  reg [31:0] _RAND_2755;
  reg [31:0] _RAND_2756;
  reg [31:0] _RAND_2757;
  reg [31:0] _RAND_2758;
  reg [31:0] _RAND_2759;
  reg [31:0] _RAND_2760;
  reg [31:0] _RAND_2761;
  reg [31:0] _RAND_2762;
  reg [31:0] _RAND_2763;
  reg [31:0] _RAND_2764;
  reg [63:0] _RAND_2765;
  reg [31:0] _RAND_2766;
  reg [31:0] _RAND_2767;
  reg [31:0] _RAND_2768;
  reg [31:0] _RAND_2769;
  reg [31:0] _RAND_2770;
  reg [31:0] _RAND_2771;
  reg [31:0] _RAND_2772;
  reg [31:0] _RAND_2773;
  reg [31:0] _RAND_2774;
  reg [31:0] _RAND_2775;
  reg [31:0] _RAND_2776;
  reg [31:0] _RAND_2777;
  reg [31:0] _RAND_2778;
  reg [31:0] _RAND_2779;
  reg [31:0] _RAND_2780;
  reg [31:0] _RAND_2781;
  reg [31:0] _RAND_2782;
  reg [31:0] _RAND_2783;
  reg [31:0] _RAND_2784;
  reg [31:0] _RAND_2785;
  reg [31:0] _RAND_2786;
  reg [31:0] _RAND_2787;
  reg [31:0] _RAND_2788;
  reg [31:0] _RAND_2789;
  reg [31:0] _RAND_2790;
  reg [31:0] _RAND_2791;
  reg [31:0] _RAND_2792;
  reg [31:0] _RAND_2793;
  reg [31:0] _RAND_2794;
  reg [31:0] _RAND_2795;
  reg [31:0] _RAND_2796;
  reg [31:0] _RAND_2797;
  reg [31:0] _RAND_2798;
  reg [31:0] _RAND_2799;
  reg [31:0] _RAND_2800;
  reg [31:0] _RAND_2801;
  reg [31:0] _RAND_2802;
  reg [31:0] _RAND_2803;
  reg [31:0] _RAND_2804;
  reg [31:0] _RAND_2805;
  reg [31:0] _RAND_2806;
  reg [31:0] _RAND_2807;
  reg [31:0] _RAND_2808;
  reg [63:0] _RAND_2809;
  reg [31:0] _RAND_2810;
  reg [31:0] _RAND_2811;
  reg [31:0] _RAND_2812;
  reg [31:0] _RAND_2813;
  reg [31:0] _RAND_2814;
  reg [31:0] _RAND_2815;
  reg [31:0] _RAND_2816;
  reg [31:0] _RAND_2817;
  reg [31:0] _RAND_2818;
  reg [31:0] _RAND_2819;
  reg [31:0] _RAND_2820;
  reg [31:0] _RAND_2821;
  reg [31:0] _RAND_2822;
  reg [31:0] _RAND_2823;
  reg [31:0] _RAND_2824;
  reg [31:0] _RAND_2825;
  reg [31:0] _RAND_2826;
  reg [31:0] _RAND_2827;
  reg [31:0] _RAND_2828;
  reg [31:0] _RAND_2829;
  reg [31:0] _RAND_2830;
  reg [31:0] _RAND_2831;
  reg [31:0] _RAND_2832;
  reg [31:0] _RAND_2833;
  reg [31:0] _RAND_2834;
  reg [31:0] _RAND_2835;
  reg [31:0] _RAND_2836;
  reg [31:0] _RAND_2837;
  reg [31:0] _RAND_2838;
  reg [31:0] _RAND_2839;
  reg [31:0] _RAND_2840;
  reg [31:0] _RAND_2841;
  reg [31:0] _RAND_2842;
  reg [31:0] _RAND_2843;
  reg [31:0] _RAND_2844;
  reg [31:0] _RAND_2845;
  reg [31:0] _RAND_2846;
  reg [31:0] _RAND_2847;
  reg [31:0] _RAND_2848;
  reg [31:0] _RAND_2849;
  reg [31:0] _RAND_2850;
  reg [31:0] _RAND_2851;
  reg [31:0] _RAND_2852;
  reg [31:0] _RAND_2853;
  reg [31:0] _RAND_2854;
  reg [31:0] _RAND_2855;
  reg [31:0] _RAND_2856;
  reg [31:0] _RAND_2857;
  reg [31:0] _RAND_2858;
  reg [31:0] _RAND_2859;
  reg [31:0] _RAND_2860;
  reg [31:0] _RAND_2861;
  reg [63:0] _RAND_2862;
  reg [31:0] _RAND_2863;
  reg [31:0] _RAND_2864;
  reg [31:0] _RAND_2865;
  reg [31:0] _RAND_2866;
  reg [31:0] _RAND_2867;
  reg [31:0] _RAND_2868;
  reg [31:0] _RAND_2869;
  reg [31:0] _RAND_2870;
  reg [31:0] _RAND_2871;
  reg [31:0] _RAND_2872;
  reg [31:0] _RAND_2873;
  reg [31:0] _RAND_2874;
  reg [31:0] _RAND_2875;
  reg [31:0] _RAND_2876;
  reg [31:0] _RAND_2877;
  reg [31:0] _RAND_2878;
  reg [31:0] _RAND_2879;
  reg [31:0] _RAND_2880;
  reg [31:0] _RAND_2881;
  reg [31:0] _RAND_2882;
  reg [31:0] _RAND_2883;
  reg [31:0] _RAND_2884;
  reg [31:0] _RAND_2885;
  reg [31:0] _RAND_2886;
  reg [31:0] _RAND_2887;
  reg [31:0] _RAND_2888;
  reg [31:0] _RAND_2889;
  reg [31:0] _RAND_2890;
  reg [31:0] _RAND_2891;
  reg [31:0] _RAND_2892;
  reg [31:0] _RAND_2893;
  reg [31:0] _RAND_2894;
  reg [31:0] _RAND_2895;
  reg [31:0] _RAND_2896;
  reg [31:0] _RAND_2897;
  reg [31:0] _RAND_2898;
  reg [31:0] _RAND_2899;
  reg [31:0] _RAND_2900;
  reg [31:0] _RAND_2901;
  reg [31:0] _RAND_2902;
  reg [31:0] _RAND_2903;
  reg [31:0] _RAND_2904;
  reg [31:0] _RAND_2905;
  reg [63:0] _RAND_2906;
  reg [31:0] _RAND_2907;
  reg [31:0] _RAND_2908;
  reg [31:0] _RAND_2909;
  reg [31:0] _RAND_2910;
  reg [31:0] _RAND_2911;
  reg [31:0] _RAND_2912;
  reg [31:0] _RAND_2913;
  reg [31:0] _RAND_2914;
  reg [31:0] _RAND_2915;
  reg [31:0] _RAND_2916;
  reg [31:0] _RAND_2917;
  reg [31:0] _RAND_2918;
  reg [31:0] _RAND_2919;
  reg [31:0] _RAND_2920;
  reg [31:0] _RAND_2921;
  reg [31:0] _RAND_2922;
  reg [31:0] _RAND_2923;
  reg [31:0] _RAND_2924;
  reg [31:0] _RAND_2925;
  reg [31:0] _RAND_2926;
  reg [31:0] _RAND_2927;
  reg [31:0] _RAND_2928;
  reg [31:0] _RAND_2929;
  reg [31:0] _RAND_2930;
  reg [31:0] _RAND_2931;
  reg [31:0] _RAND_2932;
  reg [31:0] _RAND_2933;
  reg [31:0] _RAND_2934;
  reg [31:0] _RAND_2935;
  reg [31:0] _RAND_2936;
  reg [31:0] _RAND_2937;
  reg [31:0] _RAND_2938;
  reg [31:0] _RAND_2939;
  reg [31:0] _RAND_2940;
  reg [31:0] _RAND_2941;
  reg [31:0] _RAND_2942;
  reg [31:0] _RAND_2943;
  reg [31:0] _RAND_2944;
  reg [31:0] _RAND_2945;
  reg [31:0] _RAND_2946;
  reg [31:0] _RAND_2947;
  reg [31:0] _RAND_2948;
  reg [31:0] _RAND_2949;
  reg [31:0] _RAND_2950;
  reg [31:0] _RAND_2951;
  reg [31:0] _RAND_2952;
  reg [31:0] _RAND_2953;
  reg [31:0] _RAND_2954;
  reg [31:0] _RAND_2955;
  reg [31:0] _RAND_2956;
  reg [31:0] _RAND_2957;
  reg [31:0] _RAND_2958;
  reg [63:0] _RAND_2959;
  reg [31:0] _RAND_2960;
  reg [31:0] _RAND_2961;
  reg [31:0] _RAND_2962;
  reg [31:0] _RAND_2963;
  reg [31:0] _RAND_2964;
  reg [31:0] _RAND_2965;
  reg [31:0] _RAND_2966;
  reg [31:0] _RAND_2967;
  reg [31:0] _RAND_2968;
  reg [31:0] _RAND_2969;
  reg [31:0] _RAND_2970;
  reg [31:0] _RAND_2971;
  reg [31:0] _RAND_2972;
  reg [31:0] _RAND_2973;
  reg [31:0] _RAND_2974;
  reg [31:0] _RAND_2975;
  reg [31:0] _RAND_2976;
  reg [31:0] _RAND_2977;
  reg [31:0] _RAND_2978;
  reg [31:0] _RAND_2979;
  reg [31:0] _RAND_2980;
  reg [31:0] _RAND_2981;
  reg [31:0] _RAND_2982;
  reg [31:0] _RAND_2983;
  reg [31:0] _RAND_2984;
  reg [31:0] _RAND_2985;
  reg [31:0] _RAND_2986;
  reg [31:0] _RAND_2987;
  reg [31:0] _RAND_2988;
  reg [31:0] _RAND_2989;
  reg [31:0] _RAND_2990;
  reg [31:0] _RAND_2991;
  reg [31:0] _RAND_2992;
  reg [31:0] _RAND_2993;
  reg [31:0] _RAND_2994;
  reg [31:0] _RAND_2995;
  reg [31:0] _RAND_2996;
  reg [31:0] _RAND_2997;
  reg [31:0] _RAND_2998;
  reg [31:0] _RAND_2999;
  reg [31:0] _RAND_3000;
  reg [31:0] _RAND_3001;
  reg [31:0] _RAND_3002;
  reg [63:0] _RAND_3003;
  reg [31:0] _RAND_3004;
  reg [31:0] _RAND_3005;
  reg [31:0] _RAND_3006;
  reg [31:0] _RAND_3007;
  reg [31:0] _RAND_3008;
  reg [31:0] _RAND_3009;
  reg [31:0] _RAND_3010;
  reg [31:0] _RAND_3011;
  reg [31:0] _RAND_3012;
  reg [31:0] _RAND_3013;
  reg [31:0] _RAND_3014;
  reg [31:0] _RAND_3015;
  reg [31:0] _RAND_3016;
  reg [31:0] _RAND_3017;
  reg [31:0] _RAND_3018;
  reg [31:0] _RAND_3019;
  reg [31:0] _RAND_3020;
  reg [31:0] _RAND_3021;
  reg [31:0] _RAND_3022;
  reg [31:0] _RAND_3023;
  reg [31:0] _RAND_3024;
  reg [31:0] _RAND_3025;
  reg [31:0] _RAND_3026;
  reg [31:0] _RAND_3027;
  reg [31:0] _RAND_3028;
  reg [31:0] _RAND_3029;
  reg [31:0] _RAND_3030;
  reg [31:0] _RAND_3031;
  reg [31:0] _RAND_3032;
  reg [31:0] _RAND_3033;
  reg [31:0] _RAND_3034;
  reg [31:0] _RAND_3035;
  reg [31:0] _RAND_3036;
  reg [31:0] _RAND_3037;
  reg [31:0] _RAND_3038;
  reg [31:0] _RAND_3039;
  reg [31:0] _RAND_3040;
  reg [31:0] _RAND_3041;
  reg [31:0] _RAND_3042;
  reg [31:0] _RAND_3043;
  reg [31:0] _RAND_3044;
  reg [31:0] _RAND_3045;
  reg [31:0] _RAND_3046;
  reg [31:0] _RAND_3047;
  reg [31:0] _RAND_3048;
  reg [31:0] _RAND_3049;
  reg [31:0] _RAND_3050;
  reg [31:0] _RAND_3051;
  reg [31:0] _RAND_3052;
  reg [31:0] _RAND_3053;
  reg [31:0] _RAND_3054;
  reg [31:0] _RAND_3055;
  reg [63:0] _RAND_3056;
  reg [31:0] _RAND_3057;
  reg [31:0] _RAND_3058;
  reg [31:0] _RAND_3059;
  reg [31:0] _RAND_3060;
  reg [31:0] _RAND_3061;
  reg [31:0] _RAND_3062;
  reg [31:0] _RAND_3063;
  reg [31:0] _RAND_3064;
  reg [31:0] _RAND_3065;
  reg [31:0] _RAND_3066;
  reg [31:0] _RAND_3067;
  reg [31:0] _RAND_3068;
  reg [31:0] _RAND_3069;
  reg [31:0] _RAND_3070;
  reg [31:0] _RAND_3071;
  reg [31:0] _RAND_3072;
  reg [31:0] _RAND_3073;
  reg [31:0] _RAND_3074;
  reg [31:0] _RAND_3075;
  reg [31:0] _RAND_3076;
  reg [31:0] _RAND_3077;
  reg [31:0] _RAND_3078;
  reg [31:0] _RAND_3079;
  reg [31:0] _RAND_3080;
  reg [31:0] _RAND_3081;
  reg [31:0] _RAND_3082;
  reg [31:0] _RAND_3083;
  reg [31:0] _RAND_3084;
  reg [31:0] _RAND_3085;
  reg [31:0] _RAND_3086;
  reg [31:0] _RAND_3087;
  reg [31:0] _RAND_3088;
  reg [31:0] _RAND_3089;
  reg [31:0] _RAND_3090;
  reg [31:0] _RAND_3091;
  reg [31:0] _RAND_3092;
  reg [31:0] _RAND_3093;
  reg [31:0] _RAND_3094;
  reg [31:0] _RAND_3095;
  reg [31:0] _RAND_3096;
  reg [31:0] _RAND_3097;
  reg [31:0] _RAND_3098;
  reg [31:0] _RAND_3099;
  reg [63:0] _RAND_3100;
  reg [31:0] _RAND_3101;
  reg [31:0] _RAND_3102;
  reg [31:0] _RAND_3103;
  reg [31:0] _RAND_3104;
  reg [31:0] _RAND_3105;
  reg [31:0] _RAND_3106;
  reg [31:0] _RAND_3107;
  reg [31:0] _RAND_3108;
  reg [31:0] _RAND_3109;
  reg [31:0] _RAND_3110;
  reg [31:0] _RAND_3111;
  reg [31:0] _RAND_3112;
  reg [31:0] _RAND_3113;
  reg [31:0] _RAND_3114;
  reg [31:0] _RAND_3115;
  reg [31:0] _RAND_3116;
  reg [31:0] _RAND_3117;
  reg [31:0] _RAND_3118;
  reg [31:0] _RAND_3119;
  reg [31:0] _RAND_3120;
  reg [31:0] _RAND_3121;
  reg [31:0] _RAND_3122;
  reg [31:0] _RAND_3123;
  reg [31:0] _RAND_3124;
  reg [31:0] _RAND_3125;
  reg [31:0] _RAND_3126;
  reg [31:0] _RAND_3127;
  reg [31:0] _RAND_3128;
  reg [31:0] _RAND_3129;
  reg [31:0] _RAND_3130;
  reg [31:0] _RAND_3131;
  reg [31:0] _RAND_3132;
  reg [31:0] _RAND_3133;
  reg [31:0] _RAND_3134;
  reg [31:0] _RAND_3135;
  reg [31:0] _RAND_3136;
  reg [31:0] _RAND_3137;
  reg [31:0] _RAND_3138;
  reg [31:0] _RAND_3139;
`endif // RANDOMIZE_REG_INIT
  wire  trans_buffer_clock; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_reset; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_ready; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_valid; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_switch; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_switch_off; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_is_unicore; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_enq_bits_dec_uops_0_shift; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_0_lrs3_rtype; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_rflag; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_wflag; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_0_prflag; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_0_pwflag; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_pflag_busy; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_0_stale_pflag; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_0_op1_sel; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_0_op2_sel; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_0_split_num; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_0_self_index; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_0_rob_inst_idx; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_0_address_num; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_0_uopc; // @[enq_transBuff.scala 37:31]
  wire [31:0] trans_buffer_io_enq_bits_dec_uops_0_inst; // @[enq_transBuff.scala 37:31]
  wire [31:0] trans_buffer_io_enq_bits_dec_uops_0_debug_inst; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_is_rvc; // @[enq_transBuff.scala 37:31]
  wire [39:0] trans_buffer_io_enq_bits_dec_uops_0_debug_pc; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_enq_bits_dec_uops_0_iq_type; // @[enq_transBuff.scala 37:31]
  wire [9:0] trans_buffer_io_enq_bits_dec_uops_0_fu_code; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_0_ctrl_br_type; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_0_ctrl_op1_sel; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_enq_bits_dec_uops_0_ctrl_op2_sel; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_enq_bits_dec_uops_0_ctrl_imm_sel; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_0_ctrl_op_fcn; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_ctrl_fcn_dw; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_enq_bits_dec_uops_0_ctrl_csr_cmd; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_ctrl_is_load; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_ctrl_is_sta; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_ctrl_is_std; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_0_ctrl_op3_sel; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_0_iw_state; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_iw_p1_poisoned; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_iw_p2_poisoned; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_is_br; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_is_jalr; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_is_jal; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_is_sfb; // @[enq_transBuff.scala 37:31]
  wire [11:0] trans_buffer_io_enq_bits_dec_uops_0_br_mask; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_0_br_tag; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_enq_bits_dec_uops_0_ftq_idx; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_edge_inst; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_0_pc_lob; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_taken; // @[enq_transBuff.scala 37:31]
  wire [19:0] trans_buffer_io_enq_bits_dec_uops_0_imm_packed; // @[enq_transBuff.scala 37:31]
  wire [11:0] trans_buffer_io_enq_bits_dec_uops_0_csr_addr; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_0_rob_idx; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_enq_bits_dec_uops_0_ldq_idx; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_enq_bits_dec_uops_0_stq_idx; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_0_rxq_idx; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_0_pdst; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_0_prs1; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_0_prs2; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_0_prs3; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_enq_bits_dec_uops_0_ppred; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_prs1_busy; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_prs2_busy; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_prs3_busy; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_ppred_busy; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_0_stale_pdst; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_exception; // @[enq_transBuff.scala 37:31]
  wire [63:0] trans_buffer_io_enq_bits_dec_uops_0_exc_cause; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_bypassable; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_enq_bits_dec_uops_0_mem_cmd; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_0_mem_size; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_mem_signed; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_is_fence; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_is_fencei; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_is_amo; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_uses_ldq; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_uses_stq; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_is_sys_pc2epc; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_is_unique; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_flush_on_commit; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_ldst_is_rs1; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_0_ldst; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_0_lrs1; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_0_lrs2; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_0_lrs3; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_ldst_val; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_0_dst_rtype; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_0_lrs1_rtype; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_0_lrs2_rtype; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_frs3_en; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_fp_val; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_fp_single; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_xcpt_pf_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_xcpt_ae_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_xcpt_ma_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_bp_debug_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_0_bp_xcpt_if; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_0_debug_fsrc; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_0_debug_tsrc; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_switch; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_switch_off; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_is_unicore; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_enq_bits_dec_uops_1_shift; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_1_lrs3_rtype; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_rflag; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_wflag; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_1_prflag; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_1_pwflag; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_pflag_busy; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_1_stale_pflag; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_1_op1_sel; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_1_op2_sel; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_1_split_num; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_1_self_index; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_1_rob_inst_idx; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_1_address_num; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_1_uopc; // @[enq_transBuff.scala 37:31]
  wire [31:0] trans_buffer_io_enq_bits_dec_uops_1_inst; // @[enq_transBuff.scala 37:31]
  wire [31:0] trans_buffer_io_enq_bits_dec_uops_1_debug_inst; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_is_rvc; // @[enq_transBuff.scala 37:31]
  wire [39:0] trans_buffer_io_enq_bits_dec_uops_1_debug_pc; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_enq_bits_dec_uops_1_iq_type; // @[enq_transBuff.scala 37:31]
  wire [9:0] trans_buffer_io_enq_bits_dec_uops_1_fu_code; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_1_ctrl_br_type; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_1_ctrl_op1_sel; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_enq_bits_dec_uops_1_ctrl_op2_sel; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_enq_bits_dec_uops_1_ctrl_imm_sel; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_1_ctrl_op_fcn; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_ctrl_fcn_dw; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_enq_bits_dec_uops_1_ctrl_csr_cmd; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_ctrl_is_load; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_ctrl_is_sta; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_ctrl_is_std; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_1_ctrl_op3_sel; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_1_iw_state; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_iw_p1_poisoned; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_iw_p2_poisoned; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_is_br; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_is_jalr; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_is_jal; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_is_sfb; // @[enq_transBuff.scala 37:31]
  wire [11:0] trans_buffer_io_enq_bits_dec_uops_1_br_mask; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_1_br_tag; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_enq_bits_dec_uops_1_ftq_idx; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_edge_inst; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_1_pc_lob; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_taken; // @[enq_transBuff.scala 37:31]
  wire [19:0] trans_buffer_io_enq_bits_dec_uops_1_imm_packed; // @[enq_transBuff.scala 37:31]
  wire [11:0] trans_buffer_io_enq_bits_dec_uops_1_csr_addr; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_1_rob_idx; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_enq_bits_dec_uops_1_ldq_idx; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_enq_bits_dec_uops_1_stq_idx; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_1_rxq_idx; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_1_pdst; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_1_prs1; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_1_prs2; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_1_prs3; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_enq_bits_dec_uops_1_ppred; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_prs1_busy; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_prs2_busy; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_prs3_busy; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_ppred_busy; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_1_stale_pdst; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_exception; // @[enq_transBuff.scala 37:31]
  wire [63:0] trans_buffer_io_enq_bits_dec_uops_1_exc_cause; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_bypassable; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_enq_bits_dec_uops_1_mem_cmd; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_1_mem_size; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_mem_signed; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_is_fence; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_is_fencei; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_is_amo; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_uses_ldq; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_uses_stq; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_is_sys_pc2epc; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_is_unique; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_flush_on_commit; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_ldst_is_rs1; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_1_ldst; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_1_lrs1; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_1_lrs2; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_1_lrs3; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_ldst_val; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_1_dst_rtype; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_1_lrs1_rtype; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_1_lrs2_rtype; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_frs3_en; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_fp_val; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_fp_single; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_xcpt_pf_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_xcpt_ae_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_xcpt_ma_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_bp_debug_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_1_bp_xcpt_if; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_1_debug_fsrc; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_1_debug_tsrc; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_switch; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_switch_off; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_is_unicore; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_enq_bits_dec_uops_2_shift; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_2_lrs3_rtype; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_rflag; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_wflag; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_2_prflag; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_2_pwflag; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_pflag_busy; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_2_stale_pflag; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_2_op1_sel; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_2_op2_sel; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_2_split_num; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_2_self_index; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_2_rob_inst_idx; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_2_address_num; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_2_uopc; // @[enq_transBuff.scala 37:31]
  wire [31:0] trans_buffer_io_enq_bits_dec_uops_2_inst; // @[enq_transBuff.scala 37:31]
  wire [31:0] trans_buffer_io_enq_bits_dec_uops_2_debug_inst; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_is_rvc; // @[enq_transBuff.scala 37:31]
  wire [39:0] trans_buffer_io_enq_bits_dec_uops_2_debug_pc; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_enq_bits_dec_uops_2_iq_type; // @[enq_transBuff.scala 37:31]
  wire [9:0] trans_buffer_io_enq_bits_dec_uops_2_fu_code; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_2_ctrl_br_type; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_2_ctrl_op1_sel; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_enq_bits_dec_uops_2_ctrl_op2_sel; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_enq_bits_dec_uops_2_ctrl_imm_sel; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_2_ctrl_op_fcn; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_ctrl_fcn_dw; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_enq_bits_dec_uops_2_ctrl_csr_cmd; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_ctrl_is_load; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_ctrl_is_sta; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_ctrl_is_std; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_2_ctrl_op3_sel; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_2_iw_state; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_iw_p1_poisoned; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_iw_p2_poisoned; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_is_br; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_is_jalr; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_is_jal; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_is_sfb; // @[enq_transBuff.scala 37:31]
  wire [11:0] trans_buffer_io_enq_bits_dec_uops_2_br_mask; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_2_br_tag; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_enq_bits_dec_uops_2_ftq_idx; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_edge_inst; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_2_pc_lob; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_taken; // @[enq_transBuff.scala 37:31]
  wire [19:0] trans_buffer_io_enq_bits_dec_uops_2_imm_packed; // @[enq_transBuff.scala 37:31]
  wire [11:0] trans_buffer_io_enq_bits_dec_uops_2_csr_addr; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_2_rob_idx; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_enq_bits_dec_uops_2_ldq_idx; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_enq_bits_dec_uops_2_stq_idx; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_2_rxq_idx; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_2_pdst; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_2_prs1; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_2_prs2; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_2_prs3; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_enq_bits_dec_uops_2_ppred; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_prs1_busy; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_prs2_busy; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_prs3_busy; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_ppred_busy; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_2_stale_pdst; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_exception; // @[enq_transBuff.scala 37:31]
  wire [63:0] trans_buffer_io_enq_bits_dec_uops_2_exc_cause; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_bypassable; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_enq_bits_dec_uops_2_mem_cmd; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_2_mem_size; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_mem_signed; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_is_fence; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_is_fencei; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_is_amo; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_uses_ldq; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_uses_stq; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_is_sys_pc2epc; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_is_unique; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_flush_on_commit; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_ldst_is_rs1; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_2_ldst; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_2_lrs1; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_2_lrs2; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_2_lrs3; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_ldst_val; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_2_dst_rtype; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_2_lrs1_rtype; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_2_lrs2_rtype; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_frs3_en; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_fp_val; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_fp_single; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_xcpt_pf_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_xcpt_ae_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_xcpt_ma_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_bp_debug_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_2_bp_xcpt_if; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_2_debug_fsrc; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_2_debug_tsrc; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_switch; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_switch_off; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_is_unicore; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_enq_bits_dec_uops_3_shift; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_3_lrs3_rtype; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_rflag; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_wflag; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_3_prflag; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_3_pwflag; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_pflag_busy; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_3_stale_pflag; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_3_op1_sel; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_3_op2_sel; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_3_split_num; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_3_self_index; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_3_rob_inst_idx; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_3_address_num; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_3_uopc; // @[enq_transBuff.scala 37:31]
  wire [31:0] trans_buffer_io_enq_bits_dec_uops_3_inst; // @[enq_transBuff.scala 37:31]
  wire [31:0] trans_buffer_io_enq_bits_dec_uops_3_debug_inst; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_is_rvc; // @[enq_transBuff.scala 37:31]
  wire [39:0] trans_buffer_io_enq_bits_dec_uops_3_debug_pc; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_enq_bits_dec_uops_3_iq_type; // @[enq_transBuff.scala 37:31]
  wire [9:0] trans_buffer_io_enq_bits_dec_uops_3_fu_code; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_3_ctrl_br_type; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_3_ctrl_op1_sel; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_enq_bits_dec_uops_3_ctrl_op2_sel; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_enq_bits_dec_uops_3_ctrl_imm_sel; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_3_ctrl_op_fcn; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_ctrl_fcn_dw; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_enq_bits_dec_uops_3_ctrl_csr_cmd; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_ctrl_is_load; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_ctrl_is_sta; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_ctrl_is_std; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_3_ctrl_op3_sel; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_3_iw_state; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_iw_p1_poisoned; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_iw_p2_poisoned; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_is_br; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_is_jalr; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_is_jal; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_is_sfb; // @[enq_transBuff.scala 37:31]
  wire [11:0] trans_buffer_io_enq_bits_dec_uops_3_br_mask; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_enq_bits_dec_uops_3_br_tag; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_enq_bits_dec_uops_3_ftq_idx; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_edge_inst; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_3_pc_lob; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_taken; // @[enq_transBuff.scala 37:31]
  wire [19:0] trans_buffer_io_enq_bits_dec_uops_3_imm_packed; // @[enq_transBuff.scala 37:31]
  wire [11:0] trans_buffer_io_enq_bits_dec_uops_3_csr_addr; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_3_rob_idx; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_enq_bits_dec_uops_3_ldq_idx; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_enq_bits_dec_uops_3_stq_idx; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_3_rxq_idx; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_3_pdst; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_3_prs1; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_3_prs2; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_3_prs3; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_enq_bits_dec_uops_3_ppred; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_prs1_busy; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_prs2_busy; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_prs3_busy; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_ppred_busy; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_enq_bits_dec_uops_3_stale_pdst; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_exception; // @[enq_transBuff.scala 37:31]
  wire [63:0] trans_buffer_io_enq_bits_dec_uops_3_exc_cause; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_bypassable; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_enq_bits_dec_uops_3_mem_cmd; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_3_mem_size; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_mem_signed; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_is_fence; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_is_fencei; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_is_amo; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_uses_ldq; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_uses_stq; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_is_sys_pc2epc; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_is_unique; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_flush_on_commit; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_ldst_is_rs1; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_3_ldst; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_3_lrs1; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_3_lrs2; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_enq_bits_dec_uops_3_lrs3; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_ldst_val; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_3_dst_rtype; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_3_lrs1_rtype; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_3_lrs2_rtype; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_frs3_en; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_fp_val; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_fp_single; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_xcpt_pf_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_xcpt_ae_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_xcpt_ma_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_bp_debug_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_dec_uops_3_bp_xcpt_if; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_3_debug_fsrc; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_enq_bits_dec_uops_3_debug_tsrc; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_val_mask_0; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_val_mask_1; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_val_mask_2; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_enq_bits_val_mask_3; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_ready; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_valid; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_switch; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_switch_off; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_is_unicore; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_deq_bits_tran_uops_0_shift; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_0_lrs3_rtype; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_rflag; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_wflag; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_deq_bits_tran_uops_0_prflag; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_deq_bits_tran_uops_0_pwflag; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_pflag_busy; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_deq_bits_tran_uops_0_stale_pflag; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_deq_bits_tran_uops_0_op1_sel; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_deq_bits_tran_uops_0_op2_sel; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_deq_bits_tran_uops_0_split_num; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_deq_bits_tran_uops_0_self_index; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_deq_bits_tran_uops_0_rob_inst_idx; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_deq_bits_tran_uops_0_address_num; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_deq_bits_tran_uops_0_uopc; // @[enq_transBuff.scala 37:31]
  wire [31:0] trans_buffer_io_deq_bits_tran_uops_0_inst; // @[enq_transBuff.scala 37:31]
  wire [31:0] trans_buffer_io_deq_bits_tran_uops_0_debug_inst; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_is_rvc; // @[enq_transBuff.scala 37:31]
  wire [39:0] trans_buffer_io_deq_bits_tran_uops_0_debug_pc; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_deq_bits_tran_uops_0_iq_type; // @[enq_transBuff.scala 37:31]
  wire [9:0] trans_buffer_io_deq_bits_tran_uops_0_fu_code; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_deq_bits_tran_uops_0_ctrl_br_type; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_0_ctrl_op1_sel; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_deq_bits_tran_uops_0_ctrl_op2_sel; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_deq_bits_tran_uops_0_ctrl_imm_sel; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_deq_bits_tran_uops_0_ctrl_op_fcn; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_ctrl_fcn_dw; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_deq_bits_tran_uops_0_ctrl_csr_cmd; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_ctrl_is_load; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_ctrl_is_sta; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_ctrl_is_std; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_0_ctrl_op3_sel; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_0_iw_state; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_iw_p1_poisoned; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_iw_p2_poisoned; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_is_br; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_is_jalr; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_is_jal; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_is_sfb; // @[enq_transBuff.scala 37:31]
  wire [11:0] trans_buffer_io_deq_bits_tran_uops_0_br_mask; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_deq_bits_tran_uops_0_br_tag; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_deq_bits_tran_uops_0_ftq_idx; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_edge_inst; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_deq_bits_tran_uops_0_pc_lob; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_taken; // @[enq_transBuff.scala 37:31]
  wire [19:0] trans_buffer_io_deq_bits_tran_uops_0_imm_packed; // @[enq_transBuff.scala 37:31]
  wire [11:0] trans_buffer_io_deq_bits_tran_uops_0_csr_addr; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_deq_bits_tran_uops_0_rob_idx; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_deq_bits_tran_uops_0_ldq_idx; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_deq_bits_tran_uops_0_stq_idx; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_0_rxq_idx; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_deq_bits_tran_uops_0_pdst; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_deq_bits_tran_uops_0_prs1; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_deq_bits_tran_uops_0_prs2; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_deq_bits_tran_uops_0_prs3; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_deq_bits_tran_uops_0_ppred; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_prs1_busy; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_prs2_busy; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_prs3_busy; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_ppred_busy; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_deq_bits_tran_uops_0_stale_pdst; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_exception; // @[enq_transBuff.scala 37:31]
  wire [63:0] trans_buffer_io_deq_bits_tran_uops_0_exc_cause; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_bypassable; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_deq_bits_tran_uops_0_mem_cmd; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_0_mem_size; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_mem_signed; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_is_fence; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_is_fencei; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_is_amo; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_uses_ldq; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_uses_stq; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_is_sys_pc2epc; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_is_unique; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_flush_on_commit; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_ldst_is_rs1; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_deq_bits_tran_uops_0_ldst; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_deq_bits_tran_uops_0_lrs1; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_deq_bits_tran_uops_0_lrs2; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_deq_bits_tran_uops_0_lrs3; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_ldst_val; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_0_dst_rtype; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_0_lrs1_rtype; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_0_lrs2_rtype; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_frs3_en; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_fp_val; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_fp_single; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_xcpt_pf_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_xcpt_ae_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_xcpt_ma_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_bp_debug_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_0_bp_xcpt_if; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_0_debug_fsrc; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_0_debug_tsrc; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_switch; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_switch_off; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_is_unicore; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_deq_bits_tran_uops_1_shift; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_1_lrs3_rtype; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_rflag; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_wflag; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_deq_bits_tran_uops_1_prflag; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_deq_bits_tran_uops_1_pwflag; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_pflag_busy; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_deq_bits_tran_uops_1_stale_pflag; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_deq_bits_tran_uops_1_op1_sel; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_deq_bits_tran_uops_1_op2_sel; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_deq_bits_tran_uops_1_split_num; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_deq_bits_tran_uops_1_self_index; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_deq_bits_tran_uops_1_rob_inst_idx; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_deq_bits_tran_uops_1_address_num; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_deq_bits_tran_uops_1_uopc; // @[enq_transBuff.scala 37:31]
  wire [31:0] trans_buffer_io_deq_bits_tran_uops_1_inst; // @[enq_transBuff.scala 37:31]
  wire [31:0] trans_buffer_io_deq_bits_tran_uops_1_debug_inst; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_is_rvc; // @[enq_transBuff.scala 37:31]
  wire [39:0] trans_buffer_io_deq_bits_tran_uops_1_debug_pc; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_deq_bits_tran_uops_1_iq_type; // @[enq_transBuff.scala 37:31]
  wire [9:0] trans_buffer_io_deq_bits_tran_uops_1_fu_code; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_deq_bits_tran_uops_1_ctrl_br_type; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_1_ctrl_op1_sel; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_deq_bits_tran_uops_1_ctrl_op2_sel; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_deq_bits_tran_uops_1_ctrl_imm_sel; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_deq_bits_tran_uops_1_ctrl_op_fcn; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_ctrl_fcn_dw; // @[enq_transBuff.scala 37:31]
  wire [2:0] trans_buffer_io_deq_bits_tran_uops_1_ctrl_csr_cmd; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_ctrl_is_load; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_ctrl_is_sta; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_ctrl_is_std; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_1_ctrl_op3_sel; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_1_iw_state; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_iw_p1_poisoned; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_iw_p2_poisoned; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_is_br; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_is_jalr; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_is_jal; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_is_sfb; // @[enq_transBuff.scala 37:31]
  wire [11:0] trans_buffer_io_deq_bits_tran_uops_1_br_mask; // @[enq_transBuff.scala 37:31]
  wire [3:0] trans_buffer_io_deq_bits_tran_uops_1_br_tag; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_deq_bits_tran_uops_1_ftq_idx; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_edge_inst; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_deq_bits_tran_uops_1_pc_lob; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_taken; // @[enq_transBuff.scala 37:31]
  wire [19:0] trans_buffer_io_deq_bits_tran_uops_1_imm_packed; // @[enq_transBuff.scala 37:31]
  wire [11:0] trans_buffer_io_deq_bits_tran_uops_1_csr_addr; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_deq_bits_tran_uops_1_rob_idx; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_deq_bits_tran_uops_1_ldq_idx; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_deq_bits_tran_uops_1_stq_idx; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_1_rxq_idx; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_deq_bits_tran_uops_1_pdst; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_deq_bits_tran_uops_1_prs1; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_deq_bits_tran_uops_1_prs2; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_deq_bits_tran_uops_1_prs3; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_deq_bits_tran_uops_1_ppred; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_prs1_busy; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_prs2_busy; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_prs3_busy; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_ppred_busy; // @[enq_transBuff.scala 37:31]
  wire [6:0] trans_buffer_io_deq_bits_tran_uops_1_stale_pdst; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_exception; // @[enq_transBuff.scala 37:31]
  wire [63:0] trans_buffer_io_deq_bits_tran_uops_1_exc_cause; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_bypassable; // @[enq_transBuff.scala 37:31]
  wire [4:0] trans_buffer_io_deq_bits_tran_uops_1_mem_cmd; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_1_mem_size; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_mem_signed; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_is_fence; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_is_fencei; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_is_amo; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_uses_ldq; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_uses_stq; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_is_sys_pc2epc; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_is_unique; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_flush_on_commit; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_ldst_is_rs1; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_deq_bits_tran_uops_1_ldst; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_deq_bits_tran_uops_1_lrs1; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_deq_bits_tran_uops_1_lrs2; // @[enq_transBuff.scala 37:31]
  wire [5:0] trans_buffer_io_deq_bits_tran_uops_1_lrs3; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_ldst_val; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_1_dst_rtype; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_1_lrs1_rtype; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_1_lrs2_rtype; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_frs3_en; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_fp_val; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_fp_single; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_xcpt_pf_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_xcpt_ae_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_xcpt_ma_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_bp_debug_if; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_uops_1_bp_xcpt_if; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_1_debug_fsrc; // @[enq_transBuff.scala 37:31]
  wire [1:0] trans_buffer_io_deq_bits_tran_uops_1_debug_tsrc; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_valids_0; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_deq_bits_tran_valids_1; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_clear; // @[enq_transBuff.scala 37:31]
  wire  trans_buffer_io_isUnicoreMode; // @[enq_transBuff.scala 37:31]
  reg  enq_buffer_0_dec_uops_0_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_0_dec_uops_0_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_0_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_0_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_0_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_0_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_0_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_0_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_0_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_0_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_0_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_0_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_0_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_0_dec_uops_0_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_0_dec_uops_0_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_0_dec_uops_0_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_0_dec_uops_0_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_0_dec_uops_0_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_0_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_0_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_0_dec_uops_0_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_0_dec_uops_0_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_0_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_0_dec_uops_0_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_0_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_0_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_0_dec_uops_0_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_0_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_0_dec_uops_0_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_0_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_0_dec_uops_0_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_0_dec_uops_0_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_0_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_0_dec_uops_0_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_0_dec_uops_0_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_0_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_0_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_0_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_0_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_0_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_0_dec_uops_0_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_0_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_0_dec_uops_0_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_0_dec_uops_0_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_0_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_0_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_0_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_0_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_0_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_0_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_0_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_0_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_0_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_0_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_0_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_0_dec_uops_1_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_1_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_1_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_1_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_1_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_1_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_1_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_1_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_1_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_1_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_1_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_1_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_0_dec_uops_1_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_0_dec_uops_1_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_0_dec_uops_1_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_0_dec_uops_1_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_0_dec_uops_1_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_1_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_1_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_0_dec_uops_1_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_0_dec_uops_1_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_1_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_0_dec_uops_1_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_1_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_1_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_0_dec_uops_1_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_1_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_0_dec_uops_1_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_1_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_0_dec_uops_1_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_0_dec_uops_1_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_1_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_0_dec_uops_1_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_0_dec_uops_1_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_1_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_1_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_1_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_1_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_1_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_0_dec_uops_1_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_1_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_0_dec_uops_1_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_0_dec_uops_1_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_1_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_1_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_1_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_1_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_1_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_1_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_1_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_1_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_1_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_1_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_1_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_0_dec_uops_2_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_2_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_2_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_2_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_2_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_2_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_2_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_2_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_2_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_2_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_2_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_2_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_0_dec_uops_2_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_0_dec_uops_2_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_0_dec_uops_2_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_0_dec_uops_2_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_0_dec_uops_2_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_2_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_2_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_0_dec_uops_2_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_0_dec_uops_2_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_2_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_0_dec_uops_2_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_2_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_2_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_0_dec_uops_2_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_2_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_0_dec_uops_2_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_2_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_0_dec_uops_2_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_0_dec_uops_2_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_2_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_0_dec_uops_2_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_0_dec_uops_2_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_2_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_2_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_2_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_2_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_2_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_0_dec_uops_2_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_2_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_0_dec_uops_2_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_0_dec_uops_2_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_2_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_2_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_2_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_2_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_2_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_2_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_2_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_2_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_2_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_2_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_2_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_0_dec_uops_3_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_3_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_3_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_3_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_3_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_3_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_3_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_3_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_3_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_3_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_3_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_3_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_0_dec_uops_3_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_0_dec_uops_3_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_0_dec_uops_3_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_0_dec_uops_3_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_0_dec_uops_3_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_3_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_3_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_0_dec_uops_3_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_0_dec_uops_3_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_3_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_0_dec_uops_3_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_3_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_3_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_0_dec_uops_3_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_0_dec_uops_3_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_0_dec_uops_3_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_3_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_0_dec_uops_3_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_0_dec_uops_3_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_3_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_0_dec_uops_3_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_0_dec_uops_3_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_3_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_3_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_3_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_3_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_3_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_0_dec_uops_3_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_0_dec_uops_3_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_0_dec_uops_3_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_0_dec_uops_3_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_3_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_3_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_3_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_3_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_0_dec_uops_3_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_3_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_3_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_3_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_dec_uops_3_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_3_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_0_dec_uops_3_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_val_mask_0; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_val_mask_1; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_val_mask_2; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_0_val_mask_3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_1_dec_uops_0_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_0_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_0_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_0_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_0_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_0_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_0_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_0_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_0_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_0_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_0_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_0_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_1_dec_uops_0_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_1_dec_uops_0_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_1_dec_uops_0_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_1_dec_uops_0_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_1_dec_uops_0_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_0_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_0_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_1_dec_uops_0_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_1_dec_uops_0_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_0_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_1_dec_uops_0_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_0_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_0_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_1_dec_uops_0_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_0_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_1_dec_uops_0_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_0_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_1_dec_uops_0_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_1_dec_uops_0_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_0_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_1_dec_uops_0_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_1_dec_uops_0_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_0_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_0_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_0_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_0_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_0_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_1_dec_uops_0_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_0_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_1_dec_uops_0_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_1_dec_uops_0_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_0_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_0_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_0_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_0_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_0_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_0_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_0_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_0_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_0_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_0_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_0_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_1_dec_uops_1_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_1_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_1_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_1_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_1_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_1_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_1_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_1_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_1_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_1_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_1_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_1_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_1_dec_uops_1_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_1_dec_uops_1_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_1_dec_uops_1_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_1_dec_uops_1_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_1_dec_uops_1_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_1_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_1_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_1_dec_uops_1_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_1_dec_uops_1_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_1_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_1_dec_uops_1_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_1_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_1_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_1_dec_uops_1_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_1_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_1_dec_uops_1_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_1_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_1_dec_uops_1_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_1_dec_uops_1_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_1_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_1_dec_uops_1_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_1_dec_uops_1_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_1_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_1_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_1_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_1_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_1_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_1_dec_uops_1_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_1_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_1_dec_uops_1_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_1_dec_uops_1_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_1_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_1_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_1_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_1_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_1_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_1_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_1_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_1_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_1_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_1_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_1_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_1_dec_uops_2_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_2_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_2_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_2_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_2_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_2_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_2_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_2_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_2_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_2_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_2_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_2_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_1_dec_uops_2_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_1_dec_uops_2_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_1_dec_uops_2_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_1_dec_uops_2_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_1_dec_uops_2_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_2_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_2_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_1_dec_uops_2_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_1_dec_uops_2_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_2_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_1_dec_uops_2_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_2_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_2_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_1_dec_uops_2_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_2_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_1_dec_uops_2_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_2_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_1_dec_uops_2_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_1_dec_uops_2_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_2_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_1_dec_uops_2_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_1_dec_uops_2_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_2_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_2_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_2_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_2_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_2_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_1_dec_uops_2_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_2_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_1_dec_uops_2_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_1_dec_uops_2_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_2_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_2_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_2_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_2_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_2_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_2_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_2_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_2_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_2_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_2_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_2_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_1_dec_uops_3_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_3_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_3_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_3_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_3_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_3_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_3_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_3_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_3_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_3_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_3_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_3_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_1_dec_uops_3_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_1_dec_uops_3_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_1_dec_uops_3_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_1_dec_uops_3_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_1_dec_uops_3_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_3_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_3_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_1_dec_uops_3_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_1_dec_uops_3_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_3_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_1_dec_uops_3_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_3_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_3_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_1_dec_uops_3_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_1_dec_uops_3_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_1_dec_uops_3_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_3_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_1_dec_uops_3_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_1_dec_uops_3_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_3_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_1_dec_uops_3_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_1_dec_uops_3_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_3_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_3_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_3_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_3_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_3_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_1_dec_uops_3_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_1_dec_uops_3_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_1_dec_uops_3_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_1_dec_uops_3_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_3_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_3_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_3_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_3_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_1_dec_uops_3_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_3_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_3_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_3_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_dec_uops_3_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_3_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_1_dec_uops_3_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_val_mask_0; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_val_mask_1; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_val_mask_2; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_1_val_mask_3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_2_dec_uops_0_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_0_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_0_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_0_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_0_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_0_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_0_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_0_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_0_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_0_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_0_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_0_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_2_dec_uops_0_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_2_dec_uops_0_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_2_dec_uops_0_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_2_dec_uops_0_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_2_dec_uops_0_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_0_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_0_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_2_dec_uops_0_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_2_dec_uops_0_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_0_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_2_dec_uops_0_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_0_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_0_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_2_dec_uops_0_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_0_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_2_dec_uops_0_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_0_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_2_dec_uops_0_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_2_dec_uops_0_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_0_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_2_dec_uops_0_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_2_dec_uops_0_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_0_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_0_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_0_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_0_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_0_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_2_dec_uops_0_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_0_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_2_dec_uops_0_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_2_dec_uops_0_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_0_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_0_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_0_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_0_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_0_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_0_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_0_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_0_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_0_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_0_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_0_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_2_dec_uops_1_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_1_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_1_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_1_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_1_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_1_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_1_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_1_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_1_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_1_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_1_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_1_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_2_dec_uops_1_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_2_dec_uops_1_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_2_dec_uops_1_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_2_dec_uops_1_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_2_dec_uops_1_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_1_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_1_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_2_dec_uops_1_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_2_dec_uops_1_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_1_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_2_dec_uops_1_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_1_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_1_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_2_dec_uops_1_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_1_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_2_dec_uops_1_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_1_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_2_dec_uops_1_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_2_dec_uops_1_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_1_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_2_dec_uops_1_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_2_dec_uops_1_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_1_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_1_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_1_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_1_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_1_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_2_dec_uops_1_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_1_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_2_dec_uops_1_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_2_dec_uops_1_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_1_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_1_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_1_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_1_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_1_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_1_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_1_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_1_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_1_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_1_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_1_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_2_dec_uops_2_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_2_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_2_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_2_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_2_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_2_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_2_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_2_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_2_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_2_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_2_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_2_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_2_dec_uops_2_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_2_dec_uops_2_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_2_dec_uops_2_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_2_dec_uops_2_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_2_dec_uops_2_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_2_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_2_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_2_dec_uops_2_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_2_dec_uops_2_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_2_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_2_dec_uops_2_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_2_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_2_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_2_dec_uops_2_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_2_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_2_dec_uops_2_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_2_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_2_dec_uops_2_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_2_dec_uops_2_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_2_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_2_dec_uops_2_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_2_dec_uops_2_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_2_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_2_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_2_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_2_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_2_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_2_dec_uops_2_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_2_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_2_dec_uops_2_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_2_dec_uops_2_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_2_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_2_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_2_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_2_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_2_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_2_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_2_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_2_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_2_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_2_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_2_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_2_dec_uops_3_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_3_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_3_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_3_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_3_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_3_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_3_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_3_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_3_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_3_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_3_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_3_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_2_dec_uops_3_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_2_dec_uops_3_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_2_dec_uops_3_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_2_dec_uops_3_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_2_dec_uops_3_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_3_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_3_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_2_dec_uops_3_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_2_dec_uops_3_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_3_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_2_dec_uops_3_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_3_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_3_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_2_dec_uops_3_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_2_dec_uops_3_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_2_dec_uops_3_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_3_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_2_dec_uops_3_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_2_dec_uops_3_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_3_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_2_dec_uops_3_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_2_dec_uops_3_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_3_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_3_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_3_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_3_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_3_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_2_dec_uops_3_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_2_dec_uops_3_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_2_dec_uops_3_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_2_dec_uops_3_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_3_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_3_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_3_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_3_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_2_dec_uops_3_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_3_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_3_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_3_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_dec_uops_3_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_3_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_2_dec_uops_3_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_val_mask_0; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_val_mask_1; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_val_mask_2; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_2_val_mask_3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_3_dec_uops_0_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_0_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_0_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_0_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_0_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_0_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_0_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_0_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_0_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_0_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_0_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_0_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_3_dec_uops_0_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_3_dec_uops_0_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_3_dec_uops_0_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_3_dec_uops_0_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_3_dec_uops_0_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_0_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_0_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_3_dec_uops_0_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_3_dec_uops_0_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_0_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_3_dec_uops_0_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_0_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_0_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_3_dec_uops_0_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_0_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_3_dec_uops_0_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_0_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_3_dec_uops_0_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_3_dec_uops_0_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_0_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_3_dec_uops_0_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_3_dec_uops_0_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_0_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_0_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_0_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_0_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_0_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_3_dec_uops_0_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_0_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_3_dec_uops_0_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_3_dec_uops_0_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_0_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_0_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_0_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_0_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_0_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_0_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_0_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_0_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_0_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_0_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_0_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_3_dec_uops_1_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_1_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_1_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_1_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_1_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_1_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_1_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_1_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_1_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_1_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_1_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_1_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_3_dec_uops_1_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_3_dec_uops_1_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_3_dec_uops_1_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_3_dec_uops_1_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_3_dec_uops_1_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_1_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_1_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_3_dec_uops_1_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_3_dec_uops_1_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_1_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_3_dec_uops_1_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_1_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_1_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_3_dec_uops_1_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_1_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_3_dec_uops_1_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_1_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_3_dec_uops_1_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_3_dec_uops_1_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_1_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_3_dec_uops_1_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_3_dec_uops_1_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_1_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_1_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_1_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_1_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_1_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_3_dec_uops_1_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_1_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_3_dec_uops_1_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_3_dec_uops_1_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_1_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_1_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_1_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_1_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_1_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_1_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_1_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_1_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_1_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_1_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_1_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_3_dec_uops_2_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_2_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_2_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_2_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_2_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_2_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_2_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_2_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_2_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_2_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_2_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_2_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_3_dec_uops_2_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_3_dec_uops_2_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_3_dec_uops_2_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_3_dec_uops_2_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_3_dec_uops_2_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_2_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_2_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_3_dec_uops_2_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_3_dec_uops_2_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_2_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_3_dec_uops_2_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_2_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_2_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_3_dec_uops_2_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_2_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_3_dec_uops_2_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_2_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_3_dec_uops_2_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_3_dec_uops_2_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_2_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_3_dec_uops_2_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_3_dec_uops_2_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_2_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_2_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_2_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_2_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_2_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_3_dec_uops_2_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_2_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_3_dec_uops_2_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_3_dec_uops_2_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_2_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_2_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_2_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_2_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_2_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_2_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_2_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_2_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_2_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_2_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_2_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_3_dec_uops_3_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_3_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_3_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_3_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_3_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_3_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_3_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_3_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_3_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_3_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_3_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_3_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_3_dec_uops_3_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_3_dec_uops_3_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_3_dec_uops_3_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_3_dec_uops_3_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_3_dec_uops_3_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_3_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_3_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_3_dec_uops_3_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_3_dec_uops_3_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_3_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_3_dec_uops_3_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_3_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_3_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_3_dec_uops_3_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_3_dec_uops_3_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_3_dec_uops_3_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_3_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_3_dec_uops_3_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_3_dec_uops_3_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_3_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_3_dec_uops_3_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_3_dec_uops_3_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_3_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_3_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_3_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_3_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_3_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_3_dec_uops_3_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_3_dec_uops_3_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_3_dec_uops_3_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_3_dec_uops_3_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_3_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_3_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_3_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_3_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_3_dec_uops_3_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_3_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_3_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_3_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_dec_uops_3_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_3_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_3_dec_uops_3_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_val_mask_0; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_val_mask_1; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_val_mask_2; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_3_val_mask_3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_4_dec_uops_0_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_0_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_0_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_0_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_0_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_0_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_0_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_0_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_0_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_0_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_0_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_0_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_4_dec_uops_0_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_4_dec_uops_0_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_4_dec_uops_0_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_4_dec_uops_0_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_4_dec_uops_0_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_0_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_0_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_4_dec_uops_0_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_4_dec_uops_0_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_0_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_4_dec_uops_0_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_0_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_0_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_4_dec_uops_0_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_0_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_4_dec_uops_0_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_0_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_4_dec_uops_0_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_4_dec_uops_0_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_0_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_4_dec_uops_0_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_4_dec_uops_0_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_0_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_0_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_0_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_0_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_0_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_4_dec_uops_0_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_0_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_4_dec_uops_0_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_4_dec_uops_0_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_0_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_0_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_0_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_0_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_0_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_0_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_0_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_0_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_0_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_0_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_0_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_4_dec_uops_1_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_1_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_1_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_1_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_1_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_1_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_1_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_1_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_1_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_1_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_1_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_1_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_4_dec_uops_1_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_4_dec_uops_1_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_4_dec_uops_1_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_4_dec_uops_1_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_4_dec_uops_1_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_1_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_1_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_4_dec_uops_1_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_4_dec_uops_1_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_1_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_4_dec_uops_1_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_1_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_1_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_4_dec_uops_1_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_1_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_4_dec_uops_1_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_1_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_4_dec_uops_1_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_4_dec_uops_1_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_1_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_4_dec_uops_1_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_4_dec_uops_1_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_1_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_1_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_1_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_1_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_1_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_4_dec_uops_1_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_1_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_4_dec_uops_1_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_4_dec_uops_1_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_1_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_1_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_1_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_1_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_1_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_1_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_1_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_1_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_1_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_1_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_1_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_4_dec_uops_2_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_2_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_2_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_2_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_2_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_2_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_2_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_2_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_2_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_2_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_2_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_2_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_4_dec_uops_2_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_4_dec_uops_2_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_4_dec_uops_2_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_4_dec_uops_2_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_4_dec_uops_2_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_2_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_2_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_4_dec_uops_2_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_4_dec_uops_2_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_2_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_4_dec_uops_2_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_2_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_2_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_4_dec_uops_2_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_2_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_4_dec_uops_2_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_2_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_4_dec_uops_2_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_4_dec_uops_2_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_2_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_4_dec_uops_2_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_4_dec_uops_2_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_2_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_2_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_2_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_2_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_2_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_4_dec_uops_2_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_2_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_4_dec_uops_2_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_4_dec_uops_2_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_2_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_2_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_2_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_2_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_2_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_2_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_2_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_2_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_2_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_2_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_2_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_4_dec_uops_3_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_3_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_3_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_3_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_3_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_3_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_3_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_3_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_3_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_3_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_3_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_3_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_4_dec_uops_3_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_4_dec_uops_3_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_4_dec_uops_3_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_4_dec_uops_3_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_4_dec_uops_3_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_3_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_3_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_4_dec_uops_3_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_4_dec_uops_3_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_3_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_4_dec_uops_3_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_3_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_3_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_4_dec_uops_3_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_4_dec_uops_3_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_4_dec_uops_3_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_3_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_4_dec_uops_3_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_4_dec_uops_3_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_3_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_4_dec_uops_3_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_4_dec_uops_3_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_3_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_3_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_3_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_3_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_3_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_4_dec_uops_3_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_4_dec_uops_3_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_4_dec_uops_3_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_4_dec_uops_3_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_3_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_3_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_3_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_3_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_4_dec_uops_3_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_3_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_3_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_3_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_dec_uops_3_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_3_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_4_dec_uops_3_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_val_mask_0; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_val_mask_1; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_val_mask_2; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_4_val_mask_3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_5_dec_uops_0_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_0_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_0_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_0_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_0_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_0_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_0_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_0_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_0_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_0_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_0_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_0_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_5_dec_uops_0_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_5_dec_uops_0_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_5_dec_uops_0_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_5_dec_uops_0_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_5_dec_uops_0_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_0_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_0_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_5_dec_uops_0_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_5_dec_uops_0_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_0_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_5_dec_uops_0_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_0_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_0_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_5_dec_uops_0_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_0_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_5_dec_uops_0_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_0_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_5_dec_uops_0_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_5_dec_uops_0_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_0_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_5_dec_uops_0_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_5_dec_uops_0_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_0_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_0_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_0_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_0_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_0_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_5_dec_uops_0_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_0_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_5_dec_uops_0_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_5_dec_uops_0_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_0_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_0_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_0_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_0_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_0_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_0_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_0_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_0_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_0_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_0_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_0_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_5_dec_uops_1_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_1_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_1_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_1_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_1_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_1_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_1_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_1_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_1_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_1_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_1_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_1_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_5_dec_uops_1_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_5_dec_uops_1_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_5_dec_uops_1_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_5_dec_uops_1_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_5_dec_uops_1_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_1_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_1_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_5_dec_uops_1_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_5_dec_uops_1_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_1_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_5_dec_uops_1_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_1_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_1_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_5_dec_uops_1_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_1_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_5_dec_uops_1_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_1_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_5_dec_uops_1_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_5_dec_uops_1_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_1_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_5_dec_uops_1_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_5_dec_uops_1_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_1_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_1_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_1_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_1_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_1_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_5_dec_uops_1_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_1_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_5_dec_uops_1_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_5_dec_uops_1_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_1_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_1_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_1_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_1_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_1_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_1_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_1_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_1_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_1_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_1_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_1_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_5_dec_uops_2_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_2_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_2_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_2_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_2_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_2_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_2_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_2_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_2_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_2_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_2_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_2_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_5_dec_uops_2_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_5_dec_uops_2_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_5_dec_uops_2_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_5_dec_uops_2_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_5_dec_uops_2_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_2_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_2_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_5_dec_uops_2_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_5_dec_uops_2_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_2_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_5_dec_uops_2_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_2_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_2_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_5_dec_uops_2_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_2_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_5_dec_uops_2_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_2_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_5_dec_uops_2_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_5_dec_uops_2_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_2_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_5_dec_uops_2_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_5_dec_uops_2_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_2_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_2_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_2_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_2_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_2_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_5_dec_uops_2_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_2_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_5_dec_uops_2_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_5_dec_uops_2_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_2_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_2_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_2_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_2_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_2_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_2_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_2_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_2_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_2_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_2_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_2_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_5_dec_uops_3_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_3_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_3_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_3_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_3_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_3_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_3_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_3_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_3_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_3_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_3_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_3_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_5_dec_uops_3_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_5_dec_uops_3_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_5_dec_uops_3_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_5_dec_uops_3_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_5_dec_uops_3_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_3_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_3_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_5_dec_uops_3_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_5_dec_uops_3_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_3_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_5_dec_uops_3_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_3_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_3_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_5_dec_uops_3_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_5_dec_uops_3_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_5_dec_uops_3_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_3_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_5_dec_uops_3_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_5_dec_uops_3_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_3_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_5_dec_uops_3_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_5_dec_uops_3_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_3_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_3_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_3_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_3_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_3_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_5_dec_uops_3_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_5_dec_uops_3_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_5_dec_uops_3_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_5_dec_uops_3_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_3_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_3_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_3_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_3_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_5_dec_uops_3_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_3_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_3_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_3_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_dec_uops_3_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_3_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_5_dec_uops_3_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_val_mask_0; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_val_mask_1; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_val_mask_2; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_5_val_mask_3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_6_dec_uops_0_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_0_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_0_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_0_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_0_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_0_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_0_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_0_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_0_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_0_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_0_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_0_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_6_dec_uops_0_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_6_dec_uops_0_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_6_dec_uops_0_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_6_dec_uops_0_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_6_dec_uops_0_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_0_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_0_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_6_dec_uops_0_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_6_dec_uops_0_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_0_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_6_dec_uops_0_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_0_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_0_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_6_dec_uops_0_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_0_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_6_dec_uops_0_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_0_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_6_dec_uops_0_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_6_dec_uops_0_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_0_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_6_dec_uops_0_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_6_dec_uops_0_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_0_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_0_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_0_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_0_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_0_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_6_dec_uops_0_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_0_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_6_dec_uops_0_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_6_dec_uops_0_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_0_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_0_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_0_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_0_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_0_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_0_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_0_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_0_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_0_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_0_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_0_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_6_dec_uops_1_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_1_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_1_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_1_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_1_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_1_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_1_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_1_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_1_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_1_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_1_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_1_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_6_dec_uops_1_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_6_dec_uops_1_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_6_dec_uops_1_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_6_dec_uops_1_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_6_dec_uops_1_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_1_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_1_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_6_dec_uops_1_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_6_dec_uops_1_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_1_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_6_dec_uops_1_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_1_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_1_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_6_dec_uops_1_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_1_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_6_dec_uops_1_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_1_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_6_dec_uops_1_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_6_dec_uops_1_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_1_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_6_dec_uops_1_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_6_dec_uops_1_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_1_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_1_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_1_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_1_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_1_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_6_dec_uops_1_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_1_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_6_dec_uops_1_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_6_dec_uops_1_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_1_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_1_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_1_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_1_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_1_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_1_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_1_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_1_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_1_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_1_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_1_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_6_dec_uops_2_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_2_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_2_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_2_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_2_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_2_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_2_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_2_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_2_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_2_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_2_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_2_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_6_dec_uops_2_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_6_dec_uops_2_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_6_dec_uops_2_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_6_dec_uops_2_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_6_dec_uops_2_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_2_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_2_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_6_dec_uops_2_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_6_dec_uops_2_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_2_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_6_dec_uops_2_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_2_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_2_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_6_dec_uops_2_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_2_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_6_dec_uops_2_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_2_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_6_dec_uops_2_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_6_dec_uops_2_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_2_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_6_dec_uops_2_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_6_dec_uops_2_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_2_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_2_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_2_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_2_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_2_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_6_dec_uops_2_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_2_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_6_dec_uops_2_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_6_dec_uops_2_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_2_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_2_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_2_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_2_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_2_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_2_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_2_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_2_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_2_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_2_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_2_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_6_dec_uops_3_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_3_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_3_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_3_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_3_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_3_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_3_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_3_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_3_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_3_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_3_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_3_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_6_dec_uops_3_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_6_dec_uops_3_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_6_dec_uops_3_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_6_dec_uops_3_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_6_dec_uops_3_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_3_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_3_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_6_dec_uops_3_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_6_dec_uops_3_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_3_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_6_dec_uops_3_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_3_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_3_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_6_dec_uops_3_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_6_dec_uops_3_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_6_dec_uops_3_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_3_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_6_dec_uops_3_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_6_dec_uops_3_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_3_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_6_dec_uops_3_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_6_dec_uops_3_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_3_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_3_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_3_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_3_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_3_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_6_dec_uops_3_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_6_dec_uops_3_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_6_dec_uops_3_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_6_dec_uops_3_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_3_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_3_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_3_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_3_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_6_dec_uops_3_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_3_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_3_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_3_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_dec_uops_3_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_3_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_6_dec_uops_3_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_val_mask_0; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_val_mask_1; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_val_mask_2; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_6_val_mask_3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_7_dec_uops_0_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_0_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_0_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_0_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_0_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_0_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_0_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_0_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_0_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_0_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_0_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_0_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_7_dec_uops_0_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_7_dec_uops_0_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_7_dec_uops_0_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_7_dec_uops_0_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_7_dec_uops_0_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_0_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_0_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_7_dec_uops_0_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_7_dec_uops_0_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_0_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_7_dec_uops_0_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_0_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_0_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_7_dec_uops_0_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_0_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_7_dec_uops_0_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_0_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_7_dec_uops_0_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_7_dec_uops_0_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_0_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_7_dec_uops_0_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_7_dec_uops_0_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_0_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_0_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_0_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_0_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_0_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_7_dec_uops_0_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_0_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_7_dec_uops_0_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_7_dec_uops_0_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_0_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_0_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_0_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_0_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_0_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_0_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_0_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_0_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_0_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_0_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_0_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_7_dec_uops_1_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_1_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_1_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_1_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_1_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_1_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_1_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_1_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_1_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_1_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_1_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_1_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_7_dec_uops_1_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_7_dec_uops_1_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_7_dec_uops_1_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_7_dec_uops_1_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_7_dec_uops_1_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_1_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_1_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_7_dec_uops_1_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_7_dec_uops_1_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_1_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_7_dec_uops_1_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_1_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_1_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_7_dec_uops_1_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_1_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_7_dec_uops_1_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_1_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_7_dec_uops_1_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_7_dec_uops_1_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_1_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_7_dec_uops_1_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_7_dec_uops_1_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_1_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_1_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_1_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_1_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_1_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_7_dec_uops_1_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_1_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_7_dec_uops_1_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_7_dec_uops_1_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_1_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_1_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_1_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_1_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_1_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_1_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_1_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_1_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_1_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_1_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_1_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_7_dec_uops_2_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_2_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_2_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_2_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_2_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_2_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_2_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_2_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_2_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_2_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_2_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_2_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_7_dec_uops_2_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_7_dec_uops_2_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_7_dec_uops_2_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_7_dec_uops_2_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_7_dec_uops_2_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_2_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_2_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_7_dec_uops_2_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_7_dec_uops_2_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_2_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_7_dec_uops_2_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_2_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_2_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_7_dec_uops_2_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_2_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_7_dec_uops_2_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_2_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_7_dec_uops_2_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_7_dec_uops_2_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_2_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_7_dec_uops_2_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_7_dec_uops_2_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_2_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_2_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_2_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_2_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_2_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_7_dec_uops_2_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_2_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_7_dec_uops_2_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_7_dec_uops_2_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_2_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_2_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_2_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_2_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_2_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_2_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_2_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_2_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_2_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_2_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_2_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_switch; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_switch_off; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_is_unicore; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_7_dec_uops_3_shift; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_3_lrs3_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_rflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_wflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_3_prflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_3_pwflag; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_pflag_busy; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_3_stale_pflag; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_3_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_3_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_3_split_num; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_3_self_index; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_3_rob_inst_idx; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_3_address_num; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_3_uopc; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_7_dec_uops_3_inst; // @[enq_transBuff.scala 50:25]
  reg [31:0] enq_buffer_7_dec_uops_3_debug_inst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_is_rvc; // @[enq_transBuff.scala 50:25]
  reg [39:0] enq_buffer_7_dec_uops_3_debug_pc; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_7_dec_uops_3_iq_type; // @[enq_transBuff.scala 50:25]
  reg [9:0] enq_buffer_7_dec_uops_3_fu_code; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_3_ctrl_br_type; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_3_ctrl_op1_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_7_dec_uops_3_ctrl_op2_sel; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_7_dec_uops_3_ctrl_imm_sel; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_3_ctrl_op_fcn; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_ctrl_fcn_dw; // @[enq_transBuff.scala 50:25]
  reg [2:0] enq_buffer_7_dec_uops_3_ctrl_csr_cmd; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_ctrl_is_load; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_ctrl_is_sta; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_ctrl_is_std; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_3_ctrl_op3_sel; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_3_iw_state; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_iw_p1_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_iw_p2_poisoned; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_is_br; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_is_jalr; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_is_jal; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_is_sfb; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_7_dec_uops_3_br_mask; // @[enq_transBuff.scala 50:25]
  reg [3:0] enq_buffer_7_dec_uops_3_br_tag; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_7_dec_uops_3_ftq_idx; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_edge_inst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_3_pc_lob; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_taken; // @[enq_transBuff.scala 50:25]
  reg [19:0] enq_buffer_7_dec_uops_3_imm_packed; // @[enq_transBuff.scala 50:25]
  reg [11:0] enq_buffer_7_dec_uops_3_csr_addr; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_3_rob_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_7_dec_uops_3_ldq_idx; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_7_dec_uops_3_stq_idx; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_3_rxq_idx; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_3_pdst; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_3_prs1; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_3_prs2; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_3_prs3; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_7_dec_uops_3_ppred; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_prs1_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_prs2_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_prs3_busy; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_ppred_busy; // @[enq_transBuff.scala 50:25]
  reg [6:0] enq_buffer_7_dec_uops_3_stale_pdst; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_exception; // @[enq_transBuff.scala 50:25]
  reg [63:0] enq_buffer_7_dec_uops_3_exc_cause; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_bypassable; // @[enq_transBuff.scala 50:25]
  reg [4:0] enq_buffer_7_dec_uops_3_mem_cmd; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_3_mem_size; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_mem_signed; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_is_fence; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_is_fencei; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_is_amo; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_uses_ldq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_uses_stq; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_is_sys_pc2epc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_is_unique; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_flush_on_commit; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_ldst_is_rs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_3_ldst; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_3_lrs1; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_3_lrs2; // @[enq_transBuff.scala 50:25]
  reg [5:0] enq_buffer_7_dec_uops_3_lrs3; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_ldst_val; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_3_dst_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_3_lrs1_rtype; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_3_lrs2_rtype; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_frs3_en; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_fp_val; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_fp_single; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_xcpt_pf_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_xcpt_ae_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_xcpt_ma_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_bp_debug_if; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_dec_uops_3_bp_xcpt_if; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_3_debug_fsrc; // @[enq_transBuff.scala 50:25]
  reg [1:0] enq_buffer_7_dec_uops_3_debug_tsrc; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_val_mask_0; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_val_mask_1; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_val_mask_2; // @[enq_transBuff.scala 50:25]
  reg  enq_buffer_7_val_mask_3; // @[enq_transBuff.scala 50:25]
  reg  enq_valid; // @[enq_transBuff.scala 51:24]
  reg [4:0] set_idx; // @[enq_transBuff.scala 53:26]
  reg [4:0] set_num; // @[enq_transBuff.scala 54:26]
  wire  _T = set_idx == 5'h0; // @[enq_transBuff.scala 61:44]
  wire  _T_2 = io_enq_valid & set_idx == 5'h0 & trans_buffer_io_enq_ready; // @[enq_transBuff.scala 61:52]
  wire  _T_3 = io_set_num == 5'h0; // @[enq_transBuff.scala 61:94]
  wire  _T_6 = set_idx == set_num; // @[enq_transBuff.scala 61:145]
  wire  isBound = io_enq_valid & set_idx == 5'h0 & trans_buffer_io_enq_ready ? io_set_num == 5'h0 & set_idx == 5'h0 :
    enq_valid & set_idx == set_num & trans_buffer_io_enq_ready; // @[enq_transBuff.scala 61:19]
  wire  _T_16 = enq_valid ? _T_6 & trans_buffer_io_enq_ready : 1'h1; // @[enq_transBuff.scala 79:28]
  wire  last_cycle_over = _T_2 ? _T_3 : _T_16; // @[enq_transBuff.scala 78:27]
  reg  REG; // @[enq_transBuff.scala 81:41]
  wire [4:0] _T_24 = set_idx + 5'h1; // @[enq_transBuff.scala 112:39]
  wire [4:0] _GEN_1 = isBound ? 5'h0 : _T_24; // @[enq_transBuff.scala 107:22 enq_transBuff.scala 108:21 enq_transBuff.scala 112:21]
  wire  _GEN_3144 = 3'h1 == set_idx[2:0] ? enq_buffer_1_val_mask_0 : enq_buffer_0_val_mask_0; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3145 = 3'h2 == set_idx[2:0] ? enq_buffer_2_val_mask_0 : _GEN_3144; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3146 = 3'h3 == set_idx[2:0] ? enq_buffer_3_val_mask_0 : _GEN_3145; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3147 = 3'h4 == set_idx[2:0] ? enq_buffer_4_val_mask_0 : _GEN_3146; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3148 = 3'h5 == set_idx[2:0] ? enq_buffer_5_val_mask_0 : _GEN_3147; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3149 = 3'h6 == set_idx[2:0] ? enq_buffer_6_val_mask_0 : _GEN_3148; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3150 = 3'h7 == set_idx[2:0] ? enq_buffer_7_val_mask_0 : _GEN_3149; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3152 = 3'h1 == set_idx[2:0] ? enq_buffer_1_val_mask_1 : enq_buffer_0_val_mask_1; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3153 = 3'h2 == set_idx[2:0] ? enq_buffer_2_val_mask_1 : _GEN_3152; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3154 = 3'h3 == set_idx[2:0] ? enq_buffer_3_val_mask_1 : _GEN_3153; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3155 = 3'h4 == set_idx[2:0] ? enq_buffer_4_val_mask_1 : _GEN_3154; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3156 = 3'h5 == set_idx[2:0] ? enq_buffer_5_val_mask_1 : _GEN_3155; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3157 = 3'h6 == set_idx[2:0] ? enq_buffer_6_val_mask_1 : _GEN_3156; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3158 = 3'h7 == set_idx[2:0] ? enq_buffer_7_val_mask_1 : _GEN_3157; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3160 = 3'h1 == set_idx[2:0] ? enq_buffer_1_val_mask_2 : enq_buffer_0_val_mask_2; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3161 = 3'h2 == set_idx[2:0] ? enq_buffer_2_val_mask_2 : _GEN_3160; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3162 = 3'h3 == set_idx[2:0] ? enq_buffer_3_val_mask_2 : _GEN_3161; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3163 = 3'h4 == set_idx[2:0] ? enq_buffer_4_val_mask_2 : _GEN_3162; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3164 = 3'h5 == set_idx[2:0] ? enq_buffer_5_val_mask_2 : _GEN_3163; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3165 = 3'h6 == set_idx[2:0] ? enq_buffer_6_val_mask_2 : _GEN_3164; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3166 = 3'h7 == set_idx[2:0] ? enq_buffer_7_val_mask_2 : _GEN_3165; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3168 = 3'h1 == set_idx[2:0] ? enq_buffer_1_val_mask_3 : enq_buffer_0_val_mask_3; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3169 = 3'h2 == set_idx[2:0] ? enq_buffer_2_val_mask_3 : _GEN_3168; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3170 = 3'h3 == set_idx[2:0] ? enq_buffer_3_val_mask_3 : _GEN_3169; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3171 = 3'h4 == set_idx[2:0] ? enq_buffer_4_val_mask_3 : _GEN_3170; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3172 = 3'h5 == set_idx[2:0] ? enq_buffer_5_val_mask_3 : _GEN_3171; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3173 = 3'h6 == set_idx[2:0] ? enq_buffer_6_val_mask_3 : _GEN_3172; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3174 = 3'h7 == set_idx[2:0] ? enq_buffer_7_val_mask_3 : _GEN_3173; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3176 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_debug_tsrc : enq_buffer_0_dec_uops_0_debug_tsrc; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3177 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_debug_tsrc : _GEN_3176; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3178 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_debug_tsrc : _GEN_3177; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3179 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_debug_tsrc : _GEN_3178; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3180 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_debug_tsrc : _GEN_3179; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3181 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_debug_tsrc : _GEN_3180; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3182 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_debug_tsrc : _GEN_3181; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3184 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_debug_fsrc : enq_buffer_0_dec_uops_0_debug_fsrc; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3185 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_debug_fsrc : _GEN_3184; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3186 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_debug_fsrc : _GEN_3185; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3187 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_debug_fsrc : _GEN_3186; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3188 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_debug_fsrc : _GEN_3187; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3189 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_debug_fsrc : _GEN_3188; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3190 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_debug_fsrc : _GEN_3189; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3192 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_bp_xcpt_if : enq_buffer_0_dec_uops_0_bp_xcpt_if; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3193 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_bp_xcpt_if : _GEN_3192; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3194 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_bp_xcpt_if : _GEN_3193; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3195 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_bp_xcpt_if : _GEN_3194; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3196 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_bp_xcpt_if : _GEN_3195; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3197 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_bp_xcpt_if : _GEN_3196; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3198 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_bp_xcpt_if : _GEN_3197; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3200 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_bp_debug_if : enq_buffer_0_dec_uops_0_bp_debug_if; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3201 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_bp_debug_if : _GEN_3200; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3202 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_bp_debug_if : _GEN_3201; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3203 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_bp_debug_if : _GEN_3202; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3204 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_bp_debug_if : _GEN_3203; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3205 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_bp_debug_if : _GEN_3204; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3206 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_bp_debug_if : _GEN_3205; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3208 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_xcpt_ma_if : enq_buffer_0_dec_uops_0_xcpt_ma_if; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3209 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_xcpt_ma_if : _GEN_3208; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3210 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_xcpt_ma_if : _GEN_3209; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3211 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_xcpt_ma_if : _GEN_3210; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3212 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_xcpt_ma_if : _GEN_3211; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3213 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_xcpt_ma_if : _GEN_3212; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3214 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_xcpt_ma_if : _GEN_3213; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3216 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_xcpt_ae_if : enq_buffer_0_dec_uops_0_xcpt_ae_if; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3217 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_xcpt_ae_if : _GEN_3216; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3218 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_xcpt_ae_if : _GEN_3217; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3219 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_xcpt_ae_if : _GEN_3218; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3220 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_xcpt_ae_if : _GEN_3219; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3221 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_xcpt_ae_if : _GEN_3220; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3222 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_xcpt_ae_if : _GEN_3221; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3224 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_xcpt_pf_if : enq_buffer_0_dec_uops_0_xcpt_pf_if; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3225 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_xcpt_pf_if : _GEN_3224; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3226 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_xcpt_pf_if : _GEN_3225; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3227 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_xcpt_pf_if : _GEN_3226; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3228 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_xcpt_pf_if : _GEN_3227; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3229 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_xcpt_pf_if : _GEN_3228; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3230 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_xcpt_pf_if : _GEN_3229; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3232 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_fp_single : enq_buffer_0_dec_uops_0_fp_single; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3233 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_fp_single : _GEN_3232; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3234 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_fp_single : _GEN_3233; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3235 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_fp_single : _GEN_3234; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3236 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_fp_single : _GEN_3235; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3237 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_fp_single : _GEN_3236; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3238 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_fp_single : _GEN_3237; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3240 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_fp_val : enq_buffer_0_dec_uops_0_fp_val; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3241 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_fp_val : _GEN_3240; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3242 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_fp_val : _GEN_3241; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3243 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_fp_val : _GEN_3242; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3244 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_fp_val : _GEN_3243; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3245 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_fp_val : _GEN_3244; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3246 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_fp_val : _GEN_3245; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3248 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_frs3_en : enq_buffer_0_dec_uops_0_frs3_en; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3249 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_frs3_en : _GEN_3248; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3250 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_frs3_en : _GEN_3249; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3251 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_frs3_en : _GEN_3250; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3252 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_frs3_en : _GEN_3251; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3253 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_frs3_en : _GEN_3252; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3254 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_frs3_en : _GEN_3253; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3256 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_lrs2_rtype : enq_buffer_0_dec_uops_0_lrs2_rtype; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3257 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_lrs2_rtype : _GEN_3256; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3258 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_lrs2_rtype : _GEN_3257; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3259 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_lrs2_rtype : _GEN_3258; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3260 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_lrs2_rtype : _GEN_3259; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3261 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_lrs2_rtype : _GEN_3260; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3262 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_lrs2_rtype : _GEN_3261; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3264 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_lrs1_rtype : enq_buffer_0_dec_uops_0_lrs1_rtype; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3265 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_lrs1_rtype : _GEN_3264; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3266 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_lrs1_rtype : _GEN_3265; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3267 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_lrs1_rtype : _GEN_3266; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3268 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_lrs1_rtype : _GEN_3267; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3269 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_lrs1_rtype : _GEN_3268; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3270 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_lrs1_rtype : _GEN_3269; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3272 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_dst_rtype : enq_buffer_0_dec_uops_0_dst_rtype; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3273 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_dst_rtype : _GEN_3272; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3274 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_dst_rtype : _GEN_3273; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3275 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_dst_rtype : _GEN_3274; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3276 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_dst_rtype : _GEN_3275; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3277 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_dst_rtype : _GEN_3276; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3278 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_dst_rtype : _GEN_3277; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3280 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_ldst_val : enq_buffer_0_dec_uops_0_ldst_val; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3281 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_ldst_val : _GEN_3280; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3282 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_ldst_val : _GEN_3281; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3283 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_ldst_val : _GEN_3282; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3284 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_ldst_val : _GEN_3283; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3285 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_ldst_val : _GEN_3284; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3286 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_ldst_val : _GEN_3285; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3288 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_lrs3 : enq_buffer_0_dec_uops_0_lrs3; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3289 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_lrs3 : _GEN_3288; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3290 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_lrs3 : _GEN_3289; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3291 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_lrs3 : _GEN_3290; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3292 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_lrs3 : _GEN_3291; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3293 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_lrs3 : _GEN_3292; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3294 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_lrs3 : _GEN_3293; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3296 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_lrs2 : enq_buffer_0_dec_uops_0_lrs2; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3297 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_lrs2 : _GEN_3296; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3298 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_lrs2 : _GEN_3297; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3299 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_lrs2 : _GEN_3298; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3300 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_lrs2 : _GEN_3299; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3301 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_lrs2 : _GEN_3300; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3302 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_lrs2 : _GEN_3301; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3304 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_lrs1 : enq_buffer_0_dec_uops_0_lrs1; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3305 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_lrs1 : _GEN_3304; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3306 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_lrs1 : _GEN_3305; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3307 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_lrs1 : _GEN_3306; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3308 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_lrs1 : _GEN_3307; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3309 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_lrs1 : _GEN_3308; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3310 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_lrs1 : _GEN_3309; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3312 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_ldst : enq_buffer_0_dec_uops_0_ldst; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3313 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_ldst : _GEN_3312; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3314 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_ldst : _GEN_3313; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3315 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_ldst : _GEN_3314; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3316 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_ldst : _GEN_3315; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3317 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_ldst : _GEN_3316; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3318 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_ldst : _GEN_3317; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3320 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_ldst_is_rs1 : enq_buffer_0_dec_uops_0_ldst_is_rs1; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3321 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_ldst_is_rs1 : _GEN_3320; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3322 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_ldst_is_rs1 : _GEN_3321; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3323 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_ldst_is_rs1 : _GEN_3322; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3324 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_ldst_is_rs1 : _GEN_3323; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3325 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_ldst_is_rs1 : _GEN_3324; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3326 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_ldst_is_rs1 : _GEN_3325; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3328 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_flush_on_commit :
    enq_buffer_0_dec_uops_0_flush_on_commit; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3329 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_flush_on_commit : _GEN_3328; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3330 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_flush_on_commit : _GEN_3329; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3331 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_flush_on_commit : _GEN_3330; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3332 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_flush_on_commit : _GEN_3331; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3333 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_flush_on_commit : _GEN_3332; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3334 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_flush_on_commit : _GEN_3333; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3336 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_is_unique : enq_buffer_0_dec_uops_0_is_unique; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3337 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_is_unique : _GEN_3336; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3338 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_is_unique : _GEN_3337; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3339 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_is_unique : _GEN_3338; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3340 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_is_unique : _GEN_3339; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3341 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_is_unique : _GEN_3340; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3342 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_is_unique : _GEN_3341; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3344 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_is_sys_pc2epc : enq_buffer_0_dec_uops_0_is_sys_pc2epc
    ; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3345 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_is_sys_pc2epc : _GEN_3344; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3346 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_is_sys_pc2epc : _GEN_3345; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3347 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_is_sys_pc2epc : _GEN_3346; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3348 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_is_sys_pc2epc : _GEN_3347; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3349 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_is_sys_pc2epc : _GEN_3348; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3350 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_is_sys_pc2epc : _GEN_3349; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3352 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_uses_stq : enq_buffer_0_dec_uops_0_uses_stq; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3353 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_uses_stq : _GEN_3352; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3354 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_uses_stq : _GEN_3353; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3355 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_uses_stq : _GEN_3354; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3356 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_uses_stq : _GEN_3355; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3357 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_uses_stq : _GEN_3356; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3358 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_uses_stq : _GEN_3357; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3360 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_uses_ldq : enq_buffer_0_dec_uops_0_uses_ldq; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3361 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_uses_ldq : _GEN_3360; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3362 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_uses_ldq : _GEN_3361; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3363 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_uses_ldq : _GEN_3362; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3364 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_uses_ldq : _GEN_3363; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3365 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_uses_ldq : _GEN_3364; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3366 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_uses_ldq : _GEN_3365; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3368 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_is_amo : enq_buffer_0_dec_uops_0_is_amo; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3369 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_is_amo : _GEN_3368; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3370 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_is_amo : _GEN_3369; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3371 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_is_amo : _GEN_3370; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3372 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_is_amo : _GEN_3371; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3373 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_is_amo : _GEN_3372; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3374 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_is_amo : _GEN_3373; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3376 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_is_fencei : enq_buffer_0_dec_uops_0_is_fencei; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3377 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_is_fencei : _GEN_3376; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3378 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_is_fencei : _GEN_3377; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3379 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_is_fencei : _GEN_3378; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3380 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_is_fencei : _GEN_3379; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3381 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_is_fencei : _GEN_3380; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3382 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_is_fencei : _GEN_3381; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3384 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_is_fence : enq_buffer_0_dec_uops_0_is_fence; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3385 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_is_fence : _GEN_3384; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3386 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_is_fence : _GEN_3385; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3387 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_is_fence : _GEN_3386; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3388 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_is_fence : _GEN_3387; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3389 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_is_fence : _GEN_3388; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3390 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_is_fence : _GEN_3389; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3392 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_mem_signed : enq_buffer_0_dec_uops_0_mem_signed; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3393 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_mem_signed : _GEN_3392; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3394 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_mem_signed : _GEN_3393; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3395 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_mem_signed : _GEN_3394; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3396 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_mem_signed : _GEN_3395; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3397 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_mem_signed : _GEN_3396; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3398 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_mem_signed : _GEN_3397; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3400 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_mem_size : enq_buffer_0_dec_uops_0_mem_size; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3401 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_mem_size : _GEN_3400; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3402 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_mem_size : _GEN_3401; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3403 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_mem_size : _GEN_3402; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3404 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_mem_size : _GEN_3403; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3405 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_mem_size : _GEN_3404; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3406 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_mem_size : _GEN_3405; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3408 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_mem_cmd : enq_buffer_0_dec_uops_0_mem_cmd; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3409 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_mem_cmd : _GEN_3408; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3410 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_mem_cmd : _GEN_3409; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3411 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_mem_cmd : _GEN_3410; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3412 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_mem_cmd : _GEN_3411; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3413 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_mem_cmd : _GEN_3412; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3414 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_mem_cmd : _GEN_3413; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3416 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_bypassable : enq_buffer_0_dec_uops_0_bypassable; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3417 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_bypassable : _GEN_3416; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3418 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_bypassable : _GEN_3417; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3419 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_bypassable : _GEN_3418; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3420 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_bypassable : _GEN_3419; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3421 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_bypassable : _GEN_3420; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3422 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_bypassable : _GEN_3421; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_3424 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_exc_cause : enq_buffer_0_dec_uops_0_exc_cause; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_3425 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_exc_cause : _GEN_3424; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_3426 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_exc_cause : _GEN_3425; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_3427 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_exc_cause : _GEN_3426; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_3428 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_exc_cause : _GEN_3427; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_3429 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_exc_cause : _GEN_3428; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_3430 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_exc_cause : _GEN_3429; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3432 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_exception : enq_buffer_0_dec_uops_0_exception; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3433 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_exception : _GEN_3432; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3434 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_exception : _GEN_3433; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3435 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_exception : _GEN_3434; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3436 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_exception : _GEN_3435; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3437 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_exception : _GEN_3436; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3438 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_exception : _GEN_3437; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3440 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_stale_pdst : enq_buffer_0_dec_uops_0_stale_pdst; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3441 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_stale_pdst : _GEN_3440; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3442 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_stale_pdst : _GEN_3441; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3443 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_stale_pdst : _GEN_3442; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3444 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_stale_pdst : _GEN_3443; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3445 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_stale_pdst : _GEN_3444; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3446 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_stale_pdst : _GEN_3445; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3448 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_ppred_busy : enq_buffer_0_dec_uops_0_ppred_busy; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3449 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_ppred_busy : _GEN_3448; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3450 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_ppred_busy : _GEN_3449; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3451 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_ppred_busy : _GEN_3450; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3452 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_ppred_busy : _GEN_3451; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3453 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_ppred_busy : _GEN_3452; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3454 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_ppred_busy : _GEN_3453; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3456 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_prs3_busy : enq_buffer_0_dec_uops_0_prs3_busy; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3457 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_prs3_busy : _GEN_3456; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3458 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_prs3_busy : _GEN_3457; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3459 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_prs3_busy : _GEN_3458; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3460 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_prs3_busy : _GEN_3459; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3461 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_prs3_busy : _GEN_3460; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3462 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_prs3_busy : _GEN_3461; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3464 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_prs2_busy : enq_buffer_0_dec_uops_0_prs2_busy; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3465 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_prs2_busy : _GEN_3464; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3466 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_prs2_busy : _GEN_3465; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3467 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_prs2_busy : _GEN_3466; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3468 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_prs2_busy : _GEN_3467; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3469 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_prs2_busy : _GEN_3468; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3470 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_prs2_busy : _GEN_3469; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3472 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_prs1_busy : enq_buffer_0_dec_uops_0_prs1_busy; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3473 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_prs1_busy : _GEN_3472; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3474 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_prs1_busy : _GEN_3473; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3475 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_prs1_busy : _GEN_3474; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3476 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_prs1_busy : _GEN_3475; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3477 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_prs1_busy : _GEN_3476; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3478 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_prs1_busy : _GEN_3477; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3480 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_ppred : enq_buffer_0_dec_uops_0_ppred; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3481 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_ppred : _GEN_3480; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3482 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_ppred : _GEN_3481; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3483 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_ppred : _GEN_3482; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3484 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_ppred : _GEN_3483; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3485 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_ppred : _GEN_3484; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3486 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_ppred : _GEN_3485; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3488 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_prs3 : enq_buffer_0_dec_uops_0_prs3; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3489 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_prs3 : _GEN_3488; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3490 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_prs3 : _GEN_3489; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3491 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_prs3 : _GEN_3490; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3492 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_prs3 : _GEN_3491; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3493 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_prs3 : _GEN_3492; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3494 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_prs3 : _GEN_3493; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3496 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_prs2 : enq_buffer_0_dec_uops_0_prs2; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3497 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_prs2 : _GEN_3496; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3498 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_prs2 : _GEN_3497; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3499 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_prs2 : _GEN_3498; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3500 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_prs2 : _GEN_3499; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3501 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_prs2 : _GEN_3500; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3502 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_prs2 : _GEN_3501; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3504 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_prs1 : enq_buffer_0_dec_uops_0_prs1; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3505 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_prs1 : _GEN_3504; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3506 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_prs1 : _GEN_3505; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3507 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_prs1 : _GEN_3506; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3508 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_prs1 : _GEN_3507; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3509 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_prs1 : _GEN_3508; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3510 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_prs1 : _GEN_3509; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3512 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_pdst : enq_buffer_0_dec_uops_0_pdst; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3513 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_pdst : _GEN_3512; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3514 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_pdst : _GEN_3513; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3515 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_pdst : _GEN_3514; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3516 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_pdst : _GEN_3515; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3517 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_pdst : _GEN_3516; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3518 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_pdst : _GEN_3517; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3520 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_rxq_idx : enq_buffer_0_dec_uops_0_rxq_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3521 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_rxq_idx : _GEN_3520; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3522 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_rxq_idx : _GEN_3521; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3523 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_rxq_idx : _GEN_3522; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3524 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_rxq_idx : _GEN_3523; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3525 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_rxq_idx : _GEN_3524; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3526 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_rxq_idx : _GEN_3525; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3528 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_stq_idx : enq_buffer_0_dec_uops_0_stq_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3529 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_stq_idx : _GEN_3528; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3530 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_stq_idx : _GEN_3529; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3531 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_stq_idx : _GEN_3530; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3532 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_stq_idx : _GEN_3531; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3533 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_stq_idx : _GEN_3532; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3534 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_stq_idx : _GEN_3533; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3536 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_ldq_idx : enq_buffer_0_dec_uops_0_ldq_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3537 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_ldq_idx : _GEN_3536; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3538 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_ldq_idx : _GEN_3537; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3539 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_ldq_idx : _GEN_3538; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3540 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_ldq_idx : _GEN_3539; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3541 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_ldq_idx : _GEN_3540; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3542 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_ldq_idx : _GEN_3541; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3544 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_rob_idx : enq_buffer_0_dec_uops_0_rob_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3545 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_rob_idx : _GEN_3544; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3546 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_rob_idx : _GEN_3545; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3547 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_rob_idx : _GEN_3546; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3548 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_rob_idx : _GEN_3547; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3549 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_rob_idx : _GEN_3548; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3550 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_rob_idx : _GEN_3549; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_3552 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_csr_addr : enq_buffer_0_dec_uops_0_csr_addr; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_3553 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_csr_addr : _GEN_3552; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_3554 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_csr_addr : _GEN_3553; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_3555 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_csr_addr : _GEN_3554; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_3556 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_csr_addr : _GEN_3555; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_3557 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_csr_addr : _GEN_3556; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_3558 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_csr_addr : _GEN_3557; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_3560 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_imm_packed : enq_buffer_0_dec_uops_0_imm_packed
    ; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_3561 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_imm_packed : _GEN_3560; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_3562 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_imm_packed : _GEN_3561; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_3563 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_imm_packed : _GEN_3562; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_3564 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_imm_packed : _GEN_3563; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_3565 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_imm_packed : _GEN_3564; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_3566 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_imm_packed : _GEN_3565; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3568 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_taken : enq_buffer_0_dec_uops_0_taken; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3569 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_taken : _GEN_3568; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3570 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_taken : _GEN_3569; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3571 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_taken : _GEN_3570; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3572 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_taken : _GEN_3571; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3573 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_taken : _GEN_3572; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3574 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_taken : _GEN_3573; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3576 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_pc_lob : enq_buffer_0_dec_uops_0_pc_lob; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3577 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_pc_lob : _GEN_3576; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3578 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_pc_lob : _GEN_3577; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3579 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_pc_lob : _GEN_3578; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3580 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_pc_lob : _GEN_3579; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3581 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_pc_lob : _GEN_3580; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3582 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_pc_lob : _GEN_3581; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3584 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_edge_inst : enq_buffer_0_dec_uops_0_edge_inst; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3585 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_edge_inst : _GEN_3584; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3586 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_edge_inst : _GEN_3585; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3587 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_edge_inst : _GEN_3586; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3588 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_edge_inst : _GEN_3587; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3589 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_edge_inst : _GEN_3588; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3590 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_edge_inst : _GEN_3589; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3592 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_ftq_idx : enq_buffer_0_dec_uops_0_ftq_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3593 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_ftq_idx : _GEN_3592; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3594 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_ftq_idx : _GEN_3593; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3595 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_ftq_idx : _GEN_3594; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3596 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_ftq_idx : _GEN_3595; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3597 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_ftq_idx : _GEN_3596; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_3598 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_ftq_idx : _GEN_3597; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3600 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_br_tag : enq_buffer_0_dec_uops_0_br_tag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3601 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_br_tag : _GEN_3600; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3602 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_br_tag : _GEN_3601; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3603 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_br_tag : _GEN_3602; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3604 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_br_tag : _GEN_3603; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3605 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_br_tag : _GEN_3604; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3606 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_br_tag : _GEN_3605; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_3608 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_br_mask : enq_buffer_0_dec_uops_0_br_mask; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_3609 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_br_mask : _GEN_3608; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_3610 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_br_mask : _GEN_3609; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_3611 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_br_mask : _GEN_3610; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_3612 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_br_mask : _GEN_3611; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_3613 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_br_mask : _GEN_3612; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_3614 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_br_mask : _GEN_3613; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3616 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_is_sfb : enq_buffer_0_dec_uops_0_is_sfb; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3617 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_is_sfb : _GEN_3616; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3618 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_is_sfb : _GEN_3617; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3619 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_is_sfb : _GEN_3618; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3620 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_is_sfb : _GEN_3619; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3621 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_is_sfb : _GEN_3620; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3622 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_is_sfb : _GEN_3621; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3624 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_is_jal : enq_buffer_0_dec_uops_0_is_jal; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3625 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_is_jal : _GEN_3624; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3626 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_is_jal : _GEN_3625; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3627 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_is_jal : _GEN_3626; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3628 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_is_jal : _GEN_3627; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3629 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_is_jal : _GEN_3628; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3630 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_is_jal : _GEN_3629; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3632 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_is_jalr : enq_buffer_0_dec_uops_0_is_jalr; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3633 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_is_jalr : _GEN_3632; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3634 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_is_jalr : _GEN_3633; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3635 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_is_jalr : _GEN_3634; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3636 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_is_jalr : _GEN_3635; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3637 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_is_jalr : _GEN_3636; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3638 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_is_jalr : _GEN_3637; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3640 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_is_br : enq_buffer_0_dec_uops_0_is_br; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3641 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_is_br : _GEN_3640; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3642 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_is_br : _GEN_3641; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3643 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_is_br : _GEN_3642; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3644 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_is_br : _GEN_3643; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3645 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_is_br : _GEN_3644; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3646 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_is_br : _GEN_3645; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3648 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_iw_p2_poisoned :
    enq_buffer_0_dec_uops_0_iw_p2_poisoned; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3649 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_iw_p2_poisoned : _GEN_3648; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3650 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_iw_p2_poisoned : _GEN_3649; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3651 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_iw_p2_poisoned : _GEN_3650; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3652 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_iw_p2_poisoned : _GEN_3651; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3653 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_iw_p2_poisoned : _GEN_3652; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3654 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_iw_p2_poisoned : _GEN_3653; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3656 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_iw_p1_poisoned :
    enq_buffer_0_dec_uops_0_iw_p1_poisoned; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3657 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_iw_p1_poisoned : _GEN_3656; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3658 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_iw_p1_poisoned : _GEN_3657; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3659 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_iw_p1_poisoned : _GEN_3658; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3660 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_iw_p1_poisoned : _GEN_3659; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3661 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_iw_p1_poisoned : _GEN_3660; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3662 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_iw_p1_poisoned : _GEN_3661; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3664 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_iw_state : enq_buffer_0_dec_uops_0_iw_state; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3665 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_iw_state : _GEN_3664; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3666 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_iw_state : _GEN_3665; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3667 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_iw_state : _GEN_3666; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3668 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_iw_state : _GEN_3667; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3669 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_iw_state : _GEN_3668; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3670 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_iw_state : _GEN_3669; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3672 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_ctrl_op3_sel :
    enq_buffer_0_dec_uops_0_ctrl_op3_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3673 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_ctrl_op3_sel : _GEN_3672; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3674 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_ctrl_op3_sel : _GEN_3673; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3675 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_ctrl_op3_sel : _GEN_3674; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3676 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_ctrl_op3_sel : _GEN_3675; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3677 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_ctrl_op3_sel : _GEN_3676; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3678 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_ctrl_op3_sel : _GEN_3677; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3680 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_ctrl_is_std : enq_buffer_0_dec_uops_0_ctrl_is_std; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3681 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_ctrl_is_std : _GEN_3680; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3682 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_ctrl_is_std : _GEN_3681; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3683 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_ctrl_is_std : _GEN_3682; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3684 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_ctrl_is_std : _GEN_3683; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3685 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_ctrl_is_std : _GEN_3684; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3686 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_ctrl_is_std : _GEN_3685; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3688 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_ctrl_is_sta : enq_buffer_0_dec_uops_0_ctrl_is_sta; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3689 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_ctrl_is_sta : _GEN_3688; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3690 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_ctrl_is_sta : _GEN_3689; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3691 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_ctrl_is_sta : _GEN_3690; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3692 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_ctrl_is_sta : _GEN_3691; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3693 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_ctrl_is_sta : _GEN_3692; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3694 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_ctrl_is_sta : _GEN_3693; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3696 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_ctrl_is_load : enq_buffer_0_dec_uops_0_ctrl_is_load; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3697 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_ctrl_is_load : _GEN_3696; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3698 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_ctrl_is_load : _GEN_3697; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3699 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_ctrl_is_load : _GEN_3698; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3700 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_ctrl_is_load : _GEN_3699; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3701 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_ctrl_is_load : _GEN_3700; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3702 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_ctrl_is_load : _GEN_3701; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3704 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_ctrl_csr_cmd :
    enq_buffer_0_dec_uops_0_ctrl_csr_cmd; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3705 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_ctrl_csr_cmd : _GEN_3704; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3706 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_ctrl_csr_cmd : _GEN_3705; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3707 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_ctrl_csr_cmd : _GEN_3706; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3708 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_ctrl_csr_cmd : _GEN_3707; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3709 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_ctrl_csr_cmd : _GEN_3708; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3710 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_ctrl_csr_cmd : _GEN_3709; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3712 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_ctrl_fcn_dw : enq_buffer_0_dec_uops_0_ctrl_fcn_dw; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3713 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_ctrl_fcn_dw : _GEN_3712; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3714 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_ctrl_fcn_dw : _GEN_3713; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3715 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_ctrl_fcn_dw : _GEN_3714; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3716 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_ctrl_fcn_dw : _GEN_3715; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3717 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_ctrl_fcn_dw : _GEN_3716; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3718 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_ctrl_fcn_dw : _GEN_3717; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3720 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_ctrl_op_fcn :
    enq_buffer_0_dec_uops_0_ctrl_op_fcn; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3721 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_ctrl_op_fcn : _GEN_3720; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3722 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_ctrl_op_fcn : _GEN_3721; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3723 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_ctrl_op_fcn : _GEN_3722; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3724 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_ctrl_op_fcn : _GEN_3723; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3725 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_ctrl_op_fcn : _GEN_3724; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3726 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_ctrl_op_fcn : _GEN_3725; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3728 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_ctrl_imm_sel :
    enq_buffer_0_dec_uops_0_ctrl_imm_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3729 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_ctrl_imm_sel : _GEN_3728; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3730 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_ctrl_imm_sel : _GEN_3729; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3731 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_ctrl_imm_sel : _GEN_3730; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3732 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_ctrl_imm_sel : _GEN_3731; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3733 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_ctrl_imm_sel : _GEN_3732; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3734 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_ctrl_imm_sel : _GEN_3733; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3736 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_ctrl_op2_sel :
    enq_buffer_0_dec_uops_0_ctrl_op2_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3737 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_ctrl_op2_sel : _GEN_3736; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3738 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_ctrl_op2_sel : _GEN_3737; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3739 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_ctrl_op2_sel : _GEN_3738; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3740 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_ctrl_op2_sel : _GEN_3739; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3741 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_ctrl_op2_sel : _GEN_3740; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3742 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_ctrl_op2_sel : _GEN_3741; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3744 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_ctrl_op1_sel :
    enq_buffer_0_dec_uops_0_ctrl_op1_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3745 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_ctrl_op1_sel : _GEN_3744; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3746 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_ctrl_op1_sel : _GEN_3745; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3747 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_ctrl_op1_sel : _GEN_3746; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3748 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_ctrl_op1_sel : _GEN_3747; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3749 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_ctrl_op1_sel : _GEN_3748; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3750 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_ctrl_op1_sel : _GEN_3749; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3752 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_ctrl_br_type :
    enq_buffer_0_dec_uops_0_ctrl_br_type; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3753 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_ctrl_br_type : _GEN_3752; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3754 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_ctrl_br_type : _GEN_3753; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3755 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_ctrl_br_type : _GEN_3754; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3756 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_ctrl_br_type : _GEN_3755; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3757 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_ctrl_br_type : _GEN_3756; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3758 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_ctrl_br_type : _GEN_3757; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_3760 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_fu_code : enq_buffer_0_dec_uops_0_fu_code; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_3761 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_fu_code : _GEN_3760; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_3762 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_fu_code : _GEN_3761; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_3763 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_fu_code : _GEN_3762; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_3764 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_fu_code : _GEN_3763; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_3765 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_fu_code : _GEN_3764; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_3766 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_fu_code : _GEN_3765; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3768 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_iq_type : enq_buffer_0_dec_uops_0_iq_type; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3769 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_iq_type : _GEN_3768; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3770 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_iq_type : _GEN_3769; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3771 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_iq_type : _GEN_3770; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3772 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_iq_type : _GEN_3771; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3773 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_iq_type : _GEN_3772; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3774 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_iq_type : _GEN_3773; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_3776 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_debug_pc : enq_buffer_0_dec_uops_0_debug_pc; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_3777 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_debug_pc : _GEN_3776; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_3778 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_debug_pc : _GEN_3777; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_3779 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_debug_pc : _GEN_3778; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_3780 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_debug_pc : _GEN_3779; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_3781 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_debug_pc : _GEN_3780; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_3782 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_debug_pc : _GEN_3781; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3784 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_is_rvc : enq_buffer_0_dec_uops_0_is_rvc; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3785 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_is_rvc : _GEN_3784; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3786 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_is_rvc : _GEN_3785; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3787 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_is_rvc : _GEN_3786; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3788 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_is_rvc : _GEN_3787; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3789 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_is_rvc : _GEN_3788; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3790 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_is_rvc : _GEN_3789; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_3792 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_debug_inst : enq_buffer_0_dec_uops_0_debug_inst
    ; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_3793 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_debug_inst : _GEN_3792; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_3794 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_debug_inst : _GEN_3793; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_3795 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_debug_inst : _GEN_3794; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_3796 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_debug_inst : _GEN_3795; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_3797 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_debug_inst : _GEN_3796; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_3798 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_debug_inst : _GEN_3797; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_3800 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_inst : enq_buffer_0_dec_uops_0_inst; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_3801 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_inst : _GEN_3800; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_3802 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_inst : _GEN_3801; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_3803 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_inst : _GEN_3802; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_3804 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_inst : _GEN_3803; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_3805 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_inst : _GEN_3804; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_3806 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_inst : _GEN_3805; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3808 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_uopc : enq_buffer_0_dec_uops_0_uopc; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3809 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_uopc : _GEN_3808; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3810 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_uopc : _GEN_3809; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3811 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_uopc : _GEN_3810; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3812 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_uopc : _GEN_3811; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3813 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_uopc : _GEN_3812; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_3814 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_uopc : _GEN_3813; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3816 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_address_num :
    enq_buffer_0_dec_uops_0_address_num; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3817 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_address_num : _GEN_3816; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3818 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_address_num : _GEN_3817; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3819 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_address_num : _GEN_3818; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3820 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_address_num : _GEN_3819; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3821 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_address_num : _GEN_3820; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3822 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_address_num : _GEN_3821; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3824 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_rob_inst_idx :
    enq_buffer_0_dec_uops_0_rob_inst_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3825 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_rob_inst_idx : _GEN_3824; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3826 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_rob_inst_idx : _GEN_3825; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3827 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_rob_inst_idx : _GEN_3826; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3828 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_rob_inst_idx : _GEN_3827; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3829 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_rob_inst_idx : _GEN_3828; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3830 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_rob_inst_idx : _GEN_3829; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3832 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_self_index : enq_buffer_0_dec_uops_0_self_index; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3833 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_self_index : _GEN_3832; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3834 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_self_index : _GEN_3833; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3835 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_self_index : _GEN_3834; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3836 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_self_index : _GEN_3835; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3837 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_self_index : _GEN_3836; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3838 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_self_index : _GEN_3837; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3840 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_split_num : enq_buffer_0_dec_uops_0_split_num; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3841 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_split_num : _GEN_3840; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3842 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_split_num : _GEN_3841; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3843 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_split_num : _GEN_3842; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3844 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_split_num : _GEN_3843; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3845 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_split_num : _GEN_3844; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_3846 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_split_num : _GEN_3845; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3848 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_op2_sel : enq_buffer_0_dec_uops_0_op2_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3849 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_op2_sel : _GEN_3848; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3850 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_op2_sel : _GEN_3849; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3851 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_op2_sel : _GEN_3850; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3852 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_op2_sel : _GEN_3851; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3853 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_op2_sel : _GEN_3852; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3854 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_op2_sel : _GEN_3853; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3856 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_op1_sel : enq_buffer_0_dec_uops_0_op1_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3857 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_op1_sel : _GEN_3856; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3858 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_op1_sel : _GEN_3857; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3859 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_op1_sel : _GEN_3858; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3860 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_op1_sel : _GEN_3859; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3861 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_op1_sel : _GEN_3860; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3862 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_op1_sel : _GEN_3861; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3864 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_stale_pflag :
    enq_buffer_0_dec_uops_0_stale_pflag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3865 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_stale_pflag : _GEN_3864; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3866 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_stale_pflag : _GEN_3865; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3867 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_stale_pflag : _GEN_3866; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3868 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_stale_pflag : _GEN_3867; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3869 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_stale_pflag : _GEN_3868; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3870 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_stale_pflag : _GEN_3869; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3872 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_pflag_busy : enq_buffer_0_dec_uops_0_pflag_busy; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3873 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_pflag_busy : _GEN_3872; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3874 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_pflag_busy : _GEN_3873; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3875 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_pflag_busy : _GEN_3874; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3876 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_pflag_busy : _GEN_3875; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3877 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_pflag_busy : _GEN_3876; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3878 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_pflag_busy : _GEN_3877; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3880 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_pwflag : enq_buffer_0_dec_uops_0_pwflag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3881 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_pwflag : _GEN_3880; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3882 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_pwflag : _GEN_3881; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3883 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_pwflag : _GEN_3882; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3884 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_pwflag : _GEN_3883; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3885 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_pwflag : _GEN_3884; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3886 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_pwflag : _GEN_3885; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3888 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_prflag : enq_buffer_0_dec_uops_0_prflag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3889 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_prflag : _GEN_3888; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3890 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_prflag : _GEN_3889; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3891 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_prflag : _GEN_3890; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3892 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_prflag : _GEN_3891; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3893 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_prflag : _GEN_3892; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_3894 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_prflag : _GEN_3893; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3896 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_wflag : enq_buffer_0_dec_uops_0_wflag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3897 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_wflag : _GEN_3896; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3898 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_wflag : _GEN_3897; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3899 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_wflag : _GEN_3898; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3900 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_wflag : _GEN_3899; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3901 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_wflag : _GEN_3900; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3902 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_wflag : _GEN_3901; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3904 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_rflag : enq_buffer_0_dec_uops_0_rflag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3905 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_rflag : _GEN_3904; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3906 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_rflag : _GEN_3905; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3907 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_rflag : _GEN_3906; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3908 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_rflag : _GEN_3907; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3909 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_rflag : _GEN_3908; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3910 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_rflag : _GEN_3909; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3912 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_lrs3_rtype : enq_buffer_0_dec_uops_0_lrs3_rtype; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3913 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_lrs3_rtype : _GEN_3912; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3914 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_lrs3_rtype : _GEN_3913; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3915 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_lrs3_rtype : _GEN_3914; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3916 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_lrs3_rtype : _GEN_3915; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3917 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_lrs3_rtype : _GEN_3916; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3918 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_lrs3_rtype : _GEN_3917; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3920 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_shift : enq_buffer_0_dec_uops_0_shift; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3921 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_shift : _GEN_3920; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3922 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_shift : _GEN_3921; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3923 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_shift : _GEN_3922; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3924 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_shift : _GEN_3923; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3925 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_shift : _GEN_3924; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_3926 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_shift : _GEN_3925; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3928 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_is_unicore : enq_buffer_0_dec_uops_0_is_unicore; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3929 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_is_unicore : _GEN_3928; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3930 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_is_unicore : _GEN_3929; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3931 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_is_unicore : _GEN_3930; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3932 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_is_unicore : _GEN_3931; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3933 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_is_unicore : _GEN_3932; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3934 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_is_unicore : _GEN_3933; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3936 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_switch_off : enq_buffer_0_dec_uops_0_switch_off; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3937 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_switch_off : _GEN_3936; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3938 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_switch_off : _GEN_3937; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3939 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_switch_off : _GEN_3938; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3940 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_switch_off : _GEN_3939; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3941 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_switch_off : _GEN_3940; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3942 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_switch_off : _GEN_3941; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3944 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_0_switch : enq_buffer_0_dec_uops_0_switch; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3945 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_0_switch : _GEN_3944; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3946 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_0_switch : _GEN_3945; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3947 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_0_switch : _GEN_3946; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3948 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_0_switch : _GEN_3947; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3949 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_0_switch : _GEN_3948; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3950 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_0_switch : _GEN_3949; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3952 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_debug_tsrc : enq_buffer_0_dec_uops_1_debug_tsrc; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3953 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_debug_tsrc : _GEN_3952; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3954 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_debug_tsrc : _GEN_3953; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3955 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_debug_tsrc : _GEN_3954; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3956 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_debug_tsrc : _GEN_3955; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3957 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_debug_tsrc : _GEN_3956; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3958 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_debug_tsrc : _GEN_3957; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3960 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_debug_fsrc : enq_buffer_0_dec_uops_1_debug_fsrc; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3961 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_debug_fsrc : _GEN_3960; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3962 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_debug_fsrc : _GEN_3961; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3963 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_debug_fsrc : _GEN_3962; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3964 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_debug_fsrc : _GEN_3963; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3965 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_debug_fsrc : _GEN_3964; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_3966 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_debug_fsrc : _GEN_3965; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3968 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_bp_xcpt_if : enq_buffer_0_dec_uops_1_bp_xcpt_if; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3969 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_bp_xcpt_if : _GEN_3968; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3970 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_bp_xcpt_if : _GEN_3969; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3971 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_bp_xcpt_if : _GEN_3970; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3972 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_bp_xcpt_if : _GEN_3971; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3973 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_bp_xcpt_if : _GEN_3972; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3974 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_bp_xcpt_if : _GEN_3973; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3976 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_bp_debug_if : enq_buffer_0_dec_uops_1_bp_debug_if; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3977 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_bp_debug_if : _GEN_3976; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3978 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_bp_debug_if : _GEN_3977; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3979 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_bp_debug_if : _GEN_3978; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3980 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_bp_debug_if : _GEN_3979; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3981 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_bp_debug_if : _GEN_3980; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3982 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_bp_debug_if : _GEN_3981; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3984 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_xcpt_ma_if : enq_buffer_0_dec_uops_1_xcpt_ma_if; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3985 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_xcpt_ma_if : _GEN_3984; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3986 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_xcpt_ma_if : _GEN_3985; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3987 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_xcpt_ma_if : _GEN_3986; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3988 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_xcpt_ma_if : _GEN_3987; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3989 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_xcpt_ma_if : _GEN_3988; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3990 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_xcpt_ma_if : _GEN_3989; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3992 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_xcpt_ae_if : enq_buffer_0_dec_uops_1_xcpt_ae_if; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3993 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_xcpt_ae_if : _GEN_3992; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3994 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_xcpt_ae_if : _GEN_3993; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3995 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_xcpt_ae_if : _GEN_3994; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3996 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_xcpt_ae_if : _GEN_3995; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3997 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_xcpt_ae_if : _GEN_3996; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_3998 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_xcpt_ae_if : _GEN_3997; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4000 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_xcpt_pf_if : enq_buffer_0_dec_uops_1_xcpt_pf_if; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4001 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_xcpt_pf_if : _GEN_4000; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4002 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_xcpt_pf_if : _GEN_4001; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4003 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_xcpt_pf_if : _GEN_4002; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4004 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_xcpt_pf_if : _GEN_4003; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4005 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_xcpt_pf_if : _GEN_4004; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4006 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_xcpt_pf_if : _GEN_4005; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4008 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_fp_single : enq_buffer_0_dec_uops_1_fp_single; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4009 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_fp_single : _GEN_4008; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4010 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_fp_single : _GEN_4009; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4011 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_fp_single : _GEN_4010; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4012 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_fp_single : _GEN_4011; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4013 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_fp_single : _GEN_4012; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4014 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_fp_single : _GEN_4013; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4016 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_fp_val : enq_buffer_0_dec_uops_1_fp_val; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4017 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_fp_val : _GEN_4016; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4018 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_fp_val : _GEN_4017; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4019 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_fp_val : _GEN_4018; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4020 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_fp_val : _GEN_4019; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4021 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_fp_val : _GEN_4020; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4022 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_fp_val : _GEN_4021; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4024 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_frs3_en : enq_buffer_0_dec_uops_1_frs3_en; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4025 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_frs3_en : _GEN_4024; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4026 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_frs3_en : _GEN_4025; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4027 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_frs3_en : _GEN_4026; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4028 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_frs3_en : _GEN_4027; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4029 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_frs3_en : _GEN_4028; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4030 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_frs3_en : _GEN_4029; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4032 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_lrs2_rtype : enq_buffer_0_dec_uops_1_lrs2_rtype; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4033 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_lrs2_rtype : _GEN_4032; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4034 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_lrs2_rtype : _GEN_4033; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4035 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_lrs2_rtype : _GEN_4034; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4036 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_lrs2_rtype : _GEN_4035; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4037 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_lrs2_rtype : _GEN_4036; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4038 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_lrs2_rtype : _GEN_4037; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4040 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_lrs1_rtype : enq_buffer_0_dec_uops_1_lrs1_rtype; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4041 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_lrs1_rtype : _GEN_4040; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4042 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_lrs1_rtype : _GEN_4041; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4043 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_lrs1_rtype : _GEN_4042; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4044 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_lrs1_rtype : _GEN_4043; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4045 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_lrs1_rtype : _GEN_4044; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4046 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_lrs1_rtype : _GEN_4045; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4048 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_dst_rtype : enq_buffer_0_dec_uops_1_dst_rtype; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4049 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_dst_rtype : _GEN_4048; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4050 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_dst_rtype : _GEN_4049; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4051 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_dst_rtype : _GEN_4050; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4052 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_dst_rtype : _GEN_4051; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4053 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_dst_rtype : _GEN_4052; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4054 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_dst_rtype : _GEN_4053; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4056 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_ldst_val : enq_buffer_0_dec_uops_1_ldst_val; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4057 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_ldst_val : _GEN_4056; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4058 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_ldst_val : _GEN_4057; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4059 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_ldst_val : _GEN_4058; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4060 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_ldst_val : _GEN_4059; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4061 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_ldst_val : _GEN_4060; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4062 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_ldst_val : _GEN_4061; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4064 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_lrs3 : enq_buffer_0_dec_uops_1_lrs3; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4065 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_lrs3 : _GEN_4064; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4066 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_lrs3 : _GEN_4065; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4067 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_lrs3 : _GEN_4066; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4068 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_lrs3 : _GEN_4067; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4069 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_lrs3 : _GEN_4068; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4070 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_lrs3 : _GEN_4069; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4072 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_lrs2 : enq_buffer_0_dec_uops_1_lrs2; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4073 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_lrs2 : _GEN_4072; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4074 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_lrs2 : _GEN_4073; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4075 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_lrs2 : _GEN_4074; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4076 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_lrs2 : _GEN_4075; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4077 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_lrs2 : _GEN_4076; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4078 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_lrs2 : _GEN_4077; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4080 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_lrs1 : enq_buffer_0_dec_uops_1_lrs1; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4081 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_lrs1 : _GEN_4080; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4082 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_lrs1 : _GEN_4081; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4083 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_lrs1 : _GEN_4082; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4084 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_lrs1 : _GEN_4083; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4085 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_lrs1 : _GEN_4084; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4086 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_lrs1 : _GEN_4085; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4088 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_ldst : enq_buffer_0_dec_uops_1_ldst; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4089 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_ldst : _GEN_4088; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4090 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_ldst : _GEN_4089; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4091 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_ldst : _GEN_4090; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4092 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_ldst : _GEN_4091; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4093 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_ldst : _GEN_4092; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4094 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_ldst : _GEN_4093; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4096 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_ldst_is_rs1 : enq_buffer_0_dec_uops_1_ldst_is_rs1; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4097 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_ldst_is_rs1 : _GEN_4096; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4098 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_ldst_is_rs1 : _GEN_4097; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4099 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_ldst_is_rs1 : _GEN_4098; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4100 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_ldst_is_rs1 : _GEN_4099; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4101 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_ldst_is_rs1 : _GEN_4100; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4102 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_ldst_is_rs1 : _GEN_4101; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4104 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_flush_on_commit :
    enq_buffer_0_dec_uops_1_flush_on_commit; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4105 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_flush_on_commit : _GEN_4104; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4106 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_flush_on_commit : _GEN_4105; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4107 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_flush_on_commit : _GEN_4106; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4108 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_flush_on_commit : _GEN_4107; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4109 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_flush_on_commit : _GEN_4108; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4110 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_flush_on_commit : _GEN_4109; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4112 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_is_unique : enq_buffer_0_dec_uops_1_is_unique; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4113 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_is_unique : _GEN_4112; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4114 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_is_unique : _GEN_4113; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4115 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_is_unique : _GEN_4114; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4116 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_is_unique : _GEN_4115; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4117 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_is_unique : _GEN_4116; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4118 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_is_unique : _GEN_4117; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4120 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_is_sys_pc2epc : enq_buffer_0_dec_uops_1_is_sys_pc2epc
    ; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4121 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_is_sys_pc2epc : _GEN_4120; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4122 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_is_sys_pc2epc : _GEN_4121; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4123 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_is_sys_pc2epc : _GEN_4122; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4124 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_is_sys_pc2epc : _GEN_4123; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4125 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_is_sys_pc2epc : _GEN_4124; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4126 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_is_sys_pc2epc : _GEN_4125; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4128 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_uses_stq : enq_buffer_0_dec_uops_1_uses_stq; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4129 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_uses_stq : _GEN_4128; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4130 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_uses_stq : _GEN_4129; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4131 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_uses_stq : _GEN_4130; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4132 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_uses_stq : _GEN_4131; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4133 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_uses_stq : _GEN_4132; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4134 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_uses_stq : _GEN_4133; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4136 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_uses_ldq : enq_buffer_0_dec_uops_1_uses_ldq; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4137 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_uses_ldq : _GEN_4136; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4138 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_uses_ldq : _GEN_4137; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4139 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_uses_ldq : _GEN_4138; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4140 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_uses_ldq : _GEN_4139; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4141 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_uses_ldq : _GEN_4140; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4142 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_uses_ldq : _GEN_4141; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4144 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_is_amo : enq_buffer_0_dec_uops_1_is_amo; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4145 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_is_amo : _GEN_4144; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4146 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_is_amo : _GEN_4145; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4147 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_is_amo : _GEN_4146; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4148 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_is_amo : _GEN_4147; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4149 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_is_amo : _GEN_4148; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4150 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_is_amo : _GEN_4149; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4152 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_is_fencei : enq_buffer_0_dec_uops_1_is_fencei; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4153 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_is_fencei : _GEN_4152; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4154 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_is_fencei : _GEN_4153; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4155 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_is_fencei : _GEN_4154; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4156 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_is_fencei : _GEN_4155; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4157 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_is_fencei : _GEN_4156; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4158 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_is_fencei : _GEN_4157; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4160 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_is_fence : enq_buffer_0_dec_uops_1_is_fence; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4161 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_is_fence : _GEN_4160; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4162 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_is_fence : _GEN_4161; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4163 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_is_fence : _GEN_4162; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4164 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_is_fence : _GEN_4163; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4165 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_is_fence : _GEN_4164; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4166 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_is_fence : _GEN_4165; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4168 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_mem_signed : enq_buffer_0_dec_uops_1_mem_signed; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4169 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_mem_signed : _GEN_4168; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4170 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_mem_signed : _GEN_4169; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4171 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_mem_signed : _GEN_4170; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4172 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_mem_signed : _GEN_4171; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4173 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_mem_signed : _GEN_4172; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4174 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_mem_signed : _GEN_4173; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4176 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_mem_size : enq_buffer_0_dec_uops_1_mem_size; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4177 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_mem_size : _GEN_4176; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4178 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_mem_size : _GEN_4177; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4179 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_mem_size : _GEN_4178; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4180 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_mem_size : _GEN_4179; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4181 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_mem_size : _GEN_4180; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4182 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_mem_size : _GEN_4181; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4184 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_mem_cmd : enq_buffer_0_dec_uops_1_mem_cmd; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4185 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_mem_cmd : _GEN_4184; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4186 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_mem_cmd : _GEN_4185; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4187 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_mem_cmd : _GEN_4186; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4188 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_mem_cmd : _GEN_4187; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4189 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_mem_cmd : _GEN_4188; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4190 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_mem_cmd : _GEN_4189; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4192 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_bypassable : enq_buffer_0_dec_uops_1_bypassable; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4193 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_bypassable : _GEN_4192; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4194 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_bypassable : _GEN_4193; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4195 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_bypassable : _GEN_4194; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4196 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_bypassable : _GEN_4195; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4197 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_bypassable : _GEN_4196; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4198 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_bypassable : _GEN_4197; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_4200 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_exc_cause : enq_buffer_0_dec_uops_1_exc_cause; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_4201 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_exc_cause : _GEN_4200; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_4202 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_exc_cause : _GEN_4201; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_4203 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_exc_cause : _GEN_4202; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_4204 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_exc_cause : _GEN_4203; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_4205 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_exc_cause : _GEN_4204; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_4206 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_exc_cause : _GEN_4205; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4208 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_exception : enq_buffer_0_dec_uops_1_exception; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4209 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_exception : _GEN_4208; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4210 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_exception : _GEN_4209; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4211 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_exception : _GEN_4210; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4212 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_exception : _GEN_4211; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4213 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_exception : _GEN_4212; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4214 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_exception : _GEN_4213; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4216 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_stale_pdst : enq_buffer_0_dec_uops_1_stale_pdst; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4217 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_stale_pdst : _GEN_4216; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4218 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_stale_pdst : _GEN_4217; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4219 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_stale_pdst : _GEN_4218; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4220 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_stale_pdst : _GEN_4219; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4221 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_stale_pdst : _GEN_4220; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4222 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_stale_pdst : _GEN_4221; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4224 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_ppred_busy : enq_buffer_0_dec_uops_1_ppred_busy; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4225 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_ppred_busy : _GEN_4224; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4226 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_ppred_busy : _GEN_4225; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4227 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_ppred_busy : _GEN_4226; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4228 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_ppred_busy : _GEN_4227; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4229 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_ppred_busy : _GEN_4228; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4230 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_ppred_busy : _GEN_4229; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4232 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_prs3_busy : enq_buffer_0_dec_uops_1_prs3_busy; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4233 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_prs3_busy : _GEN_4232; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4234 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_prs3_busy : _GEN_4233; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4235 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_prs3_busy : _GEN_4234; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4236 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_prs3_busy : _GEN_4235; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4237 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_prs3_busy : _GEN_4236; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4238 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_prs3_busy : _GEN_4237; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4240 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_prs2_busy : enq_buffer_0_dec_uops_1_prs2_busy; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4241 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_prs2_busy : _GEN_4240; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4242 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_prs2_busy : _GEN_4241; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4243 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_prs2_busy : _GEN_4242; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4244 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_prs2_busy : _GEN_4243; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4245 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_prs2_busy : _GEN_4244; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4246 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_prs2_busy : _GEN_4245; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4248 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_prs1_busy : enq_buffer_0_dec_uops_1_prs1_busy; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4249 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_prs1_busy : _GEN_4248; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4250 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_prs1_busy : _GEN_4249; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4251 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_prs1_busy : _GEN_4250; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4252 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_prs1_busy : _GEN_4251; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4253 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_prs1_busy : _GEN_4252; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4254 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_prs1_busy : _GEN_4253; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4256 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_ppred : enq_buffer_0_dec_uops_1_ppred; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4257 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_ppred : _GEN_4256; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4258 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_ppred : _GEN_4257; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4259 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_ppred : _GEN_4258; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4260 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_ppred : _GEN_4259; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4261 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_ppred : _GEN_4260; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4262 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_ppred : _GEN_4261; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4264 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_prs3 : enq_buffer_0_dec_uops_1_prs3; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4265 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_prs3 : _GEN_4264; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4266 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_prs3 : _GEN_4265; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4267 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_prs3 : _GEN_4266; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4268 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_prs3 : _GEN_4267; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4269 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_prs3 : _GEN_4268; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4270 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_prs3 : _GEN_4269; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4272 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_prs2 : enq_buffer_0_dec_uops_1_prs2; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4273 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_prs2 : _GEN_4272; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4274 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_prs2 : _GEN_4273; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4275 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_prs2 : _GEN_4274; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4276 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_prs2 : _GEN_4275; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4277 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_prs2 : _GEN_4276; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4278 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_prs2 : _GEN_4277; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4280 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_prs1 : enq_buffer_0_dec_uops_1_prs1; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4281 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_prs1 : _GEN_4280; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4282 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_prs1 : _GEN_4281; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4283 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_prs1 : _GEN_4282; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4284 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_prs1 : _GEN_4283; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4285 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_prs1 : _GEN_4284; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4286 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_prs1 : _GEN_4285; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4288 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_pdst : enq_buffer_0_dec_uops_1_pdst; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4289 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_pdst : _GEN_4288; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4290 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_pdst : _GEN_4289; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4291 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_pdst : _GEN_4290; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4292 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_pdst : _GEN_4291; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4293 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_pdst : _GEN_4292; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4294 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_pdst : _GEN_4293; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4296 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_rxq_idx : enq_buffer_0_dec_uops_1_rxq_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4297 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_rxq_idx : _GEN_4296; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4298 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_rxq_idx : _GEN_4297; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4299 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_rxq_idx : _GEN_4298; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4300 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_rxq_idx : _GEN_4299; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4301 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_rxq_idx : _GEN_4300; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4302 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_rxq_idx : _GEN_4301; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4304 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_stq_idx : enq_buffer_0_dec_uops_1_stq_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4305 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_stq_idx : _GEN_4304; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4306 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_stq_idx : _GEN_4305; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4307 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_stq_idx : _GEN_4306; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4308 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_stq_idx : _GEN_4307; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4309 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_stq_idx : _GEN_4308; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4310 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_stq_idx : _GEN_4309; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4312 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_ldq_idx : enq_buffer_0_dec_uops_1_ldq_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4313 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_ldq_idx : _GEN_4312; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4314 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_ldq_idx : _GEN_4313; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4315 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_ldq_idx : _GEN_4314; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4316 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_ldq_idx : _GEN_4315; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4317 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_ldq_idx : _GEN_4316; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4318 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_ldq_idx : _GEN_4317; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4320 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_rob_idx : enq_buffer_0_dec_uops_1_rob_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4321 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_rob_idx : _GEN_4320; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4322 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_rob_idx : _GEN_4321; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4323 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_rob_idx : _GEN_4322; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4324 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_rob_idx : _GEN_4323; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4325 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_rob_idx : _GEN_4324; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4326 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_rob_idx : _GEN_4325; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_4328 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_csr_addr : enq_buffer_0_dec_uops_1_csr_addr; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_4329 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_csr_addr : _GEN_4328; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_4330 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_csr_addr : _GEN_4329; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_4331 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_csr_addr : _GEN_4330; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_4332 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_csr_addr : _GEN_4331; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_4333 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_csr_addr : _GEN_4332; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_4334 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_csr_addr : _GEN_4333; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_4336 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_imm_packed : enq_buffer_0_dec_uops_1_imm_packed
    ; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_4337 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_imm_packed : _GEN_4336; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_4338 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_imm_packed : _GEN_4337; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_4339 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_imm_packed : _GEN_4338; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_4340 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_imm_packed : _GEN_4339; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_4341 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_imm_packed : _GEN_4340; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_4342 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_imm_packed : _GEN_4341; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4344 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_taken : enq_buffer_0_dec_uops_1_taken; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4345 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_taken : _GEN_4344; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4346 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_taken : _GEN_4345; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4347 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_taken : _GEN_4346; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4348 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_taken : _GEN_4347; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4349 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_taken : _GEN_4348; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4350 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_taken : _GEN_4349; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4352 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_pc_lob : enq_buffer_0_dec_uops_1_pc_lob; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4353 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_pc_lob : _GEN_4352; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4354 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_pc_lob : _GEN_4353; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4355 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_pc_lob : _GEN_4354; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4356 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_pc_lob : _GEN_4355; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4357 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_pc_lob : _GEN_4356; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4358 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_pc_lob : _GEN_4357; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4360 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_edge_inst : enq_buffer_0_dec_uops_1_edge_inst; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4361 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_edge_inst : _GEN_4360; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4362 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_edge_inst : _GEN_4361; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4363 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_edge_inst : _GEN_4362; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4364 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_edge_inst : _GEN_4363; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4365 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_edge_inst : _GEN_4364; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4366 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_edge_inst : _GEN_4365; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4368 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_ftq_idx : enq_buffer_0_dec_uops_1_ftq_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4369 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_ftq_idx : _GEN_4368; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4370 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_ftq_idx : _GEN_4369; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4371 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_ftq_idx : _GEN_4370; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4372 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_ftq_idx : _GEN_4371; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4373 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_ftq_idx : _GEN_4372; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4374 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_ftq_idx : _GEN_4373; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4376 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_br_tag : enq_buffer_0_dec_uops_1_br_tag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4377 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_br_tag : _GEN_4376; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4378 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_br_tag : _GEN_4377; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4379 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_br_tag : _GEN_4378; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4380 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_br_tag : _GEN_4379; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4381 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_br_tag : _GEN_4380; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4382 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_br_tag : _GEN_4381; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_4384 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_br_mask : enq_buffer_0_dec_uops_1_br_mask; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_4385 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_br_mask : _GEN_4384; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_4386 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_br_mask : _GEN_4385; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_4387 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_br_mask : _GEN_4386; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_4388 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_br_mask : _GEN_4387; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_4389 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_br_mask : _GEN_4388; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_4390 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_br_mask : _GEN_4389; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4392 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_is_sfb : enq_buffer_0_dec_uops_1_is_sfb; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4393 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_is_sfb : _GEN_4392; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4394 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_is_sfb : _GEN_4393; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4395 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_is_sfb : _GEN_4394; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4396 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_is_sfb : _GEN_4395; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4397 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_is_sfb : _GEN_4396; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4398 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_is_sfb : _GEN_4397; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4400 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_is_jal : enq_buffer_0_dec_uops_1_is_jal; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4401 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_is_jal : _GEN_4400; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4402 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_is_jal : _GEN_4401; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4403 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_is_jal : _GEN_4402; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4404 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_is_jal : _GEN_4403; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4405 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_is_jal : _GEN_4404; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4406 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_is_jal : _GEN_4405; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4408 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_is_jalr : enq_buffer_0_dec_uops_1_is_jalr; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4409 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_is_jalr : _GEN_4408; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4410 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_is_jalr : _GEN_4409; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4411 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_is_jalr : _GEN_4410; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4412 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_is_jalr : _GEN_4411; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4413 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_is_jalr : _GEN_4412; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4414 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_is_jalr : _GEN_4413; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4416 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_is_br : enq_buffer_0_dec_uops_1_is_br; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4417 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_is_br : _GEN_4416; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4418 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_is_br : _GEN_4417; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4419 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_is_br : _GEN_4418; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4420 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_is_br : _GEN_4419; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4421 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_is_br : _GEN_4420; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4422 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_is_br : _GEN_4421; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4424 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_iw_p2_poisoned :
    enq_buffer_0_dec_uops_1_iw_p2_poisoned; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4425 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_iw_p2_poisoned : _GEN_4424; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4426 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_iw_p2_poisoned : _GEN_4425; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4427 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_iw_p2_poisoned : _GEN_4426; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4428 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_iw_p2_poisoned : _GEN_4427; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4429 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_iw_p2_poisoned : _GEN_4428; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4430 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_iw_p2_poisoned : _GEN_4429; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4432 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_iw_p1_poisoned :
    enq_buffer_0_dec_uops_1_iw_p1_poisoned; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4433 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_iw_p1_poisoned : _GEN_4432; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4434 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_iw_p1_poisoned : _GEN_4433; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4435 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_iw_p1_poisoned : _GEN_4434; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4436 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_iw_p1_poisoned : _GEN_4435; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4437 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_iw_p1_poisoned : _GEN_4436; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4438 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_iw_p1_poisoned : _GEN_4437; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4440 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_iw_state : enq_buffer_0_dec_uops_1_iw_state; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4441 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_iw_state : _GEN_4440; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4442 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_iw_state : _GEN_4441; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4443 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_iw_state : _GEN_4442; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4444 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_iw_state : _GEN_4443; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4445 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_iw_state : _GEN_4444; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4446 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_iw_state : _GEN_4445; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4448 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_ctrl_op3_sel :
    enq_buffer_0_dec_uops_1_ctrl_op3_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4449 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_ctrl_op3_sel : _GEN_4448; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4450 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_ctrl_op3_sel : _GEN_4449; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4451 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_ctrl_op3_sel : _GEN_4450; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4452 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_ctrl_op3_sel : _GEN_4451; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4453 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_ctrl_op3_sel : _GEN_4452; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4454 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_ctrl_op3_sel : _GEN_4453; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4456 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_ctrl_is_std : enq_buffer_0_dec_uops_1_ctrl_is_std; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4457 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_ctrl_is_std : _GEN_4456; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4458 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_ctrl_is_std : _GEN_4457; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4459 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_ctrl_is_std : _GEN_4458; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4460 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_ctrl_is_std : _GEN_4459; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4461 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_ctrl_is_std : _GEN_4460; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4462 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_ctrl_is_std : _GEN_4461; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4464 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_ctrl_is_sta : enq_buffer_0_dec_uops_1_ctrl_is_sta; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4465 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_ctrl_is_sta : _GEN_4464; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4466 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_ctrl_is_sta : _GEN_4465; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4467 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_ctrl_is_sta : _GEN_4466; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4468 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_ctrl_is_sta : _GEN_4467; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4469 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_ctrl_is_sta : _GEN_4468; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4470 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_ctrl_is_sta : _GEN_4469; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4472 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_ctrl_is_load : enq_buffer_0_dec_uops_1_ctrl_is_load; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4473 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_ctrl_is_load : _GEN_4472; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4474 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_ctrl_is_load : _GEN_4473; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4475 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_ctrl_is_load : _GEN_4474; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4476 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_ctrl_is_load : _GEN_4475; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4477 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_ctrl_is_load : _GEN_4476; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4478 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_ctrl_is_load : _GEN_4477; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4480 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_ctrl_csr_cmd :
    enq_buffer_0_dec_uops_1_ctrl_csr_cmd; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4481 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_ctrl_csr_cmd : _GEN_4480; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4482 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_ctrl_csr_cmd : _GEN_4481; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4483 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_ctrl_csr_cmd : _GEN_4482; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4484 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_ctrl_csr_cmd : _GEN_4483; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4485 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_ctrl_csr_cmd : _GEN_4484; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4486 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_ctrl_csr_cmd : _GEN_4485; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4488 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_ctrl_fcn_dw : enq_buffer_0_dec_uops_1_ctrl_fcn_dw; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4489 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_ctrl_fcn_dw : _GEN_4488; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4490 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_ctrl_fcn_dw : _GEN_4489; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4491 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_ctrl_fcn_dw : _GEN_4490; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4492 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_ctrl_fcn_dw : _GEN_4491; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4493 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_ctrl_fcn_dw : _GEN_4492; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4494 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_ctrl_fcn_dw : _GEN_4493; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4496 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_ctrl_op_fcn :
    enq_buffer_0_dec_uops_1_ctrl_op_fcn; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4497 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_ctrl_op_fcn : _GEN_4496; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4498 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_ctrl_op_fcn : _GEN_4497; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4499 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_ctrl_op_fcn : _GEN_4498; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4500 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_ctrl_op_fcn : _GEN_4499; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4501 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_ctrl_op_fcn : _GEN_4500; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4502 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_ctrl_op_fcn : _GEN_4501; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4504 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_ctrl_imm_sel :
    enq_buffer_0_dec_uops_1_ctrl_imm_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4505 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_ctrl_imm_sel : _GEN_4504; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4506 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_ctrl_imm_sel : _GEN_4505; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4507 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_ctrl_imm_sel : _GEN_4506; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4508 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_ctrl_imm_sel : _GEN_4507; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4509 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_ctrl_imm_sel : _GEN_4508; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4510 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_ctrl_imm_sel : _GEN_4509; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4512 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_ctrl_op2_sel :
    enq_buffer_0_dec_uops_1_ctrl_op2_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4513 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_ctrl_op2_sel : _GEN_4512; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4514 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_ctrl_op2_sel : _GEN_4513; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4515 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_ctrl_op2_sel : _GEN_4514; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4516 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_ctrl_op2_sel : _GEN_4515; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4517 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_ctrl_op2_sel : _GEN_4516; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4518 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_ctrl_op2_sel : _GEN_4517; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4520 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_ctrl_op1_sel :
    enq_buffer_0_dec_uops_1_ctrl_op1_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4521 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_ctrl_op1_sel : _GEN_4520; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4522 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_ctrl_op1_sel : _GEN_4521; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4523 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_ctrl_op1_sel : _GEN_4522; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4524 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_ctrl_op1_sel : _GEN_4523; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4525 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_ctrl_op1_sel : _GEN_4524; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4526 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_ctrl_op1_sel : _GEN_4525; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4528 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_ctrl_br_type :
    enq_buffer_0_dec_uops_1_ctrl_br_type; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4529 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_ctrl_br_type : _GEN_4528; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4530 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_ctrl_br_type : _GEN_4529; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4531 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_ctrl_br_type : _GEN_4530; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4532 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_ctrl_br_type : _GEN_4531; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4533 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_ctrl_br_type : _GEN_4532; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4534 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_ctrl_br_type : _GEN_4533; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_4536 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_fu_code : enq_buffer_0_dec_uops_1_fu_code; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_4537 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_fu_code : _GEN_4536; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_4538 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_fu_code : _GEN_4537; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_4539 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_fu_code : _GEN_4538; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_4540 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_fu_code : _GEN_4539; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_4541 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_fu_code : _GEN_4540; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_4542 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_fu_code : _GEN_4541; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4544 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_iq_type : enq_buffer_0_dec_uops_1_iq_type; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4545 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_iq_type : _GEN_4544; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4546 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_iq_type : _GEN_4545; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4547 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_iq_type : _GEN_4546; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4548 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_iq_type : _GEN_4547; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4549 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_iq_type : _GEN_4548; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4550 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_iq_type : _GEN_4549; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_4552 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_debug_pc : enq_buffer_0_dec_uops_1_debug_pc; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_4553 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_debug_pc : _GEN_4552; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_4554 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_debug_pc : _GEN_4553; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_4555 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_debug_pc : _GEN_4554; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_4556 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_debug_pc : _GEN_4555; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_4557 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_debug_pc : _GEN_4556; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_4558 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_debug_pc : _GEN_4557; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4560 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_is_rvc : enq_buffer_0_dec_uops_1_is_rvc; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4561 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_is_rvc : _GEN_4560; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4562 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_is_rvc : _GEN_4561; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4563 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_is_rvc : _GEN_4562; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4564 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_is_rvc : _GEN_4563; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4565 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_is_rvc : _GEN_4564; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4566 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_is_rvc : _GEN_4565; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_4568 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_debug_inst : enq_buffer_0_dec_uops_1_debug_inst
    ; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_4569 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_debug_inst : _GEN_4568; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_4570 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_debug_inst : _GEN_4569; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_4571 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_debug_inst : _GEN_4570; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_4572 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_debug_inst : _GEN_4571; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_4573 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_debug_inst : _GEN_4572; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_4574 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_debug_inst : _GEN_4573; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_4576 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_inst : enq_buffer_0_dec_uops_1_inst; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_4577 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_inst : _GEN_4576; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_4578 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_inst : _GEN_4577; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_4579 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_inst : _GEN_4578; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_4580 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_inst : _GEN_4579; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_4581 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_inst : _GEN_4580; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_4582 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_inst : _GEN_4581; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4584 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_uopc : enq_buffer_0_dec_uops_1_uopc; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4585 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_uopc : _GEN_4584; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4586 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_uopc : _GEN_4585; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4587 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_uopc : _GEN_4586; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4588 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_uopc : _GEN_4587; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4589 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_uopc : _GEN_4588; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4590 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_uopc : _GEN_4589; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4592 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_address_num :
    enq_buffer_0_dec_uops_1_address_num; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4593 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_address_num : _GEN_4592; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4594 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_address_num : _GEN_4593; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4595 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_address_num : _GEN_4594; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4596 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_address_num : _GEN_4595; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4597 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_address_num : _GEN_4596; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4598 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_address_num : _GEN_4597; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4600 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_rob_inst_idx :
    enq_buffer_0_dec_uops_1_rob_inst_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4601 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_rob_inst_idx : _GEN_4600; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4602 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_rob_inst_idx : _GEN_4601; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4603 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_rob_inst_idx : _GEN_4602; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4604 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_rob_inst_idx : _GEN_4603; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4605 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_rob_inst_idx : _GEN_4604; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4606 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_rob_inst_idx : _GEN_4605; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4608 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_self_index : enq_buffer_0_dec_uops_1_self_index; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4609 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_self_index : _GEN_4608; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4610 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_self_index : _GEN_4609; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4611 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_self_index : _GEN_4610; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4612 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_self_index : _GEN_4611; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4613 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_self_index : _GEN_4612; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4614 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_self_index : _GEN_4613; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4616 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_split_num : enq_buffer_0_dec_uops_1_split_num; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4617 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_split_num : _GEN_4616; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4618 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_split_num : _GEN_4617; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4619 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_split_num : _GEN_4618; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4620 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_split_num : _GEN_4619; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4621 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_split_num : _GEN_4620; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4622 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_split_num : _GEN_4621; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4624 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_op2_sel : enq_buffer_0_dec_uops_1_op2_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4625 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_op2_sel : _GEN_4624; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4626 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_op2_sel : _GEN_4625; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4627 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_op2_sel : _GEN_4626; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4628 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_op2_sel : _GEN_4627; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4629 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_op2_sel : _GEN_4628; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4630 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_op2_sel : _GEN_4629; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4632 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_op1_sel : enq_buffer_0_dec_uops_1_op1_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4633 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_op1_sel : _GEN_4632; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4634 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_op1_sel : _GEN_4633; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4635 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_op1_sel : _GEN_4634; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4636 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_op1_sel : _GEN_4635; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4637 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_op1_sel : _GEN_4636; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4638 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_op1_sel : _GEN_4637; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4640 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_stale_pflag :
    enq_buffer_0_dec_uops_1_stale_pflag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4641 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_stale_pflag : _GEN_4640; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4642 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_stale_pflag : _GEN_4641; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4643 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_stale_pflag : _GEN_4642; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4644 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_stale_pflag : _GEN_4643; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4645 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_stale_pflag : _GEN_4644; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4646 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_stale_pflag : _GEN_4645; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4648 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_pflag_busy : enq_buffer_0_dec_uops_1_pflag_busy; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4649 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_pflag_busy : _GEN_4648; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4650 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_pflag_busy : _GEN_4649; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4651 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_pflag_busy : _GEN_4650; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4652 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_pflag_busy : _GEN_4651; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4653 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_pflag_busy : _GEN_4652; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4654 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_pflag_busy : _GEN_4653; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4656 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_pwflag : enq_buffer_0_dec_uops_1_pwflag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4657 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_pwflag : _GEN_4656; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4658 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_pwflag : _GEN_4657; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4659 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_pwflag : _GEN_4658; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4660 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_pwflag : _GEN_4659; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4661 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_pwflag : _GEN_4660; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4662 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_pwflag : _GEN_4661; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4664 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_prflag : enq_buffer_0_dec_uops_1_prflag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4665 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_prflag : _GEN_4664; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4666 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_prflag : _GEN_4665; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4667 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_prflag : _GEN_4666; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4668 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_prflag : _GEN_4667; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4669 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_prflag : _GEN_4668; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_4670 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_prflag : _GEN_4669; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4672 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_wflag : enq_buffer_0_dec_uops_1_wflag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4673 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_wflag : _GEN_4672; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4674 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_wflag : _GEN_4673; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4675 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_wflag : _GEN_4674; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4676 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_wflag : _GEN_4675; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4677 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_wflag : _GEN_4676; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4678 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_wflag : _GEN_4677; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4680 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_rflag : enq_buffer_0_dec_uops_1_rflag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4681 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_rflag : _GEN_4680; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4682 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_rflag : _GEN_4681; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4683 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_rflag : _GEN_4682; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4684 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_rflag : _GEN_4683; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4685 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_rflag : _GEN_4684; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4686 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_rflag : _GEN_4685; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4688 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_lrs3_rtype : enq_buffer_0_dec_uops_1_lrs3_rtype; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4689 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_lrs3_rtype : _GEN_4688; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4690 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_lrs3_rtype : _GEN_4689; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4691 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_lrs3_rtype : _GEN_4690; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4692 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_lrs3_rtype : _GEN_4691; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4693 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_lrs3_rtype : _GEN_4692; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4694 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_lrs3_rtype : _GEN_4693; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4696 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_shift : enq_buffer_0_dec_uops_1_shift; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4697 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_shift : _GEN_4696; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4698 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_shift : _GEN_4697; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4699 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_shift : _GEN_4698; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4700 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_shift : _GEN_4699; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4701 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_shift : _GEN_4700; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_4702 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_shift : _GEN_4701; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4704 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_is_unicore : enq_buffer_0_dec_uops_1_is_unicore; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4705 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_is_unicore : _GEN_4704; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4706 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_is_unicore : _GEN_4705; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4707 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_is_unicore : _GEN_4706; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4708 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_is_unicore : _GEN_4707; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4709 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_is_unicore : _GEN_4708; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4710 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_is_unicore : _GEN_4709; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4712 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_switch_off : enq_buffer_0_dec_uops_1_switch_off; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4713 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_switch_off : _GEN_4712; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4714 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_switch_off : _GEN_4713; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4715 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_switch_off : _GEN_4714; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4716 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_switch_off : _GEN_4715; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4717 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_switch_off : _GEN_4716; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4718 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_switch_off : _GEN_4717; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4720 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_1_switch : enq_buffer_0_dec_uops_1_switch; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4721 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_1_switch : _GEN_4720; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4722 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_1_switch : _GEN_4721; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4723 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_1_switch : _GEN_4722; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4724 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_1_switch : _GEN_4723; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4725 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_1_switch : _GEN_4724; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4726 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_1_switch : _GEN_4725; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4728 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_debug_tsrc : enq_buffer_0_dec_uops_2_debug_tsrc; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4729 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_debug_tsrc : _GEN_4728; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4730 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_debug_tsrc : _GEN_4729; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4731 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_debug_tsrc : _GEN_4730; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4732 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_debug_tsrc : _GEN_4731; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4733 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_debug_tsrc : _GEN_4732; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4734 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_debug_tsrc : _GEN_4733; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4736 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_debug_fsrc : enq_buffer_0_dec_uops_2_debug_fsrc; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4737 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_debug_fsrc : _GEN_4736; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4738 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_debug_fsrc : _GEN_4737; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4739 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_debug_fsrc : _GEN_4738; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4740 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_debug_fsrc : _GEN_4739; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4741 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_debug_fsrc : _GEN_4740; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4742 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_debug_fsrc : _GEN_4741; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4744 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_bp_xcpt_if : enq_buffer_0_dec_uops_2_bp_xcpt_if; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4745 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_bp_xcpt_if : _GEN_4744; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4746 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_bp_xcpt_if : _GEN_4745; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4747 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_bp_xcpt_if : _GEN_4746; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4748 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_bp_xcpt_if : _GEN_4747; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4749 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_bp_xcpt_if : _GEN_4748; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4750 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_bp_xcpt_if : _GEN_4749; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4752 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_bp_debug_if : enq_buffer_0_dec_uops_2_bp_debug_if; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4753 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_bp_debug_if : _GEN_4752; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4754 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_bp_debug_if : _GEN_4753; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4755 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_bp_debug_if : _GEN_4754; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4756 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_bp_debug_if : _GEN_4755; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4757 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_bp_debug_if : _GEN_4756; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4758 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_bp_debug_if : _GEN_4757; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4760 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_xcpt_ma_if : enq_buffer_0_dec_uops_2_xcpt_ma_if; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4761 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_xcpt_ma_if : _GEN_4760; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4762 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_xcpt_ma_if : _GEN_4761; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4763 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_xcpt_ma_if : _GEN_4762; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4764 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_xcpt_ma_if : _GEN_4763; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4765 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_xcpt_ma_if : _GEN_4764; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4766 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_xcpt_ma_if : _GEN_4765; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4768 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_xcpt_ae_if : enq_buffer_0_dec_uops_2_xcpt_ae_if; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4769 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_xcpt_ae_if : _GEN_4768; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4770 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_xcpt_ae_if : _GEN_4769; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4771 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_xcpt_ae_if : _GEN_4770; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4772 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_xcpt_ae_if : _GEN_4771; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4773 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_xcpt_ae_if : _GEN_4772; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4774 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_xcpt_ae_if : _GEN_4773; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4776 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_xcpt_pf_if : enq_buffer_0_dec_uops_2_xcpt_pf_if; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4777 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_xcpt_pf_if : _GEN_4776; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4778 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_xcpt_pf_if : _GEN_4777; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4779 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_xcpt_pf_if : _GEN_4778; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4780 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_xcpt_pf_if : _GEN_4779; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4781 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_xcpt_pf_if : _GEN_4780; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4782 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_xcpt_pf_if : _GEN_4781; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4784 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_fp_single : enq_buffer_0_dec_uops_2_fp_single; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4785 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_fp_single : _GEN_4784; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4786 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_fp_single : _GEN_4785; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4787 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_fp_single : _GEN_4786; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4788 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_fp_single : _GEN_4787; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4789 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_fp_single : _GEN_4788; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4790 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_fp_single : _GEN_4789; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4792 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_fp_val : enq_buffer_0_dec_uops_2_fp_val; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4793 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_fp_val : _GEN_4792; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4794 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_fp_val : _GEN_4793; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4795 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_fp_val : _GEN_4794; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4796 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_fp_val : _GEN_4795; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4797 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_fp_val : _GEN_4796; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4798 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_fp_val : _GEN_4797; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4800 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_frs3_en : enq_buffer_0_dec_uops_2_frs3_en; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4801 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_frs3_en : _GEN_4800; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4802 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_frs3_en : _GEN_4801; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4803 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_frs3_en : _GEN_4802; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4804 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_frs3_en : _GEN_4803; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4805 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_frs3_en : _GEN_4804; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4806 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_frs3_en : _GEN_4805; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4808 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_lrs2_rtype : enq_buffer_0_dec_uops_2_lrs2_rtype; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4809 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_lrs2_rtype : _GEN_4808; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4810 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_lrs2_rtype : _GEN_4809; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4811 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_lrs2_rtype : _GEN_4810; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4812 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_lrs2_rtype : _GEN_4811; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4813 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_lrs2_rtype : _GEN_4812; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4814 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_lrs2_rtype : _GEN_4813; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4816 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_lrs1_rtype : enq_buffer_0_dec_uops_2_lrs1_rtype; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4817 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_lrs1_rtype : _GEN_4816; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4818 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_lrs1_rtype : _GEN_4817; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4819 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_lrs1_rtype : _GEN_4818; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4820 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_lrs1_rtype : _GEN_4819; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4821 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_lrs1_rtype : _GEN_4820; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4822 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_lrs1_rtype : _GEN_4821; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4824 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_dst_rtype : enq_buffer_0_dec_uops_2_dst_rtype; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4825 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_dst_rtype : _GEN_4824; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4826 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_dst_rtype : _GEN_4825; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4827 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_dst_rtype : _GEN_4826; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4828 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_dst_rtype : _GEN_4827; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4829 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_dst_rtype : _GEN_4828; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4830 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_dst_rtype : _GEN_4829; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4832 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_ldst_val : enq_buffer_0_dec_uops_2_ldst_val; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4833 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_ldst_val : _GEN_4832; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4834 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_ldst_val : _GEN_4833; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4835 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_ldst_val : _GEN_4834; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4836 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_ldst_val : _GEN_4835; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4837 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_ldst_val : _GEN_4836; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4838 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_ldst_val : _GEN_4837; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4840 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_lrs3 : enq_buffer_0_dec_uops_2_lrs3; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4841 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_lrs3 : _GEN_4840; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4842 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_lrs3 : _GEN_4841; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4843 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_lrs3 : _GEN_4842; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4844 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_lrs3 : _GEN_4843; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4845 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_lrs3 : _GEN_4844; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4846 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_lrs3 : _GEN_4845; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4848 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_lrs2 : enq_buffer_0_dec_uops_2_lrs2; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4849 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_lrs2 : _GEN_4848; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4850 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_lrs2 : _GEN_4849; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4851 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_lrs2 : _GEN_4850; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4852 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_lrs2 : _GEN_4851; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4853 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_lrs2 : _GEN_4852; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4854 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_lrs2 : _GEN_4853; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4856 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_lrs1 : enq_buffer_0_dec_uops_2_lrs1; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4857 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_lrs1 : _GEN_4856; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4858 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_lrs1 : _GEN_4857; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4859 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_lrs1 : _GEN_4858; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4860 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_lrs1 : _GEN_4859; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4861 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_lrs1 : _GEN_4860; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4862 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_lrs1 : _GEN_4861; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4864 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_ldst : enq_buffer_0_dec_uops_2_ldst; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4865 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_ldst : _GEN_4864; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4866 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_ldst : _GEN_4865; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4867 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_ldst : _GEN_4866; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4868 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_ldst : _GEN_4867; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4869 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_ldst : _GEN_4868; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_4870 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_ldst : _GEN_4869; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4872 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_ldst_is_rs1 : enq_buffer_0_dec_uops_2_ldst_is_rs1; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4873 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_ldst_is_rs1 : _GEN_4872; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4874 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_ldst_is_rs1 : _GEN_4873; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4875 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_ldst_is_rs1 : _GEN_4874; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4876 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_ldst_is_rs1 : _GEN_4875; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4877 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_ldst_is_rs1 : _GEN_4876; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4878 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_ldst_is_rs1 : _GEN_4877; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4880 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_flush_on_commit :
    enq_buffer_0_dec_uops_2_flush_on_commit; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4881 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_flush_on_commit : _GEN_4880; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4882 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_flush_on_commit : _GEN_4881; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4883 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_flush_on_commit : _GEN_4882; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4884 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_flush_on_commit : _GEN_4883; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4885 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_flush_on_commit : _GEN_4884; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4886 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_flush_on_commit : _GEN_4885; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4888 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_is_unique : enq_buffer_0_dec_uops_2_is_unique; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4889 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_is_unique : _GEN_4888; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4890 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_is_unique : _GEN_4889; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4891 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_is_unique : _GEN_4890; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4892 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_is_unique : _GEN_4891; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4893 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_is_unique : _GEN_4892; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4894 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_is_unique : _GEN_4893; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4896 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_is_sys_pc2epc : enq_buffer_0_dec_uops_2_is_sys_pc2epc
    ; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4897 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_is_sys_pc2epc : _GEN_4896; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4898 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_is_sys_pc2epc : _GEN_4897; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4899 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_is_sys_pc2epc : _GEN_4898; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4900 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_is_sys_pc2epc : _GEN_4899; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4901 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_is_sys_pc2epc : _GEN_4900; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4902 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_is_sys_pc2epc : _GEN_4901; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4904 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_uses_stq : enq_buffer_0_dec_uops_2_uses_stq; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4905 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_uses_stq : _GEN_4904; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4906 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_uses_stq : _GEN_4905; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4907 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_uses_stq : _GEN_4906; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4908 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_uses_stq : _GEN_4907; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4909 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_uses_stq : _GEN_4908; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4910 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_uses_stq : _GEN_4909; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4912 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_uses_ldq : enq_buffer_0_dec_uops_2_uses_ldq; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4913 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_uses_ldq : _GEN_4912; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4914 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_uses_ldq : _GEN_4913; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4915 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_uses_ldq : _GEN_4914; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4916 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_uses_ldq : _GEN_4915; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4917 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_uses_ldq : _GEN_4916; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4918 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_uses_ldq : _GEN_4917; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4920 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_is_amo : enq_buffer_0_dec_uops_2_is_amo; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4921 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_is_amo : _GEN_4920; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4922 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_is_amo : _GEN_4921; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4923 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_is_amo : _GEN_4922; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4924 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_is_amo : _GEN_4923; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4925 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_is_amo : _GEN_4924; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4926 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_is_amo : _GEN_4925; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4928 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_is_fencei : enq_buffer_0_dec_uops_2_is_fencei; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4929 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_is_fencei : _GEN_4928; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4930 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_is_fencei : _GEN_4929; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4931 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_is_fencei : _GEN_4930; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4932 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_is_fencei : _GEN_4931; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4933 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_is_fencei : _GEN_4932; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4934 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_is_fencei : _GEN_4933; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4936 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_is_fence : enq_buffer_0_dec_uops_2_is_fence; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4937 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_is_fence : _GEN_4936; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4938 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_is_fence : _GEN_4937; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4939 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_is_fence : _GEN_4938; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4940 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_is_fence : _GEN_4939; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4941 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_is_fence : _GEN_4940; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4942 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_is_fence : _GEN_4941; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4944 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_mem_signed : enq_buffer_0_dec_uops_2_mem_signed; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4945 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_mem_signed : _GEN_4944; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4946 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_mem_signed : _GEN_4945; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4947 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_mem_signed : _GEN_4946; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4948 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_mem_signed : _GEN_4947; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4949 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_mem_signed : _GEN_4948; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4950 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_mem_signed : _GEN_4949; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4952 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_mem_size : enq_buffer_0_dec_uops_2_mem_size; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4953 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_mem_size : _GEN_4952; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4954 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_mem_size : _GEN_4953; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4955 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_mem_size : _GEN_4954; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4956 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_mem_size : _GEN_4955; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4957 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_mem_size : _GEN_4956; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_4958 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_mem_size : _GEN_4957; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4960 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_mem_cmd : enq_buffer_0_dec_uops_2_mem_cmd; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4961 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_mem_cmd : _GEN_4960; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4962 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_mem_cmd : _GEN_4961; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4963 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_mem_cmd : _GEN_4962; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4964 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_mem_cmd : _GEN_4963; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4965 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_mem_cmd : _GEN_4964; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_4966 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_mem_cmd : _GEN_4965; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4968 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_bypassable : enq_buffer_0_dec_uops_2_bypassable; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4969 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_bypassable : _GEN_4968; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4970 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_bypassable : _GEN_4969; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4971 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_bypassable : _GEN_4970; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4972 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_bypassable : _GEN_4971; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4973 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_bypassable : _GEN_4972; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4974 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_bypassable : _GEN_4973; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_4976 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_exc_cause : enq_buffer_0_dec_uops_2_exc_cause; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_4977 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_exc_cause : _GEN_4976; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_4978 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_exc_cause : _GEN_4977; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_4979 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_exc_cause : _GEN_4978; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_4980 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_exc_cause : _GEN_4979; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_4981 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_exc_cause : _GEN_4980; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_4982 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_exc_cause : _GEN_4981; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4984 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_exception : enq_buffer_0_dec_uops_2_exception; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4985 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_exception : _GEN_4984; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4986 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_exception : _GEN_4985; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4987 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_exception : _GEN_4986; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4988 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_exception : _GEN_4987; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4989 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_exception : _GEN_4988; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_4990 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_exception : _GEN_4989; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4992 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_stale_pdst : enq_buffer_0_dec_uops_2_stale_pdst; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4993 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_stale_pdst : _GEN_4992; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4994 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_stale_pdst : _GEN_4993; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4995 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_stale_pdst : _GEN_4994; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4996 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_stale_pdst : _GEN_4995; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4997 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_stale_pdst : _GEN_4996; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_4998 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_stale_pdst : _GEN_4997; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5000 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_ppred_busy : enq_buffer_0_dec_uops_2_ppred_busy; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5001 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_ppred_busy : _GEN_5000; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5002 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_ppred_busy : _GEN_5001; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5003 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_ppred_busy : _GEN_5002; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5004 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_ppred_busy : _GEN_5003; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5005 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_ppred_busy : _GEN_5004; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5006 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_ppred_busy : _GEN_5005; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5008 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_prs3_busy : enq_buffer_0_dec_uops_2_prs3_busy; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5009 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_prs3_busy : _GEN_5008; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5010 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_prs3_busy : _GEN_5009; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5011 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_prs3_busy : _GEN_5010; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5012 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_prs3_busy : _GEN_5011; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5013 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_prs3_busy : _GEN_5012; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5014 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_prs3_busy : _GEN_5013; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5016 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_prs2_busy : enq_buffer_0_dec_uops_2_prs2_busy; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5017 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_prs2_busy : _GEN_5016; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5018 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_prs2_busy : _GEN_5017; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5019 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_prs2_busy : _GEN_5018; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5020 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_prs2_busy : _GEN_5019; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5021 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_prs2_busy : _GEN_5020; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5022 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_prs2_busy : _GEN_5021; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5024 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_prs1_busy : enq_buffer_0_dec_uops_2_prs1_busy; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5025 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_prs1_busy : _GEN_5024; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5026 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_prs1_busy : _GEN_5025; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5027 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_prs1_busy : _GEN_5026; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5028 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_prs1_busy : _GEN_5027; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5029 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_prs1_busy : _GEN_5028; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5030 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_prs1_busy : _GEN_5029; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5032 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_ppred : enq_buffer_0_dec_uops_2_ppred; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5033 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_ppred : _GEN_5032; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5034 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_ppred : _GEN_5033; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5035 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_ppred : _GEN_5034; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5036 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_ppred : _GEN_5035; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5037 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_ppred : _GEN_5036; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5038 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_ppred : _GEN_5037; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5040 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_prs3 : enq_buffer_0_dec_uops_2_prs3; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5041 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_prs3 : _GEN_5040; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5042 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_prs3 : _GEN_5041; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5043 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_prs3 : _GEN_5042; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5044 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_prs3 : _GEN_5043; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5045 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_prs3 : _GEN_5044; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5046 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_prs3 : _GEN_5045; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5048 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_prs2 : enq_buffer_0_dec_uops_2_prs2; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5049 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_prs2 : _GEN_5048; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5050 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_prs2 : _GEN_5049; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5051 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_prs2 : _GEN_5050; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5052 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_prs2 : _GEN_5051; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5053 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_prs2 : _GEN_5052; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5054 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_prs2 : _GEN_5053; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5056 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_prs1 : enq_buffer_0_dec_uops_2_prs1; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5057 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_prs1 : _GEN_5056; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5058 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_prs1 : _GEN_5057; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5059 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_prs1 : _GEN_5058; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5060 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_prs1 : _GEN_5059; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5061 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_prs1 : _GEN_5060; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5062 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_prs1 : _GEN_5061; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5064 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_pdst : enq_buffer_0_dec_uops_2_pdst; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5065 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_pdst : _GEN_5064; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5066 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_pdst : _GEN_5065; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5067 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_pdst : _GEN_5066; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5068 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_pdst : _GEN_5067; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5069 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_pdst : _GEN_5068; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5070 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_pdst : _GEN_5069; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5072 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_rxq_idx : enq_buffer_0_dec_uops_2_rxq_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5073 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_rxq_idx : _GEN_5072; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5074 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_rxq_idx : _GEN_5073; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5075 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_rxq_idx : _GEN_5074; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5076 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_rxq_idx : _GEN_5075; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5077 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_rxq_idx : _GEN_5076; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5078 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_rxq_idx : _GEN_5077; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5080 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_stq_idx : enq_buffer_0_dec_uops_2_stq_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5081 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_stq_idx : _GEN_5080; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5082 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_stq_idx : _GEN_5081; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5083 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_stq_idx : _GEN_5082; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5084 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_stq_idx : _GEN_5083; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5085 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_stq_idx : _GEN_5084; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5086 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_stq_idx : _GEN_5085; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5088 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_ldq_idx : enq_buffer_0_dec_uops_2_ldq_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5089 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_ldq_idx : _GEN_5088; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5090 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_ldq_idx : _GEN_5089; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5091 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_ldq_idx : _GEN_5090; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5092 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_ldq_idx : _GEN_5091; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5093 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_ldq_idx : _GEN_5092; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5094 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_ldq_idx : _GEN_5093; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5096 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_rob_idx : enq_buffer_0_dec_uops_2_rob_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5097 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_rob_idx : _GEN_5096; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5098 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_rob_idx : _GEN_5097; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5099 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_rob_idx : _GEN_5098; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5100 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_rob_idx : _GEN_5099; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5101 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_rob_idx : _GEN_5100; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5102 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_rob_idx : _GEN_5101; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5104 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_csr_addr : enq_buffer_0_dec_uops_2_csr_addr; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5105 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_csr_addr : _GEN_5104; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5106 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_csr_addr : _GEN_5105; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5107 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_csr_addr : _GEN_5106; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5108 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_csr_addr : _GEN_5107; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5109 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_csr_addr : _GEN_5108; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5110 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_csr_addr : _GEN_5109; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_5112 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_imm_packed : enq_buffer_0_dec_uops_2_imm_packed
    ; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_5113 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_imm_packed : _GEN_5112; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_5114 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_imm_packed : _GEN_5113; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_5115 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_imm_packed : _GEN_5114; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_5116 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_imm_packed : _GEN_5115; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_5117 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_imm_packed : _GEN_5116; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_5118 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_imm_packed : _GEN_5117; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5120 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_taken : enq_buffer_0_dec_uops_2_taken; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5121 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_taken : _GEN_5120; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5122 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_taken : _GEN_5121; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5123 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_taken : _GEN_5122; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5124 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_taken : _GEN_5123; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5125 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_taken : _GEN_5124; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5126 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_taken : _GEN_5125; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5128 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_pc_lob : enq_buffer_0_dec_uops_2_pc_lob; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5129 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_pc_lob : _GEN_5128; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5130 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_pc_lob : _GEN_5129; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5131 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_pc_lob : _GEN_5130; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5132 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_pc_lob : _GEN_5131; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5133 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_pc_lob : _GEN_5132; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5134 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_pc_lob : _GEN_5133; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5136 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_edge_inst : enq_buffer_0_dec_uops_2_edge_inst; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5137 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_edge_inst : _GEN_5136; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5138 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_edge_inst : _GEN_5137; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5139 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_edge_inst : _GEN_5138; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5140 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_edge_inst : _GEN_5139; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5141 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_edge_inst : _GEN_5140; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5142 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_edge_inst : _GEN_5141; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5144 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_ftq_idx : enq_buffer_0_dec_uops_2_ftq_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5145 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_ftq_idx : _GEN_5144; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5146 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_ftq_idx : _GEN_5145; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5147 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_ftq_idx : _GEN_5146; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5148 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_ftq_idx : _GEN_5147; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5149 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_ftq_idx : _GEN_5148; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5150 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_ftq_idx : _GEN_5149; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5152 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_br_tag : enq_buffer_0_dec_uops_2_br_tag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5153 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_br_tag : _GEN_5152; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5154 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_br_tag : _GEN_5153; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5155 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_br_tag : _GEN_5154; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5156 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_br_tag : _GEN_5155; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5157 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_br_tag : _GEN_5156; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5158 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_br_tag : _GEN_5157; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5160 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_br_mask : enq_buffer_0_dec_uops_2_br_mask; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5161 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_br_mask : _GEN_5160; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5162 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_br_mask : _GEN_5161; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5163 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_br_mask : _GEN_5162; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5164 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_br_mask : _GEN_5163; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5165 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_br_mask : _GEN_5164; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5166 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_br_mask : _GEN_5165; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5168 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_is_sfb : enq_buffer_0_dec_uops_2_is_sfb; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5169 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_is_sfb : _GEN_5168; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5170 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_is_sfb : _GEN_5169; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5171 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_is_sfb : _GEN_5170; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5172 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_is_sfb : _GEN_5171; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5173 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_is_sfb : _GEN_5172; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5174 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_is_sfb : _GEN_5173; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5176 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_is_jal : enq_buffer_0_dec_uops_2_is_jal; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5177 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_is_jal : _GEN_5176; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5178 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_is_jal : _GEN_5177; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5179 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_is_jal : _GEN_5178; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5180 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_is_jal : _GEN_5179; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5181 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_is_jal : _GEN_5180; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5182 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_is_jal : _GEN_5181; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5184 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_is_jalr : enq_buffer_0_dec_uops_2_is_jalr; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5185 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_is_jalr : _GEN_5184; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5186 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_is_jalr : _GEN_5185; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5187 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_is_jalr : _GEN_5186; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5188 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_is_jalr : _GEN_5187; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5189 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_is_jalr : _GEN_5188; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5190 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_is_jalr : _GEN_5189; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5192 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_is_br : enq_buffer_0_dec_uops_2_is_br; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5193 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_is_br : _GEN_5192; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5194 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_is_br : _GEN_5193; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5195 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_is_br : _GEN_5194; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5196 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_is_br : _GEN_5195; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5197 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_is_br : _GEN_5196; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5198 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_is_br : _GEN_5197; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5200 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_iw_p2_poisoned :
    enq_buffer_0_dec_uops_2_iw_p2_poisoned; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5201 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_iw_p2_poisoned : _GEN_5200; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5202 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_iw_p2_poisoned : _GEN_5201; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5203 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_iw_p2_poisoned : _GEN_5202; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5204 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_iw_p2_poisoned : _GEN_5203; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5205 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_iw_p2_poisoned : _GEN_5204; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5206 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_iw_p2_poisoned : _GEN_5205; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5208 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_iw_p1_poisoned :
    enq_buffer_0_dec_uops_2_iw_p1_poisoned; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5209 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_iw_p1_poisoned : _GEN_5208; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5210 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_iw_p1_poisoned : _GEN_5209; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5211 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_iw_p1_poisoned : _GEN_5210; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5212 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_iw_p1_poisoned : _GEN_5211; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5213 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_iw_p1_poisoned : _GEN_5212; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5214 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_iw_p1_poisoned : _GEN_5213; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5216 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_iw_state : enq_buffer_0_dec_uops_2_iw_state; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5217 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_iw_state : _GEN_5216; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5218 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_iw_state : _GEN_5217; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5219 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_iw_state : _GEN_5218; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5220 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_iw_state : _GEN_5219; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5221 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_iw_state : _GEN_5220; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5222 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_iw_state : _GEN_5221; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5224 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_ctrl_op3_sel :
    enq_buffer_0_dec_uops_2_ctrl_op3_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5225 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_ctrl_op3_sel : _GEN_5224; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5226 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_ctrl_op3_sel : _GEN_5225; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5227 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_ctrl_op3_sel : _GEN_5226; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5228 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_ctrl_op3_sel : _GEN_5227; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5229 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_ctrl_op3_sel : _GEN_5228; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5230 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_ctrl_op3_sel : _GEN_5229; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5232 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_ctrl_is_std : enq_buffer_0_dec_uops_2_ctrl_is_std; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5233 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_ctrl_is_std : _GEN_5232; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5234 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_ctrl_is_std : _GEN_5233; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5235 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_ctrl_is_std : _GEN_5234; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5236 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_ctrl_is_std : _GEN_5235; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5237 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_ctrl_is_std : _GEN_5236; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5238 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_ctrl_is_std : _GEN_5237; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5240 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_ctrl_is_sta : enq_buffer_0_dec_uops_2_ctrl_is_sta; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5241 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_ctrl_is_sta : _GEN_5240; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5242 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_ctrl_is_sta : _GEN_5241; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5243 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_ctrl_is_sta : _GEN_5242; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5244 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_ctrl_is_sta : _GEN_5243; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5245 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_ctrl_is_sta : _GEN_5244; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5246 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_ctrl_is_sta : _GEN_5245; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5248 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_ctrl_is_load : enq_buffer_0_dec_uops_2_ctrl_is_load; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5249 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_ctrl_is_load : _GEN_5248; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5250 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_ctrl_is_load : _GEN_5249; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5251 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_ctrl_is_load : _GEN_5250; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5252 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_ctrl_is_load : _GEN_5251; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5253 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_ctrl_is_load : _GEN_5252; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5254 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_ctrl_is_load : _GEN_5253; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5256 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_ctrl_csr_cmd :
    enq_buffer_0_dec_uops_2_ctrl_csr_cmd; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5257 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_ctrl_csr_cmd : _GEN_5256; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5258 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_ctrl_csr_cmd : _GEN_5257; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5259 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_ctrl_csr_cmd : _GEN_5258; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5260 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_ctrl_csr_cmd : _GEN_5259; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5261 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_ctrl_csr_cmd : _GEN_5260; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5262 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_ctrl_csr_cmd : _GEN_5261; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5264 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_ctrl_fcn_dw : enq_buffer_0_dec_uops_2_ctrl_fcn_dw; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5265 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_ctrl_fcn_dw : _GEN_5264; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5266 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_ctrl_fcn_dw : _GEN_5265; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5267 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_ctrl_fcn_dw : _GEN_5266; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5268 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_ctrl_fcn_dw : _GEN_5267; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5269 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_ctrl_fcn_dw : _GEN_5268; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5270 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_ctrl_fcn_dw : _GEN_5269; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5272 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_ctrl_op_fcn :
    enq_buffer_0_dec_uops_2_ctrl_op_fcn; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5273 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_ctrl_op_fcn : _GEN_5272; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5274 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_ctrl_op_fcn : _GEN_5273; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5275 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_ctrl_op_fcn : _GEN_5274; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5276 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_ctrl_op_fcn : _GEN_5275; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5277 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_ctrl_op_fcn : _GEN_5276; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5278 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_ctrl_op_fcn : _GEN_5277; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5280 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_ctrl_imm_sel :
    enq_buffer_0_dec_uops_2_ctrl_imm_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5281 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_ctrl_imm_sel : _GEN_5280; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5282 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_ctrl_imm_sel : _GEN_5281; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5283 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_ctrl_imm_sel : _GEN_5282; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5284 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_ctrl_imm_sel : _GEN_5283; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5285 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_ctrl_imm_sel : _GEN_5284; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5286 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_ctrl_imm_sel : _GEN_5285; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5288 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_ctrl_op2_sel :
    enq_buffer_0_dec_uops_2_ctrl_op2_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5289 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_ctrl_op2_sel : _GEN_5288; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5290 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_ctrl_op2_sel : _GEN_5289; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5291 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_ctrl_op2_sel : _GEN_5290; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5292 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_ctrl_op2_sel : _GEN_5291; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5293 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_ctrl_op2_sel : _GEN_5292; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5294 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_ctrl_op2_sel : _GEN_5293; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5296 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_ctrl_op1_sel :
    enq_buffer_0_dec_uops_2_ctrl_op1_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5297 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_ctrl_op1_sel : _GEN_5296; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5298 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_ctrl_op1_sel : _GEN_5297; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5299 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_ctrl_op1_sel : _GEN_5298; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5300 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_ctrl_op1_sel : _GEN_5299; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5301 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_ctrl_op1_sel : _GEN_5300; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5302 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_ctrl_op1_sel : _GEN_5301; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5304 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_ctrl_br_type :
    enq_buffer_0_dec_uops_2_ctrl_br_type; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5305 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_ctrl_br_type : _GEN_5304; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5306 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_ctrl_br_type : _GEN_5305; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5307 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_ctrl_br_type : _GEN_5306; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5308 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_ctrl_br_type : _GEN_5307; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5309 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_ctrl_br_type : _GEN_5308; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5310 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_ctrl_br_type : _GEN_5309; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_5312 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_fu_code : enq_buffer_0_dec_uops_2_fu_code; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_5313 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_fu_code : _GEN_5312; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_5314 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_fu_code : _GEN_5313; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_5315 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_fu_code : _GEN_5314; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_5316 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_fu_code : _GEN_5315; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_5317 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_fu_code : _GEN_5316; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_5318 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_fu_code : _GEN_5317; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5320 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_iq_type : enq_buffer_0_dec_uops_2_iq_type; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5321 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_iq_type : _GEN_5320; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5322 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_iq_type : _GEN_5321; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5323 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_iq_type : _GEN_5322; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5324 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_iq_type : _GEN_5323; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5325 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_iq_type : _GEN_5324; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5326 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_iq_type : _GEN_5325; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_5328 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_debug_pc : enq_buffer_0_dec_uops_2_debug_pc; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_5329 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_debug_pc : _GEN_5328; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_5330 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_debug_pc : _GEN_5329; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_5331 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_debug_pc : _GEN_5330; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_5332 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_debug_pc : _GEN_5331; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_5333 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_debug_pc : _GEN_5332; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_5334 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_debug_pc : _GEN_5333; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5336 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_is_rvc : enq_buffer_0_dec_uops_2_is_rvc; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5337 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_is_rvc : _GEN_5336; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5338 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_is_rvc : _GEN_5337; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5339 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_is_rvc : _GEN_5338; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5340 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_is_rvc : _GEN_5339; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5341 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_is_rvc : _GEN_5340; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5342 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_is_rvc : _GEN_5341; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_5344 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_debug_inst : enq_buffer_0_dec_uops_2_debug_inst
    ; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_5345 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_debug_inst : _GEN_5344; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_5346 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_debug_inst : _GEN_5345; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_5347 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_debug_inst : _GEN_5346; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_5348 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_debug_inst : _GEN_5347; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_5349 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_debug_inst : _GEN_5348; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_5350 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_debug_inst : _GEN_5349; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_5352 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_inst : enq_buffer_0_dec_uops_2_inst; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_5353 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_inst : _GEN_5352; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_5354 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_inst : _GEN_5353; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_5355 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_inst : _GEN_5354; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_5356 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_inst : _GEN_5355; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_5357 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_inst : _GEN_5356; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_5358 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_inst : _GEN_5357; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5360 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_uopc : enq_buffer_0_dec_uops_2_uopc; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5361 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_uopc : _GEN_5360; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5362 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_uopc : _GEN_5361; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5363 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_uopc : _GEN_5362; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5364 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_uopc : _GEN_5363; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5365 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_uopc : _GEN_5364; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5366 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_uopc : _GEN_5365; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5368 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_address_num :
    enq_buffer_0_dec_uops_2_address_num; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5369 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_address_num : _GEN_5368; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5370 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_address_num : _GEN_5369; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5371 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_address_num : _GEN_5370; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5372 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_address_num : _GEN_5371; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5373 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_address_num : _GEN_5372; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5374 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_address_num : _GEN_5373; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5376 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_rob_inst_idx :
    enq_buffer_0_dec_uops_2_rob_inst_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5377 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_rob_inst_idx : _GEN_5376; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5378 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_rob_inst_idx : _GEN_5377; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5379 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_rob_inst_idx : _GEN_5378; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5380 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_rob_inst_idx : _GEN_5379; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5381 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_rob_inst_idx : _GEN_5380; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5382 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_rob_inst_idx : _GEN_5381; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5384 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_self_index : enq_buffer_0_dec_uops_2_self_index; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5385 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_self_index : _GEN_5384; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5386 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_self_index : _GEN_5385; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5387 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_self_index : _GEN_5386; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5388 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_self_index : _GEN_5387; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5389 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_self_index : _GEN_5388; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5390 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_self_index : _GEN_5389; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5392 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_split_num : enq_buffer_0_dec_uops_2_split_num; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5393 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_split_num : _GEN_5392; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5394 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_split_num : _GEN_5393; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5395 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_split_num : _GEN_5394; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5396 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_split_num : _GEN_5395; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5397 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_split_num : _GEN_5396; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5398 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_split_num : _GEN_5397; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5400 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_op2_sel : enq_buffer_0_dec_uops_2_op2_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5401 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_op2_sel : _GEN_5400; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5402 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_op2_sel : _GEN_5401; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5403 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_op2_sel : _GEN_5402; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5404 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_op2_sel : _GEN_5403; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5405 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_op2_sel : _GEN_5404; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5406 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_op2_sel : _GEN_5405; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5408 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_op1_sel : enq_buffer_0_dec_uops_2_op1_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5409 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_op1_sel : _GEN_5408; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5410 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_op1_sel : _GEN_5409; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5411 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_op1_sel : _GEN_5410; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5412 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_op1_sel : _GEN_5411; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5413 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_op1_sel : _GEN_5412; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5414 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_op1_sel : _GEN_5413; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5416 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_stale_pflag :
    enq_buffer_0_dec_uops_2_stale_pflag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5417 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_stale_pflag : _GEN_5416; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5418 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_stale_pflag : _GEN_5417; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5419 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_stale_pflag : _GEN_5418; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5420 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_stale_pflag : _GEN_5419; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5421 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_stale_pflag : _GEN_5420; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5422 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_stale_pflag : _GEN_5421; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5424 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_pflag_busy : enq_buffer_0_dec_uops_2_pflag_busy; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5425 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_pflag_busy : _GEN_5424; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5426 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_pflag_busy : _GEN_5425; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5427 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_pflag_busy : _GEN_5426; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5428 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_pflag_busy : _GEN_5427; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5429 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_pflag_busy : _GEN_5428; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5430 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_pflag_busy : _GEN_5429; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5432 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_pwflag : enq_buffer_0_dec_uops_2_pwflag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5433 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_pwflag : _GEN_5432; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5434 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_pwflag : _GEN_5433; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5435 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_pwflag : _GEN_5434; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5436 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_pwflag : _GEN_5435; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5437 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_pwflag : _GEN_5436; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5438 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_pwflag : _GEN_5437; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5440 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_prflag : enq_buffer_0_dec_uops_2_prflag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5441 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_prflag : _GEN_5440; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5442 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_prflag : _GEN_5441; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5443 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_prflag : _GEN_5442; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5444 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_prflag : _GEN_5443; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5445 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_prflag : _GEN_5444; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5446 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_prflag : _GEN_5445; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5448 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_wflag : enq_buffer_0_dec_uops_2_wflag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5449 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_wflag : _GEN_5448; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5450 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_wflag : _GEN_5449; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5451 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_wflag : _GEN_5450; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5452 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_wflag : _GEN_5451; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5453 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_wflag : _GEN_5452; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5454 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_wflag : _GEN_5453; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5456 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_rflag : enq_buffer_0_dec_uops_2_rflag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5457 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_rflag : _GEN_5456; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5458 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_rflag : _GEN_5457; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5459 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_rflag : _GEN_5458; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5460 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_rflag : _GEN_5459; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5461 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_rflag : _GEN_5460; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5462 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_rflag : _GEN_5461; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5464 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_lrs3_rtype : enq_buffer_0_dec_uops_2_lrs3_rtype; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5465 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_lrs3_rtype : _GEN_5464; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5466 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_lrs3_rtype : _GEN_5465; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5467 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_lrs3_rtype : _GEN_5466; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5468 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_lrs3_rtype : _GEN_5467; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5469 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_lrs3_rtype : _GEN_5468; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5470 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_lrs3_rtype : _GEN_5469; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5472 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_shift : enq_buffer_0_dec_uops_2_shift; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5473 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_shift : _GEN_5472; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5474 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_shift : _GEN_5473; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5475 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_shift : _GEN_5474; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5476 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_shift : _GEN_5475; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5477 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_shift : _GEN_5476; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_5478 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_shift : _GEN_5477; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5480 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_is_unicore : enq_buffer_0_dec_uops_2_is_unicore; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5481 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_is_unicore : _GEN_5480; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5482 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_is_unicore : _GEN_5481; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5483 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_is_unicore : _GEN_5482; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5484 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_is_unicore : _GEN_5483; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5485 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_is_unicore : _GEN_5484; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5486 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_is_unicore : _GEN_5485; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5488 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_switch_off : enq_buffer_0_dec_uops_2_switch_off; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5489 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_switch_off : _GEN_5488; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5490 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_switch_off : _GEN_5489; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5491 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_switch_off : _GEN_5490; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5492 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_switch_off : _GEN_5491; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5493 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_switch_off : _GEN_5492; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5494 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_switch_off : _GEN_5493; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5496 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_2_switch : enq_buffer_0_dec_uops_2_switch; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5497 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_2_switch : _GEN_5496; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5498 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_2_switch : _GEN_5497; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5499 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_2_switch : _GEN_5498; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5500 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_2_switch : _GEN_5499; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5501 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_2_switch : _GEN_5500; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5502 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_2_switch : _GEN_5501; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5504 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_debug_tsrc : enq_buffer_0_dec_uops_3_debug_tsrc; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5505 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_debug_tsrc : _GEN_5504; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5506 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_debug_tsrc : _GEN_5505; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5507 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_debug_tsrc : _GEN_5506; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5508 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_debug_tsrc : _GEN_5507; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5509 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_debug_tsrc : _GEN_5508; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5510 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_debug_tsrc : _GEN_5509; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5512 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_debug_fsrc : enq_buffer_0_dec_uops_3_debug_fsrc; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5513 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_debug_fsrc : _GEN_5512; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5514 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_debug_fsrc : _GEN_5513; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5515 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_debug_fsrc : _GEN_5514; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5516 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_debug_fsrc : _GEN_5515; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5517 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_debug_fsrc : _GEN_5516; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5518 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_debug_fsrc : _GEN_5517; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5520 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_bp_xcpt_if : enq_buffer_0_dec_uops_3_bp_xcpt_if; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5521 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_bp_xcpt_if : _GEN_5520; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5522 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_bp_xcpt_if : _GEN_5521; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5523 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_bp_xcpt_if : _GEN_5522; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5524 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_bp_xcpt_if : _GEN_5523; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5525 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_bp_xcpt_if : _GEN_5524; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5526 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_bp_xcpt_if : _GEN_5525; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5528 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_bp_debug_if : enq_buffer_0_dec_uops_3_bp_debug_if; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5529 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_bp_debug_if : _GEN_5528; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5530 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_bp_debug_if : _GEN_5529; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5531 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_bp_debug_if : _GEN_5530; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5532 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_bp_debug_if : _GEN_5531; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5533 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_bp_debug_if : _GEN_5532; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5534 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_bp_debug_if : _GEN_5533; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5536 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_xcpt_ma_if : enq_buffer_0_dec_uops_3_xcpt_ma_if; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5537 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_xcpt_ma_if : _GEN_5536; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5538 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_xcpt_ma_if : _GEN_5537; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5539 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_xcpt_ma_if : _GEN_5538; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5540 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_xcpt_ma_if : _GEN_5539; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5541 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_xcpt_ma_if : _GEN_5540; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5542 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_xcpt_ma_if : _GEN_5541; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5544 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_xcpt_ae_if : enq_buffer_0_dec_uops_3_xcpt_ae_if; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5545 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_xcpt_ae_if : _GEN_5544; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5546 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_xcpt_ae_if : _GEN_5545; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5547 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_xcpt_ae_if : _GEN_5546; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5548 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_xcpt_ae_if : _GEN_5547; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5549 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_xcpt_ae_if : _GEN_5548; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5550 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_xcpt_ae_if : _GEN_5549; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5552 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_xcpt_pf_if : enq_buffer_0_dec_uops_3_xcpt_pf_if; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5553 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_xcpt_pf_if : _GEN_5552; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5554 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_xcpt_pf_if : _GEN_5553; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5555 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_xcpt_pf_if : _GEN_5554; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5556 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_xcpt_pf_if : _GEN_5555; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5557 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_xcpt_pf_if : _GEN_5556; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5558 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_xcpt_pf_if : _GEN_5557; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5560 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_fp_single : enq_buffer_0_dec_uops_3_fp_single; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5561 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_fp_single : _GEN_5560; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5562 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_fp_single : _GEN_5561; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5563 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_fp_single : _GEN_5562; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5564 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_fp_single : _GEN_5563; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5565 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_fp_single : _GEN_5564; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5566 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_fp_single : _GEN_5565; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5568 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_fp_val : enq_buffer_0_dec_uops_3_fp_val; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5569 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_fp_val : _GEN_5568; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5570 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_fp_val : _GEN_5569; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5571 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_fp_val : _GEN_5570; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5572 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_fp_val : _GEN_5571; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5573 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_fp_val : _GEN_5572; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5574 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_fp_val : _GEN_5573; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5576 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_frs3_en : enq_buffer_0_dec_uops_3_frs3_en; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5577 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_frs3_en : _GEN_5576; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5578 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_frs3_en : _GEN_5577; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5579 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_frs3_en : _GEN_5578; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5580 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_frs3_en : _GEN_5579; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5581 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_frs3_en : _GEN_5580; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5582 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_frs3_en : _GEN_5581; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5584 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_lrs2_rtype : enq_buffer_0_dec_uops_3_lrs2_rtype; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5585 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_lrs2_rtype : _GEN_5584; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5586 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_lrs2_rtype : _GEN_5585; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5587 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_lrs2_rtype : _GEN_5586; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5588 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_lrs2_rtype : _GEN_5587; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5589 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_lrs2_rtype : _GEN_5588; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5590 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_lrs2_rtype : _GEN_5589; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5592 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_lrs1_rtype : enq_buffer_0_dec_uops_3_lrs1_rtype; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5593 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_lrs1_rtype : _GEN_5592; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5594 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_lrs1_rtype : _GEN_5593; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5595 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_lrs1_rtype : _GEN_5594; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5596 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_lrs1_rtype : _GEN_5595; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5597 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_lrs1_rtype : _GEN_5596; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5598 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_lrs1_rtype : _GEN_5597; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5600 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_dst_rtype : enq_buffer_0_dec_uops_3_dst_rtype; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5601 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_dst_rtype : _GEN_5600; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5602 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_dst_rtype : _GEN_5601; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5603 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_dst_rtype : _GEN_5602; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5604 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_dst_rtype : _GEN_5603; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5605 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_dst_rtype : _GEN_5604; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5606 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_dst_rtype : _GEN_5605; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5608 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_ldst_val : enq_buffer_0_dec_uops_3_ldst_val; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5609 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_ldst_val : _GEN_5608; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5610 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_ldst_val : _GEN_5609; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5611 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_ldst_val : _GEN_5610; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5612 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_ldst_val : _GEN_5611; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5613 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_ldst_val : _GEN_5612; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5614 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_ldst_val : _GEN_5613; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5616 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_lrs3 : enq_buffer_0_dec_uops_3_lrs3; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5617 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_lrs3 : _GEN_5616; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5618 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_lrs3 : _GEN_5617; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5619 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_lrs3 : _GEN_5618; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5620 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_lrs3 : _GEN_5619; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5621 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_lrs3 : _GEN_5620; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5622 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_lrs3 : _GEN_5621; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5624 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_lrs2 : enq_buffer_0_dec_uops_3_lrs2; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5625 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_lrs2 : _GEN_5624; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5626 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_lrs2 : _GEN_5625; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5627 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_lrs2 : _GEN_5626; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5628 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_lrs2 : _GEN_5627; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5629 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_lrs2 : _GEN_5628; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5630 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_lrs2 : _GEN_5629; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5632 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_lrs1 : enq_buffer_0_dec_uops_3_lrs1; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5633 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_lrs1 : _GEN_5632; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5634 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_lrs1 : _GEN_5633; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5635 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_lrs1 : _GEN_5634; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5636 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_lrs1 : _GEN_5635; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5637 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_lrs1 : _GEN_5636; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5638 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_lrs1 : _GEN_5637; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5640 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_ldst : enq_buffer_0_dec_uops_3_ldst; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5641 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_ldst : _GEN_5640; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5642 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_ldst : _GEN_5641; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5643 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_ldst : _GEN_5642; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5644 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_ldst : _GEN_5643; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5645 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_ldst : _GEN_5644; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5646 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_ldst : _GEN_5645; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5648 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_ldst_is_rs1 : enq_buffer_0_dec_uops_3_ldst_is_rs1; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5649 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_ldst_is_rs1 : _GEN_5648; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5650 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_ldst_is_rs1 : _GEN_5649; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5651 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_ldst_is_rs1 : _GEN_5650; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5652 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_ldst_is_rs1 : _GEN_5651; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5653 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_ldst_is_rs1 : _GEN_5652; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5654 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_ldst_is_rs1 : _GEN_5653; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5656 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_flush_on_commit :
    enq_buffer_0_dec_uops_3_flush_on_commit; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5657 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_flush_on_commit : _GEN_5656; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5658 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_flush_on_commit : _GEN_5657; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5659 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_flush_on_commit : _GEN_5658; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5660 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_flush_on_commit : _GEN_5659; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5661 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_flush_on_commit : _GEN_5660; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5662 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_flush_on_commit : _GEN_5661; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5664 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_is_unique : enq_buffer_0_dec_uops_3_is_unique; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5665 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_is_unique : _GEN_5664; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5666 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_is_unique : _GEN_5665; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5667 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_is_unique : _GEN_5666; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5668 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_is_unique : _GEN_5667; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5669 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_is_unique : _GEN_5668; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5670 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_is_unique : _GEN_5669; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5672 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_is_sys_pc2epc : enq_buffer_0_dec_uops_3_is_sys_pc2epc
    ; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5673 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_is_sys_pc2epc : _GEN_5672; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5674 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_is_sys_pc2epc : _GEN_5673; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5675 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_is_sys_pc2epc : _GEN_5674; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5676 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_is_sys_pc2epc : _GEN_5675; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5677 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_is_sys_pc2epc : _GEN_5676; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5678 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_is_sys_pc2epc : _GEN_5677; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5680 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_uses_stq : enq_buffer_0_dec_uops_3_uses_stq; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5681 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_uses_stq : _GEN_5680; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5682 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_uses_stq : _GEN_5681; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5683 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_uses_stq : _GEN_5682; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5684 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_uses_stq : _GEN_5683; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5685 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_uses_stq : _GEN_5684; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5686 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_uses_stq : _GEN_5685; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5688 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_uses_ldq : enq_buffer_0_dec_uops_3_uses_ldq; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5689 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_uses_ldq : _GEN_5688; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5690 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_uses_ldq : _GEN_5689; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5691 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_uses_ldq : _GEN_5690; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5692 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_uses_ldq : _GEN_5691; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5693 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_uses_ldq : _GEN_5692; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5694 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_uses_ldq : _GEN_5693; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5696 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_is_amo : enq_buffer_0_dec_uops_3_is_amo; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5697 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_is_amo : _GEN_5696; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5698 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_is_amo : _GEN_5697; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5699 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_is_amo : _GEN_5698; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5700 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_is_amo : _GEN_5699; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5701 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_is_amo : _GEN_5700; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5702 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_is_amo : _GEN_5701; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5704 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_is_fencei : enq_buffer_0_dec_uops_3_is_fencei; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5705 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_is_fencei : _GEN_5704; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5706 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_is_fencei : _GEN_5705; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5707 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_is_fencei : _GEN_5706; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5708 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_is_fencei : _GEN_5707; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5709 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_is_fencei : _GEN_5708; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5710 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_is_fencei : _GEN_5709; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5712 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_is_fence : enq_buffer_0_dec_uops_3_is_fence; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5713 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_is_fence : _GEN_5712; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5714 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_is_fence : _GEN_5713; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5715 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_is_fence : _GEN_5714; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5716 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_is_fence : _GEN_5715; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5717 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_is_fence : _GEN_5716; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5718 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_is_fence : _GEN_5717; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5720 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_mem_signed : enq_buffer_0_dec_uops_3_mem_signed; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5721 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_mem_signed : _GEN_5720; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5722 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_mem_signed : _GEN_5721; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5723 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_mem_signed : _GEN_5722; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5724 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_mem_signed : _GEN_5723; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5725 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_mem_signed : _GEN_5724; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5726 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_mem_signed : _GEN_5725; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5728 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_mem_size : enq_buffer_0_dec_uops_3_mem_size; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5729 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_mem_size : _GEN_5728; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5730 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_mem_size : _GEN_5729; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5731 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_mem_size : _GEN_5730; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5732 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_mem_size : _GEN_5731; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5733 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_mem_size : _GEN_5732; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5734 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_mem_size : _GEN_5733; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5736 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_mem_cmd : enq_buffer_0_dec_uops_3_mem_cmd; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5737 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_mem_cmd : _GEN_5736; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5738 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_mem_cmd : _GEN_5737; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5739 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_mem_cmd : _GEN_5738; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5740 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_mem_cmd : _GEN_5739; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5741 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_mem_cmd : _GEN_5740; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5742 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_mem_cmd : _GEN_5741; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5744 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_bypassable : enq_buffer_0_dec_uops_3_bypassable; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5745 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_bypassable : _GEN_5744; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5746 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_bypassable : _GEN_5745; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5747 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_bypassable : _GEN_5746; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5748 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_bypassable : _GEN_5747; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5749 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_bypassable : _GEN_5748; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5750 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_bypassable : _GEN_5749; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_5752 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_exc_cause : enq_buffer_0_dec_uops_3_exc_cause; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_5753 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_exc_cause : _GEN_5752; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_5754 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_exc_cause : _GEN_5753; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_5755 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_exc_cause : _GEN_5754; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_5756 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_exc_cause : _GEN_5755; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_5757 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_exc_cause : _GEN_5756; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [63:0] _GEN_5758 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_exc_cause : _GEN_5757; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5760 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_exception : enq_buffer_0_dec_uops_3_exception; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5761 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_exception : _GEN_5760; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5762 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_exception : _GEN_5761; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5763 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_exception : _GEN_5762; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5764 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_exception : _GEN_5763; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5765 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_exception : _GEN_5764; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5766 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_exception : _GEN_5765; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5768 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_stale_pdst : enq_buffer_0_dec_uops_3_stale_pdst; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5769 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_stale_pdst : _GEN_5768; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5770 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_stale_pdst : _GEN_5769; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5771 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_stale_pdst : _GEN_5770; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5772 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_stale_pdst : _GEN_5771; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5773 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_stale_pdst : _GEN_5772; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5774 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_stale_pdst : _GEN_5773; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5776 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_ppred_busy : enq_buffer_0_dec_uops_3_ppred_busy; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5777 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_ppred_busy : _GEN_5776; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5778 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_ppred_busy : _GEN_5777; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5779 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_ppred_busy : _GEN_5778; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5780 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_ppred_busy : _GEN_5779; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5781 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_ppred_busy : _GEN_5780; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5782 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_ppred_busy : _GEN_5781; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5784 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_prs3_busy : enq_buffer_0_dec_uops_3_prs3_busy; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5785 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_prs3_busy : _GEN_5784; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5786 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_prs3_busy : _GEN_5785; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5787 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_prs3_busy : _GEN_5786; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5788 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_prs3_busy : _GEN_5787; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5789 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_prs3_busy : _GEN_5788; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5790 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_prs3_busy : _GEN_5789; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5792 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_prs2_busy : enq_buffer_0_dec_uops_3_prs2_busy; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5793 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_prs2_busy : _GEN_5792; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5794 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_prs2_busy : _GEN_5793; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5795 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_prs2_busy : _GEN_5794; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5796 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_prs2_busy : _GEN_5795; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5797 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_prs2_busy : _GEN_5796; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5798 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_prs2_busy : _GEN_5797; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5800 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_prs1_busy : enq_buffer_0_dec_uops_3_prs1_busy; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5801 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_prs1_busy : _GEN_5800; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5802 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_prs1_busy : _GEN_5801; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5803 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_prs1_busy : _GEN_5802; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5804 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_prs1_busy : _GEN_5803; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5805 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_prs1_busy : _GEN_5804; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5806 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_prs1_busy : _GEN_5805; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5808 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_ppred : enq_buffer_0_dec_uops_3_ppred; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5809 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_ppred : _GEN_5808; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5810 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_ppred : _GEN_5809; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5811 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_ppred : _GEN_5810; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5812 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_ppred : _GEN_5811; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5813 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_ppred : _GEN_5812; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5814 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_ppred : _GEN_5813; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5816 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_prs3 : enq_buffer_0_dec_uops_3_prs3; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5817 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_prs3 : _GEN_5816; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5818 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_prs3 : _GEN_5817; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5819 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_prs3 : _GEN_5818; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5820 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_prs3 : _GEN_5819; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5821 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_prs3 : _GEN_5820; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5822 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_prs3 : _GEN_5821; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5824 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_prs2 : enq_buffer_0_dec_uops_3_prs2; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5825 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_prs2 : _GEN_5824; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5826 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_prs2 : _GEN_5825; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5827 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_prs2 : _GEN_5826; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5828 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_prs2 : _GEN_5827; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5829 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_prs2 : _GEN_5828; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5830 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_prs2 : _GEN_5829; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5832 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_prs1 : enq_buffer_0_dec_uops_3_prs1; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5833 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_prs1 : _GEN_5832; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5834 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_prs1 : _GEN_5833; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5835 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_prs1 : _GEN_5834; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5836 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_prs1 : _GEN_5835; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5837 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_prs1 : _GEN_5836; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5838 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_prs1 : _GEN_5837; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5840 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_pdst : enq_buffer_0_dec_uops_3_pdst; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5841 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_pdst : _GEN_5840; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5842 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_pdst : _GEN_5841; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5843 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_pdst : _GEN_5842; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5844 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_pdst : _GEN_5843; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5845 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_pdst : _GEN_5844; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_5846 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_pdst : _GEN_5845; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5848 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_rxq_idx : enq_buffer_0_dec_uops_3_rxq_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5849 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_rxq_idx : _GEN_5848; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5850 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_rxq_idx : _GEN_5849; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5851 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_rxq_idx : _GEN_5850; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5852 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_rxq_idx : _GEN_5851; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5853 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_rxq_idx : _GEN_5852; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5854 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_rxq_idx : _GEN_5853; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5856 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_stq_idx : enq_buffer_0_dec_uops_3_stq_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5857 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_stq_idx : _GEN_5856; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5858 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_stq_idx : _GEN_5857; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5859 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_stq_idx : _GEN_5858; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5860 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_stq_idx : _GEN_5859; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5861 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_stq_idx : _GEN_5860; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5862 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_stq_idx : _GEN_5861; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5864 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_ldq_idx : enq_buffer_0_dec_uops_3_ldq_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5865 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_ldq_idx : _GEN_5864; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5866 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_ldq_idx : _GEN_5865; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5867 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_ldq_idx : _GEN_5866; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5868 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_ldq_idx : _GEN_5867; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5869 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_ldq_idx : _GEN_5868; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5870 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_ldq_idx : _GEN_5869; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5872 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_rob_idx : enq_buffer_0_dec_uops_3_rob_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5873 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_rob_idx : _GEN_5872; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5874 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_rob_idx : _GEN_5873; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5875 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_rob_idx : _GEN_5874; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5876 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_rob_idx : _GEN_5875; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5877 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_rob_idx : _GEN_5876; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5878 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_rob_idx : _GEN_5877; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5880 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_csr_addr : enq_buffer_0_dec_uops_3_csr_addr; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5881 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_csr_addr : _GEN_5880; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5882 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_csr_addr : _GEN_5881; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5883 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_csr_addr : _GEN_5882; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5884 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_csr_addr : _GEN_5883; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5885 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_csr_addr : _GEN_5884; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5886 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_csr_addr : _GEN_5885; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_5888 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_imm_packed : enq_buffer_0_dec_uops_3_imm_packed
    ; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_5889 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_imm_packed : _GEN_5888; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_5890 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_imm_packed : _GEN_5889; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_5891 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_imm_packed : _GEN_5890; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_5892 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_imm_packed : _GEN_5891; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_5893 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_imm_packed : _GEN_5892; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [19:0] _GEN_5894 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_imm_packed : _GEN_5893; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5896 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_taken : enq_buffer_0_dec_uops_3_taken; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5897 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_taken : _GEN_5896; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5898 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_taken : _GEN_5897; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5899 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_taken : _GEN_5898; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5900 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_taken : _GEN_5899; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5901 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_taken : _GEN_5900; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5902 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_taken : _GEN_5901; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5904 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_pc_lob : enq_buffer_0_dec_uops_3_pc_lob; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5905 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_pc_lob : _GEN_5904; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5906 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_pc_lob : _GEN_5905; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5907 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_pc_lob : _GEN_5906; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5908 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_pc_lob : _GEN_5907; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5909 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_pc_lob : _GEN_5908; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_5910 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_pc_lob : _GEN_5909; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5912 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_edge_inst : enq_buffer_0_dec_uops_3_edge_inst; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5913 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_edge_inst : _GEN_5912; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5914 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_edge_inst : _GEN_5913; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5915 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_edge_inst : _GEN_5914; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5916 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_edge_inst : _GEN_5915; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5917 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_edge_inst : _GEN_5916; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5918 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_edge_inst : _GEN_5917; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5920 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_ftq_idx : enq_buffer_0_dec_uops_3_ftq_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5921 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_ftq_idx : _GEN_5920; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5922 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_ftq_idx : _GEN_5921; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5923 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_ftq_idx : _GEN_5922; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5924 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_ftq_idx : _GEN_5923; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5925 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_ftq_idx : _GEN_5924; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [4:0] _GEN_5926 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_ftq_idx : _GEN_5925; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5928 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_br_tag : enq_buffer_0_dec_uops_3_br_tag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5929 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_br_tag : _GEN_5928; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5930 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_br_tag : _GEN_5929; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5931 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_br_tag : _GEN_5930; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5932 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_br_tag : _GEN_5931; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5933 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_br_tag : _GEN_5932; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_5934 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_br_tag : _GEN_5933; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5936 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_br_mask : enq_buffer_0_dec_uops_3_br_mask; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5937 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_br_mask : _GEN_5936; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5938 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_br_mask : _GEN_5937; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5939 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_br_mask : _GEN_5938; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5940 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_br_mask : _GEN_5939; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5941 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_br_mask : _GEN_5940; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [11:0] _GEN_5942 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_br_mask : _GEN_5941; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5944 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_is_sfb : enq_buffer_0_dec_uops_3_is_sfb; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5945 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_is_sfb : _GEN_5944; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5946 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_is_sfb : _GEN_5945; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5947 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_is_sfb : _GEN_5946; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5948 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_is_sfb : _GEN_5947; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5949 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_is_sfb : _GEN_5948; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5950 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_is_sfb : _GEN_5949; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5952 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_is_jal : enq_buffer_0_dec_uops_3_is_jal; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5953 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_is_jal : _GEN_5952; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5954 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_is_jal : _GEN_5953; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5955 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_is_jal : _GEN_5954; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5956 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_is_jal : _GEN_5955; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5957 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_is_jal : _GEN_5956; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5958 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_is_jal : _GEN_5957; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5960 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_is_jalr : enq_buffer_0_dec_uops_3_is_jalr; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5961 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_is_jalr : _GEN_5960; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5962 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_is_jalr : _GEN_5961; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5963 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_is_jalr : _GEN_5962; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5964 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_is_jalr : _GEN_5963; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5965 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_is_jalr : _GEN_5964; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5966 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_is_jalr : _GEN_5965; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5968 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_is_br : enq_buffer_0_dec_uops_3_is_br; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5969 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_is_br : _GEN_5968; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5970 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_is_br : _GEN_5969; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5971 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_is_br : _GEN_5970; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5972 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_is_br : _GEN_5971; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5973 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_is_br : _GEN_5972; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5974 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_is_br : _GEN_5973; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5976 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_iw_p2_poisoned :
    enq_buffer_0_dec_uops_3_iw_p2_poisoned; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5977 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_iw_p2_poisoned : _GEN_5976; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5978 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_iw_p2_poisoned : _GEN_5977; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5979 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_iw_p2_poisoned : _GEN_5978; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5980 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_iw_p2_poisoned : _GEN_5979; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5981 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_iw_p2_poisoned : _GEN_5980; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5982 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_iw_p2_poisoned : _GEN_5981; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5984 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_iw_p1_poisoned :
    enq_buffer_0_dec_uops_3_iw_p1_poisoned; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5985 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_iw_p1_poisoned : _GEN_5984; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5986 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_iw_p1_poisoned : _GEN_5985; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5987 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_iw_p1_poisoned : _GEN_5986; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5988 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_iw_p1_poisoned : _GEN_5987; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5989 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_iw_p1_poisoned : _GEN_5988; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_5990 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_iw_p1_poisoned : _GEN_5989; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5992 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_iw_state : enq_buffer_0_dec_uops_3_iw_state; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5993 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_iw_state : _GEN_5992; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5994 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_iw_state : _GEN_5993; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5995 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_iw_state : _GEN_5994; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5996 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_iw_state : _GEN_5995; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5997 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_iw_state : _GEN_5996; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_5998 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_iw_state : _GEN_5997; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_6000 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_ctrl_op3_sel :
    enq_buffer_0_dec_uops_3_ctrl_op3_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_6001 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_ctrl_op3_sel : _GEN_6000; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_6002 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_ctrl_op3_sel : _GEN_6001; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_6003 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_ctrl_op3_sel : _GEN_6002; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_6004 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_ctrl_op3_sel : _GEN_6003; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_6005 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_ctrl_op3_sel : _GEN_6004; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_6006 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_ctrl_op3_sel : _GEN_6005; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6008 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_ctrl_is_std : enq_buffer_0_dec_uops_3_ctrl_is_std; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6009 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_ctrl_is_std : _GEN_6008; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6010 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_ctrl_is_std : _GEN_6009; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6011 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_ctrl_is_std : _GEN_6010; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6012 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_ctrl_is_std : _GEN_6011; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6013 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_ctrl_is_std : _GEN_6012; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6014 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_ctrl_is_std : _GEN_6013; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6016 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_ctrl_is_sta : enq_buffer_0_dec_uops_3_ctrl_is_sta; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6017 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_ctrl_is_sta : _GEN_6016; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6018 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_ctrl_is_sta : _GEN_6017; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6019 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_ctrl_is_sta : _GEN_6018; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6020 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_ctrl_is_sta : _GEN_6019; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6021 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_ctrl_is_sta : _GEN_6020; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6022 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_ctrl_is_sta : _GEN_6021; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6024 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_ctrl_is_load : enq_buffer_0_dec_uops_3_ctrl_is_load; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6025 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_ctrl_is_load : _GEN_6024; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6026 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_ctrl_is_load : _GEN_6025; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6027 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_ctrl_is_load : _GEN_6026; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6028 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_ctrl_is_load : _GEN_6027; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6029 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_ctrl_is_load : _GEN_6028; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6030 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_ctrl_is_load : _GEN_6029; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6032 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_ctrl_csr_cmd :
    enq_buffer_0_dec_uops_3_ctrl_csr_cmd; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6033 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_ctrl_csr_cmd : _GEN_6032; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6034 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_ctrl_csr_cmd : _GEN_6033; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6035 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_ctrl_csr_cmd : _GEN_6034; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6036 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_ctrl_csr_cmd : _GEN_6035; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6037 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_ctrl_csr_cmd : _GEN_6036; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6038 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_ctrl_csr_cmd : _GEN_6037; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6040 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_ctrl_fcn_dw : enq_buffer_0_dec_uops_3_ctrl_fcn_dw; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6041 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_ctrl_fcn_dw : _GEN_6040; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6042 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_ctrl_fcn_dw : _GEN_6041; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6043 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_ctrl_fcn_dw : _GEN_6042; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6044 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_ctrl_fcn_dw : _GEN_6043; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6045 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_ctrl_fcn_dw : _GEN_6044; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6046 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_ctrl_fcn_dw : _GEN_6045; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6048 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_ctrl_op_fcn :
    enq_buffer_0_dec_uops_3_ctrl_op_fcn; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6049 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_ctrl_op_fcn : _GEN_6048; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6050 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_ctrl_op_fcn : _GEN_6049; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6051 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_ctrl_op_fcn : _GEN_6050; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6052 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_ctrl_op_fcn : _GEN_6051; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6053 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_ctrl_op_fcn : _GEN_6052; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6054 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_ctrl_op_fcn : _GEN_6053; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6056 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_ctrl_imm_sel :
    enq_buffer_0_dec_uops_3_ctrl_imm_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6057 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_ctrl_imm_sel : _GEN_6056; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6058 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_ctrl_imm_sel : _GEN_6057; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6059 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_ctrl_imm_sel : _GEN_6058; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6060 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_ctrl_imm_sel : _GEN_6059; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6061 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_ctrl_imm_sel : _GEN_6060; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6062 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_ctrl_imm_sel : _GEN_6061; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6064 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_ctrl_op2_sel :
    enq_buffer_0_dec_uops_3_ctrl_op2_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6065 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_ctrl_op2_sel : _GEN_6064; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6066 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_ctrl_op2_sel : _GEN_6065; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6067 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_ctrl_op2_sel : _GEN_6066; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6068 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_ctrl_op2_sel : _GEN_6067; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6069 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_ctrl_op2_sel : _GEN_6068; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6070 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_ctrl_op2_sel : _GEN_6069; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_6072 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_ctrl_op1_sel :
    enq_buffer_0_dec_uops_3_ctrl_op1_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_6073 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_ctrl_op1_sel : _GEN_6072; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_6074 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_ctrl_op1_sel : _GEN_6073; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_6075 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_ctrl_op1_sel : _GEN_6074; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_6076 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_ctrl_op1_sel : _GEN_6075; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_6077 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_ctrl_op1_sel : _GEN_6076; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_6078 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_ctrl_op1_sel : _GEN_6077; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6080 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_ctrl_br_type :
    enq_buffer_0_dec_uops_3_ctrl_br_type; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6081 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_ctrl_br_type : _GEN_6080; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6082 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_ctrl_br_type : _GEN_6081; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6083 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_ctrl_br_type : _GEN_6082; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6084 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_ctrl_br_type : _GEN_6083; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6085 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_ctrl_br_type : _GEN_6084; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6086 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_ctrl_br_type : _GEN_6085; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_6088 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_fu_code : enq_buffer_0_dec_uops_3_fu_code; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_6089 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_fu_code : _GEN_6088; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_6090 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_fu_code : _GEN_6089; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_6091 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_fu_code : _GEN_6090; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_6092 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_fu_code : _GEN_6091; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_6093 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_fu_code : _GEN_6092; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [9:0] _GEN_6094 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_fu_code : _GEN_6093; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6096 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_iq_type : enq_buffer_0_dec_uops_3_iq_type; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6097 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_iq_type : _GEN_6096; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6098 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_iq_type : _GEN_6097; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6099 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_iq_type : _GEN_6098; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6100 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_iq_type : _GEN_6099; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6101 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_iq_type : _GEN_6100; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6102 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_iq_type : _GEN_6101; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_6104 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_debug_pc : enq_buffer_0_dec_uops_3_debug_pc; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_6105 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_debug_pc : _GEN_6104; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_6106 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_debug_pc : _GEN_6105; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_6107 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_debug_pc : _GEN_6106; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_6108 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_debug_pc : _GEN_6107; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_6109 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_debug_pc : _GEN_6108; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [39:0] _GEN_6110 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_debug_pc : _GEN_6109; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6112 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_is_rvc : enq_buffer_0_dec_uops_3_is_rvc; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6113 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_is_rvc : _GEN_6112; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6114 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_is_rvc : _GEN_6113; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6115 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_is_rvc : _GEN_6114; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6116 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_is_rvc : _GEN_6115; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6117 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_is_rvc : _GEN_6116; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6118 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_is_rvc : _GEN_6117; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_6120 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_debug_inst : enq_buffer_0_dec_uops_3_debug_inst
    ; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_6121 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_debug_inst : _GEN_6120; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_6122 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_debug_inst : _GEN_6121; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_6123 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_debug_inst : _GEN_6122; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_6124 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_debug_inst : _GEN_6123; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_6125 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_debug_inst : _GEN_6124; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_6126 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_debug_inst : _GEN_6125; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_6128 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_inst : enq_buffer_0_dec_uops_3_inst; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_6129 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_inst : _GEN_6128; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_6130 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_inst : _GEN_6129; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_6131 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_inst : _GEN_6130; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_6132 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_inst : _GEN_6131; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_6133 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_inst : _GEN_6132; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [31:0] _GEN_6134 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_inst : _GEN_6133; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_6136 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_uopc : enq_buffer_0_dec_uops_3_uopc; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_6137 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_uopc : _GEN_6136; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_6138 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_uopc : _GEN_6137; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_6139 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_uopc : _GEN_6138; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_6140 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_uopc : _GEN_6139; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_6141 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_uopc : _GEN_6140; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [6:0] _GEN_6142 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_uopc : _GEN_6141; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6144 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_address_num :
    enq_buffer_0_dec_uops_3_address_num; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6145 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_address_num : _GEN_6144; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6146 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_address_num : _GEN_6145; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6147 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_address_num : _GEN_6146; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6148 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_address_num : _GEN_6147; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6149 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_address_num : _GEN_6148; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6150 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_address_num : _GEN_6149; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6152 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_rob_inst_idx :
    enq_buffer_0_dec_uops_3_rob_inst_idx; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6153 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_rob_inst_idx : _GEN_6152; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6154 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_rob_inst_idx : _GEN_6153; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6155 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_rob_inst_idx : _GEN_6154; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6156 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_rob_inst_idx : _GEN_6155; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6157 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_rob_inst_idx : _GEN_6156; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6158 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_rob_inst_idx : _GEN_6157; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6160 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_self_index : enq_buffer_0_dec_uops_3_self_index; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6161 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_self_index : _GEN_6160; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6162 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_self_index : _GEN_6161; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6163 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_self_index : _GEN_6162; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6164 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_self_index : _GEN_6163; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6165 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_self_index : _GEN_6164; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6166 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_self_index : _GEN_6165; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6168 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_split_num : enq_buffer_0_dec_uops_3_split_num; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6169 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_split_num : _GEN_6168; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6170 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_split_num : _GEN_6169; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6171 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_split_num : _GEN_6170; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6172 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_split_num : _GEN_6171; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6173 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_split_num : _GEN_6172; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [5:0] _GEN_6174 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_split_num : _GEN_6173; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6176 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_op2_sel : enq_buffer_0_dec_uops_3_op2_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6177 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_op2_sel : _GEN_6176; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6178 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_op2_sel : _GEN_6177; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6179 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_op2_sel : _GEN_6178; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6180 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_op2_sel : _GEN_6179; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6181 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_op2_sel : _GEN_6180; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6182 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_op2_sel : _GEN_6181; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6184 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_op1_sel : enq_buffer_0_dec_uops_3_op1_sel; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6185 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_op1_sel : _GEN_6184; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6186 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_op1_sel : _GEN_6185; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6187 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_op1_sel : _GEN_6186; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6188 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_op1_sel : _GEN_6187; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6189 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_op1_sel : _GEN_6188; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6190 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_op1_sel : _GEN_6189; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6192 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_stale_pflag :
    enq_buffer_0_dec_uops_3_stale_pflag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6193 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_stale_pflag : _GEN_6192; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6194 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_stale_pflag : _GEN_6193; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6195 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_stale_pflag : _GEN_6194; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6196 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_stale_pflag : _GEN_6195; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6197 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_stale_pflag : _GEN_6196; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6198 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_stale_pflag : _GEN_6197; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6200 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_pflag_busy : enq_buffer_0_dec_uops_3_pflag_busy; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6201 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_pflag_busy : _GEN_6200; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6202 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_pflag_busy : _GEN_6201; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6203 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_pflag_busy : _GEN_6202; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6204 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_pflag_busy : _GEN_6203; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6205 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_pflag_busy : _GEN_6204; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6206 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_pflag_busy : _GEN_6205; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6208 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_pwflag : enq_buffer_0_dec_uops_3_pwflag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6209 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_pwflag : _GEN_6208; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6210 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_pwflag : _GEN_6209; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6211 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_pwflag : _GEN_6210; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6212 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_pwflag : _GEN_6211; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6213 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_pwflag : _GEN_6212; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6214 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_pwflag : _GEN_6213; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6216 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_prflag : enq_buffer_0_dec_uops_3_prflag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6217 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_prflag : _GEN_6216; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6218 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_prflag : _GEN_6217; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6219 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_prflag : _GEN_6218; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6220 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_prflag : _GEN_6219; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6221 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_prflag : _GEN_6220; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [3:0] _GEN_6222 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_prflag : _GEN_6221; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6224 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_wflag : enq_buffer_0_dec_uops_3_wflag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6225 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_wflag : _GEN_6224; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6226 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_wflag : _GEN_6225; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6227 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_wflag : _GEN_6226; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6228 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_wflag : _GEN_6227; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6229 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_wflag : _GEN_6228; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6230 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_wflag : _GEN_6229; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6232 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_rflag : enq_buffer_0_dec_uops_3_rflag; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6233 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_rflag : _GEN_6232; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6234 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_rflag : _GEN_6233; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6235 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_rflag : _GEN_6234; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6236 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_rflag : _GEN_6235; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6237 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_rflag : _GEN_6236; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6238 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_rflag : _GEN_6237; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_6240 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_lrs3_rtype : enq_buffer_0_dec_uops_3_lrs3_rtype; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_6241 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_lrs3_rtype : _GEN_6240; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_6242 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_lrs3_rtype : _GEN_6241; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_6243 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_lrs3_rtype : _GEN_6242; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_6244 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_lrs3_rtype : _GEN_6243; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_6245 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_lrs3_rtype : _GEN_6244; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [1:0] _GEN_6246 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_lrs3_rtype : _GEN_6245; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6248 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_shift : enq_buffer_0_dec_uops_3_shift; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6249 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_shift : _GEN_6248; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6250 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_shift : _GEN_6249; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6251 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_shift : _GEN_6250; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6252 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_shift : _GEN_6251; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6253 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_shift : _GEN_6252; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire [2:0] _GEN_6254 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_shift : _GEN_6253; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6256 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_is_unicore : enq_buffer_0_dec_uops_3_is_unicore; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6257 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_is_unicore : _GEN_6256; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6258 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_is_unicore : _GEN_6257; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6259 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_is_unicore : _GEN_6258; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6260 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_is_unicore : _GEN_6259; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6261 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_is_unicore : _GEN_6260; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6262 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_is_unicore : _GEN_6261; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6264 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_switch_off : enq_buffer_0_dec_uops_3_switch_off; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6265 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_switch_off : _GEN_6264; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6266 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_switch_off : _GEN_6265; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6267 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_switch_off : _GEN_6266; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6268 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_switch_off : _GEN_6267; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6269 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_switch_off : _GEN_6268; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6270 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_switch_off : _GEN_6269; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6272 = 3'h1 == set_idx[2:0] ? enq_buffer_1_dec_uops_3_switch : enq_buffer_0_dec_uops_3_switch; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6273 = 3'h2 == set_idx[2:0] ? enq_buffer_2_dec_uops_3_switch : _GEN_6272; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6274 = 3'h3 == set_idx[2:0] ? enq_buffer_3_dec_uops_3_switch : _GEN_6273; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6275 = 3'h4 == set_idx[2:0] ? enq_buffer_4_dec_uops_3_switch : _GEN_6274; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6276 = 3'h5 == set_idx[2:0] ? enq_buffer_5_dec_uops_3_switch : _GEN_6275; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6277 = 3'h6 == set_idx[2:0] ? enq_buffer_6_dec_uops_3_switch : _GEN_6276; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  wire  _GEN_6278 = 3'h7 == set_idx[2:0] ? enq_buffer_7_dec_uops_3_switch : _GEN_6277; // @[enq_transBuff.scala 130:34 enq_transBuff.scala 130:34]
  TransBuffer trans_buffer ( // @[enq_transBuff.scala 37:31]
    .clock(trans_buffer_clock),
    .reset(trans_buffer_reset),
    .io_enq_ready(trans_buffer_io_enq_ready),
    .io_enq_valid(trans_buffer_io_enq_valid),
    .io_enq_bits_dec_uops_0_switch(trans_buffer_io_enq_bits_dec_uops_0_switch),
    .io_enq_bits_dec_uops_0_switch_off(trans_buffer_io_enq_bits_dec_uops_0_switch_off),
    .io_enq_bits_dec_uops_0_is_unicore(trans_buffer_io_enq_bits_dec_uops_0_is_unicore),
    .io_enq_bits_dec_uops_0_shift(trans_buffer_io_enq_bits_dec_uops_0_shift),
    .io_enq_bits_dec_uops_0_lrs3_rtype(trans_buffer_io_enq_bits_dec_uops_0_lrs3_rtype),
    .io_enq_bits_dec_uops_0_rflag(trans_buffer_io_enq_bits_dec_uops_0_rflag),
    .io_enq_bits_dec_uops_0_wflag(trans_buffer_io_enq_bits_dec_uops_0_wflag),
    .io_enq_bits_dec_uops_0_prflag(trans_buffer_io_enq_bits_dec_uops_0_prflag),
    .io_enq_bits_dec_uops_0_pwflag(trans_buffer_io_enq_bits_dec_uops_0_pwflag),
    .io_enq_bits_dec_uops_0_pflag_busy(trans_buffer_io_enq_bits_dec_uops_0_pflag_busy),
    .io_enq_bits_dec_uops_0_stale_pflag(trans_buffer_io_enq_bits_dec_uops_0_stale_pflag),
    .io_enq_bits_dec_uops_0_op1_sel(trans_buffer_io_enq_bits_dec_uops_0_op1_sel),
    .io_enq_bits_dec_uops_0_op2_sel(trans_buffer_io_enq_bits_dec_uops_0_op2_sel),
    .io_enq_bits_dec_uops_0_split_num(trans_buffer_io_enq_bits_dec_uops_0_split_num),
    .io_enq_bits_dec_uops_0_self_index(trans_buffer_io_enq_bits_dec_uops_0_self_index),
    .io_enq_bits_dec_uops_0_rob_inst_idx(trans_buffer_io_enq_bits_dec_uops_0_rob_inst_idx),
    .io_enq_bits_dec_uops_0_address_num(trans_buffer_io_enq_bits_dec_uops_0_address_num),
    .io_enq_bits_dec_uops_0_uopc(trans_buffer_io_enq_bits_dec_uops_0_uopc),
    .io_enq_bits_dec_uops_0_inst(trans_buffer_io_enq_bits_dec_uops_0_inst),
    .io_enq_bits_dec_uops_0_debug_inst(trans_buffer_io_enq_bits_dec_uops_0_debug_inst),
    .io_enq_bits_dec_uops_0_is_rvc(trans_buffer_io_enq_bits_dec_uops_0_is_rvc),
    .io_enq_bits_dec_uops_0_debug_pc(trans_buffer_io_enq_bits_dec_uops_0_debug_pc),
    .io_enq_bits_dec_uops_0_iq_type(trans_buffer_io_enq_bits_dec_uops_0_iq_type),
    .io_enq_bits_dec_uops_0_fu_code(trans_buffer_io_enq_bits_dec_uops_0_fu_code),
    .io_enq_bits_dec_uops_0_ctrl_br_type(trans_buffer_io_enq_bits_dec_uops_0_ctrl_br_type),
    .io_enq_bits_dec_uops_0_ctrl_op1_sel(trans_buffer_io_enq_bits_dec_uops_0_ctrl_op1_sel),
    .io_enq_bits_dec_uops_0_ctrl_op2_sel(trans_buffer_io_enq_bits_dec_uops_0_ctrl_op2_sel),
    .io_enq_bits_dec_uops_0_ctrl_imm_sel(trans_buffer_io_enq_bits_dec_uops_0_ctrl_imm_sel),
    .io_enq_bits_dec_uops_0_ctrl_op_fcn(trans_buffer_io_enq_bits_dec_uops_0_ctrl_op_fcn),
    .io_enq_bits_dec_uops_0_ctrl_fcn_dw(trans_buffer_io_enq_bits_dec_uops_0_ctrl_fcn_dw),
    .io_enq_bits_dec_uops_0_ctrl_csr_cmd(trans_buffer_io_enq_bits_dec_uops_0_ctrl_csr_cmd),
    .io_enq_bits_dec_uops_0_ctrl_is_load(trans_buffer_io_enq_bits_dec_uops_0_ctrl_is_load),
    .io_enq_bits_dec_uops_0_ctrl_is_sta(trans_buffer_io_enq_bits_dec_uops_0_ctrl_is_sta),
    .io_enq_bits_dec_uops_0_ctrl_is_std(trans_buffer_io_enq_bits_dec_uops_0_ctrl_is_std),
    .io_enq_bits_dec_uops_0_ctrl_op3_sel(trans_buffer_io_enq_bits_dec_uops_0_ctrl_op3_sel),
    .io_enq_bits_dec_uops_0_iw_state(trans_buffer_io_enq_bits_dec_uops_0_iw_state),
    .io_enq_bits_dec_uops_0_iw_p1_poisoned(trans_buffer_io_enq_bits_dec_uops_0_iw_p1_poisoned),
    .io_enq_bits_dec_uops_0_iw_p2_poisoned(trans_buffer_io_enq_bits_dec_uops_0_iw_p2_poisoned),
    .io_enq_bits_dec_uops_0_is_br(trans_buffer_io_enq_bits_dec_uops_0_is_br),
    .io_enq_bits_dec_uops_0_is_jalr(trans_buffer_io_enq_bits_dec_uops_0_is_jalr),
    .io_enq_bits_dec_uops_0_is_jal(trans_buffer_io_enq_bits_dec_uops_0_is_jal),
    .io_enq_bits_dec_uops_0_is_sfb(trans_buffer_io_enq_bits_dec_uops_0_is_sfb),
    .io_enq_bits_dec_uops_0_br_mask(trans_buffer_io_enq_bits_dec_uops_0_br_mask),
    .io_enq_bits_dec_uops_0_br_tag(trans_buffer_io_enq_bits_dec_uops_0_br_tag),
    .io_enq_bits_dec_uops_0_ftq_idx(trans_buffer_io_enq_bits_dec_uops_0_ftq_idx),
    .io_enq_bits_dec_uops_0_edge_inst(trans_buffer_io_enq_bits_dec_uops_0_edge_inst),
    .io_enq_bits_dec_uops_0_pc_lob(trans_buffer_io_enq_bits_dec_uops_0_pc_lob),
    .io_enq_bits_dec_uops_0_taken(trans_buffer_io_enq_bits_dec_uops_0_taken),
    .io_enq_bits_dec_uops_0_imm_packed(trans_buffer_io_enq_bits_dec_uops_0_imm_packed),
    .io_enq_bits_dec_uops_0_csr_addr(trans_buffer_io_enq_bits_dec_uops_0_csr_addr),
    .io_enq_bits_dec_uops_0_rob_idx(trans_buffer_io_enq_bits_dec_uops_0_rob_idx),
    .io_enq_bits_dec_uops_0_ldq_idx(trans_buffer_io_enq_bits_dec_uops_0_ldq_idx),
    .io_enq_bits_dec_uops_0_stq_idx(trans_buffer_io_enq_bits_dec_uops_0_stq_idx),
    .io_enq_bits_dec_uops_0_rxq_idx(trans_buffer_io_enq_bits_dec_uops_0_rxq_idx),
    .io_enq_bits_dec_uops_0_pdst(trans_buffer_io_enq_bits_dec_uops_0_pdst),
    .io_enq_bits_dec_uops_0_prs1(trans_buffer_io_enq_bits_dec_uops_0_prs1),
    .io_enq_bits_dec_uops_0_prs2(trans_buffer_io_enq_bits_dec_uops_0_prs2),
    .io_enq_bits_dec_uops_0_prs3(trans_buffer_io_enq_bits_dec_uops_0_prs3),
    .io_enq_bits_dec_uops_0_ppred(trans_buffer_io_enq_bits_dec_uops_0_ppred),
    .io_enq_bits_dec_uops_0_prs1_busy(trans_buffer_io_enq_bits_dec_uops_0_prs1_busy),
    .io_enq_bits_dec_uops_0_prs2_busy(trans_buffer_io_enq_bits_dec_uops_0_prs2_busy),
    .io_enq_bits_dec_uops_0_prs3_busy(trans_buffer_io_enq_bits_dec_uops_0_prs3_busy),
    .io_enq_bits_dec_uops_0_ppred_busy(trans_buffer_io_enq_bits_dec_uops_0_ppred_busy),
    .io_enq_bits_dec_uops_0_stale_pdst(trans_buffer_io_enq_bits_dec_uops_0_stale_pdst),
    .io_enq_bits_dec_uops_0_exception(trans_buffer_io_enq_bits_dec_uops_0_exception),
    .io_enq_bits_dec_uops_0_exc_cause(trans_buffer_io_enq_bits_dec_uops_0_exc_cause),
    .io_enq_bits_dec_uops_0_bypassable(trans_buffer_io_enq_bits_dec_uops_0_bypassable),
    .io_enq_bits_dec_uops_0_mem_cmd(trans_buffer_io_enq_bits_dec_uops_0_mem_cmd),
    .io_enq_bits_dec_uops_0_mem_size(trans_buffer_io_enq_bits_dec_uops_0_mem_size),
    .io_enq_bits_dec_uops_0_mem_signed(trans_buffer_io_enq_bits_dec_uops_0_mem_signed),
    .io_enq_bits_dec_uops_0_is_fence(trans_buffer_io_enq_bits_dec_uops_0_is_fence),
    .io_enq_bits_dec_uops_0_is_fencei(trans_buffer_io_enq_bits_dec_uops_0_is_fencei),
    .io_enq_bits_dec_uops_0_is_amo(trans_buffer_io_enq_bits_dec_uops_0_is_amo),
    .io_enq_bits_dec_uops_0_uses_ldq(trans_buffer_io_enq_bits_dec_uops_0_uses_ldq),
    .io_enq_bits_dec_uops_0_uses_stq(trans_buffer_io_enq_bits_dec_uops_0_uses_stq),
    .io_enq_bits_dec_uops_0_is_sys_pc2epc(trans_buffer_io_enq_bits_dec_uops_0_is_sys_pc2epc),
    .io_enq_bits_dec_uops_0_is_unique(trans_buffer_io_enq_bits_dec_uops_0_is_unique),
    .io_enq_bits_dec_uops_0_flush_on_commit(trans_buffer_io_enq_bits_dec_uops_0_flush_on_commit),
    .io_enq_bits_dec_uops_0_ldst_is_rs1(trans_buffer_io_enq_bits_dec_uops_0_ldst_is_rs1),
    .io_enq_bits_dec_uops_0_ldst(trans_buffer_io_enq_bits_dec_uops_0_ldst),
    .io_enq_bits_dec_uops_0_lrs1(trans_buffer_io_enq_bits_dec_uops_0_lrs1),
    .io_enq_bits_dec_uops_0_lrs2(trans_buffer_io_enq_bits_dec_uops_0_lrs2),
    .io_enq_bits_dec_uops_0_lrs3(trans_buffer_io_enq_bits_dec_uops_0_lrs3),
    .io_enq_bits_dec_uops_0_ldst_val(trans_buffer_io_enq_bits_dec_uops_0_ldst_val),
    .io_enq_bits_dec_uops_0_dst_rtype(trans_buffer_io_enq_bits_dec_uops_0_dst_rtype),
    .io_enq_bits_dec_uops_0_lrs1_rtype(trans_buffer_io_enq_bits_dec_uops_0_lrs1_rtype),
    .io_enq_bits_dec_uops_0_lrs2_rtype(trans_buffer_io_enq_bits_dec_uops_0_lrs2_rtype),
    .io_enq_bits_dec_uops_0_frs3_en(trans_buffer_io_enq_bits_dec_uops_0_frs3_en),
    .io_enq_bits_dec_uops_0_fp_val(trans_buffer_io_enq_bits_dec_uops_0_fp_val),
    .io_enq_bits_dec_uops_0_fp_single(trans_buffer_io_enq_bits_dec_uops_0_fp_single),
    .io_enq_bits_dec_uops_0_xcpt_pf_if(trans_buffer_io_enq_bits_dec_uops_0_xcpt_pf_if),
    .io_enq_bits_dec_uops_0_xcpt_ae_if(trans_buffer_io_enq_bits_dec_uops_0_xcpt_ae_if),
    .io_enq_bits_dec_uops_0_xcpt_ma_if(trans_buffer_io_enq_bits_dec_uops_0_xcpt_ma_if),
    .io_enq_bits_dec_uops_0_bp_debug_if(trans_buffer_io_enq_bits_dec_uops_0_bp_debug_if),
    .io_enq_bits_dec_uops_0_bp_xcpt_if(trans_buffer_io_enq_bits_dec_uops_0_bp_xcpt_if),
    .io_enq_bits_dec_uops_0_debug_fsrc(trans_buffer_io_enq_bits_dec_uops_0_debug_fsrc),
    .io_enq_bits_dec_uops_0_debug_tsrc(trans_buffer_io_enq_bits_dec_uops_0_debug_tsrc),
    .io_enq_bits_dec_uops_1_switch(trans_buffer_io_enq_bits_dec_uops_1_switch),
    .io_enq_bits_dec_uops_1_switch_off(trans_buffer_io_enq_bits_dec_uops_1_switch_off),
    .io_enq_bits_dec_uops_1_is_unicore(trans_buffer_io_enq_bits_dec_uops_1_is_unicore),
    .io_enq_bits_dec_uops_1_shift(trans_buffer_io_enq_bits_dec_uops_1_shift),
    .io_enq_bits_dec_uops_1_lrs3_rtype(trans_buffer_io_enq_bits_dec_uops_1_lrs3_rtype),
    .io_enq_bits_dec_uops_1_rflag(trans_buffer_io_enq_bits_dec_uops_1_rflag),
    .io_enq_bits_dec_uops_1_wflag(trans_buffer_io_enq_bits_dec_uops_1_wflag),
    .io_enq_bits_dec_uops_1_prflag(trans_buffer_io_enq_bits_dec_uops_1_prflag),
    .io_enq_bits_dec_uops_1_pwflag(trans_buffer_io_enq_bits_dec_uops_1_pwflag),
    .io_enq_bits_dec_uops_1_pflag_busy(trans_buffer_io_enq_bits_dec_uops_1_pflag_busy),
    .io_enq_bits_dec_uops_1_stale_pflag(trans_buffer_io_enq_bits_dec_uops_1_stale_pflag),
    .io_enq_bits_dec_uops_1_op1_sel(trans_buffer_io_enq_bits_dec_uops_1_op1_sel),
    .io_enq_bits_dec_uops_1_op2_sel(trans_buffer_io_enq_bits_dec_uops_1_op2_sel),
    .io_enq_bits_dec_uops_1_split_num(trans_buffer_io_enq_bits_dec_uops_1_split_num),
    .io_enq_bits_dec_uops_1_self_index(trans_buffer_io_enq_bits_dec_uops_1_self_index),
    .io_enq_bits_dec_uops_1_rob_inst_idx(trans_buffer_io_enq_bits_dec_uops_1_rob_inst_idx),
    .io_enq_bits_dec_uops_1_address_num(trans_buffer_io_enq_bits_dec_uops_1_address_num),
    .io_enq_bits_dec_uops_1_uopc(trans_buffer_io_enq_bits_dec_uops_1_uopc),
    .io_enq_bits_dec_uops_1_inst(trans_buffer_io_enq_bits_dec_uops_1_inst),
    .io_enq_bits_dec_uops_1_debug_inst(trans_buffer_io_enq_bits_dec_uops_1_debug_inst),
    .io_enq_bits_dec_uops_1_is_rvc(trans_buffer_io_enq_bits_dec_uops_1_is_rvc),
    .io_enq_bits_dec_uops_1_debug_pc(trans_buffer_io_enq_bits_dec_uops_1_debug_pc),
    .io_enq_bits_dec_uops_1_iq_type(trans_buffer_io_enq_bits_dec_uops_1_iq_type),
    .io_enq_bits_dec_uops_1_fu_code(trans_buffer_io_enq_bits_dec_uops_1_fu_code),
    .io_enq_bits_dec_uops_1_ctrl_br_type(trans_buffer_io_enq_bits_dec_uops_1_ctrl_br_type),
    .io_enq_bits_dec_uops_1_ctrl_op1_sel(trans_buffer_io_enq_bits_dec_uops_1_ctrl_op1_sel),
    .io_enq_bits_dec_uops_1_ctrl_op2_sel(trans_buffer_io_enq_bits_dec_uops_1_ctrl_op2_sel),
    .io_enq_bits_dec_uops_1_ctrl_imm_sel(trans_buffer_io_enq_bits_dec_uops_1_ctrl_imm_sel),
    .io_enq_bits_dec_uops_1_ctrl_op_fcn(trans_buffer_io_enq_bits_dec_uops_1_ctrl_op_fcn),
    .io_enq_bits_dec_uops_1_ctrl_fcn_dw(trans_buffer_io_enq_bits_dec_uops_1_ctrl_fcn_dw),
    .io_enq_bits_dec_uops_1_ctrl_csr_cmd(trans_buffer_io_enq_bits_dec_uops_1_ctrl_csr_cmd),
    .io_enq_bits_dec_uops_1_ctrl_is_load(trans_buffer_io_enq_bits_dec_uops_1_ctrl_is_load),
    .io_enq_bits_dec_uops_1_ctrl_is_sta(trans_buffer_io_enq_bits_dec_uops_1_ctrl_is_sta),
    .io_enq_bits_dec_uops_1_ctrl_is_std(trans_buffer_io_enq_bits_dec_uops_1_ctrl_is_std),
    .io_enq_bits_dec_uops_1_ctrl_op3_sel(trans_buffer_io_enq_bits_dec_uops_1_ctrl_op3_sel),
    .io_enq_bits_dec_uops_1_iw_state(trans_buffer_io_enq_bits_dec_uops_1_iw_state),
    .io_enq_bits_dec_uops_1_iw_p1_poisoned(trans_buffer_io_enq_bits_dec_uops_1_iw_p1_poisoned),
    .io_enq_bits_dec_uops_1_iw_p2_poisoned(trans_buffer_io_enq_bits_dec_uops_1_iw_p2_poisoned),
    .io_enq_bits_dec_uops_1_is_br(trans_buffer_io_enq_bits_dec_uops_1_is_br),
    .io_enq_bits_dec_uops_1_is_jalr(trans_buffer_io_enq_bits_dec_uops_1_is_jalr),
    .io_enq_bits_dec_uops_1_is_jal(trans_buffer_io_enq_bits_dec_uops_1_is_jal),
    .io_enq_bits_dec_uops_1_is_sfb(trans_buffer_io_enq_bits_dec_uops_1_is_sfb),
    .io_enq_bits_dec_uops_1_br_mask(trans_buffer_io_enq_bits_dec_uops_1_br_mask),
    .io_enq_bits_dec_uops_1_br_tag(trans_buffer_io_enq_bits_dec_uops_1_br_tag),
    .io_enq_bits_dec_uops_1_ftq_idx(trans_buffer_io_enq_bits_dec_uops_1_ftq_idx),
    .io_enq_bits_dec_uops_1_edge_inst(trans_buffer_io_enq_bits_dec_uops_1_edge_inst),
    .io_enq_bits_dec_uops_1_pc_lob(trans_buffer_io_enq_bits_dec_uops_1_pc_lob),
    .io_enq_bits_dec_uops_1_taken(trans_buffer_io_enq_bits_dec_uops_1_taken),
    .io_enq_bits_dec_uops_1_imm_packed(trans_buffer_io_enq_bits_dec_uops_1_imm_packed),
    .io_enq_bits_dec_uops_1_csr_addr(trans_buffer_io_enq_bits_dec_uops_1_csr_addr),
    .io_enq_bits_dec_uops_1_rob_idx(trans_buffer_io_enq_bits_dec_uops_1_rob_idx),
    .io_enq_bits_dec_uops_1_ldq_idx(trans_buffer_io_enq_bits_dec_uops_1_ldq_idx),
    .io_enq_bits_dec_uops_1_stq_idx(trans_buffer_io_enq_bits_dec_uops_1_stq_idx),
    .io_enq_bits_dec_uops_1_rxq_idx(trans_buffer_io_enq_bits_dec_uops_1_rxq_idx),
    .io_enq_bits_dec_uops_1_pdst(trans_buffer_io_enq_bits_dec_uops_1_pdst),
    .io_enq_bits_dec_uops_1_prs1(trans_buffer_io_enq_bits_dec_uops_1_prs1),
    .io_enq_bits_dec_uops_1_prs2(trans_buffer_io_enq_bits_dec_uops_1_prs2),
    .io_enq_bits_dec_uops_1_prs3(trans_buffer_io_enq_bits_dec_uops_1_prs3),
    .io_enq_bits_dec_uops_1_ppred(trans_buffer_io_enq_bits_dec_uops_1_ppred),
    .io_enq_bits_dec_uops_1_prs1_busy(trans_buffer_io_enq_bits_dec_uops_1_prs1_busy),
    .io_enq_bits_dec_uops_1_prs2_busy(trans_buffer_io_enq_bits_dec_uops_1_prs2_busy),
    .io_enq_bits_dec_uops_1_prs3_busy(trans_buffer_io_enq_bits_dec_uops_1_prs3_busy),
    .io_enq_bits_dec_uops_1_ppred_busy(trans_buffer_io_enq_bits_dec_uops_1_ppred_busy),
    .io_enq_bits_dec_uops_1_stale_pdst(trans_buffer_io_enq_bits_dec_uops_1_stale_pdst),
    .io_enq_bits_dec_uops_1_exception(trans_buffer_io_enq_bits_dec_uops_1_exception),
    .io_enq_bits_dec_uops_1_exc_cause(trans_buffer_io_enq_bits_dec_uops_1_exc_cause),
    .io_enq_bits_dec_uops_1_bypassable(trans_buffer_io_enq_bits_dec_uops_1_bypassable),
    .io_enq_bits_dec_uops_1_mem_cmd(trans_buffer_io_enq_bits_dec_uops_1_mem_cmd),
    .io_enq_bits_dec_uops_1_mem_size(trans_buffer_io_enq_bits_dec_uops_1_mem_size),
    .io_enq_bits_dec_uops_1_mem_signed(trans_buffer_io_enq_bits_dec_uops_1_mem_signed),
    .io_enq_bits_dec_uops_1_is_fence(trans_buffer_io_enq_bits_dec_uops_1_is_fence),
    .io_enq_bits_dec_uops_1_is_fencei(trans_buffer_io_enq_bits_dec_uops_1_is_fencei),
    .io_enq_bits_dec_uops_1_is_amo(trans_buffer_io_enq_bits_dec_uops_1_is_amo),
    .io_enq_bits_dec_uops_1_uses_ldq(trans_buffer_io_enq_bits_dec_uops_1_uses_ldq),
    .io_enq_bits_dec_uops_1_uses_stq(trans_buffer_io_enq_bits_dec_uops_1_uses_stq),
    .io_enq_bits_dec_uops_1_is_sys_pc2epc(trans_buffer_io_enq_bits_dec_uops_1_is_sys_pc2epc),
    .io_enq_bits_dec_uops_1_is_unique(trans_buffer_io_enq_bits_dec_uops_1_is_unique),
    .io_enq_bits_dec_uops_1_flush_on_commit(trans_buffer_io_enq_bits_dec_uops_1_flush_on_commit),
    .io_enq_bits_dec_uops_1_ldst_is_rs1(trans_buffer_io_enq_bits_dec_uops_1_ldst_is_rs1),
    .io_enq_bits_dec_uops_1_ldst(trans_buffer_io_enq_bits_dec_uops_1_ldst),
    .io_enq_bits_dec_uops_1_lrs1(trans_buffer_io_enq_bits_dec_uops_1_lrs1),
    .io_enq_bits_dec_uops_1_lrs2(trans_buffer_io_enq_bits_dec_uops_1_lrs2),
    .io_enq_bits_dec_uops_1_lrs3(trans_buffer_io_enq_bits_dec_uops_1_lrs3),
    .io_enq_bits_dec_uops_1_ldst_val(trans_buffer_io_enq_bits_dec_uops_1_ldst_val),
    .io_enq_bits_dec_uops_1_dst_rtype(trans_buffer_io_enq_bits_dec_uops_1_dst_rtype),
    .io_enq_bits_dec_uops_1_lrs1_rtype(trans_buffer_io_enq_bits_dec_uops_1_lrs1_rtype),
    .io_enq_bits_dec_uops_1_lrs2_rtype(trans_buffer_io_enq_bits_dec_uops_1_lrs2_rtype),
    .io_enq_bits_dec_uops_1_frs3_en(trans_buffer_io_enq_bits_dec_uops_1_frs3_en),
    .io_enq_bits_dec_uops_1_fp_val(trans_buffer_io_enq_bits_dec_uops_1_fp_val),
    .io_enq_bits_dec_uops_1_fp_single(trans_buffer_io_enq_bits_dec_uops_1_fp_single),
    .io_enq_bits_dec_uops_1_xcpt_pf_if(trans_buffer_io_enq_bits_dec_uops_1_xcpt_pf_if),
    .io_enq_bits_dec_uops_1_xcpt_ae_if(trans_buffer_io_enq_bits_dec_uops_1_xcpt_ae_if),
    .io_enq_bits_dec_uops_1_xcpt_ma_if(trans_buffer_io_enq_bits_dec_uops_1_xcpt_ma_if),
    .io_enq_bits_dec_uops_1_bp_debug_if(trans_buffer_io_enq_bits_dec_uops_1_bp_debug_if),
    .io_enq_bits_dec_uops_1_bp_xcpt_if(trans_buffer_io_enq_bits_dec_uops_1_bp_xcpt_if),
    .io_enq_bits_dec_uops_1_debug_fsrc(trans_buffer_io_enq_bits_dec_uops_1_debug_fsrc),
    .io_enq_bits_dec_uops_1_debug_tsrc(trans_buffer_io_enq_bits_dec_uops_1_debug_tsrc),
    .io_enq_bits_dec_uops_2_switch(trans_buffer_io_enq_bits_dec_uops_2_switch),
    .io_enq_bits_dec_uops_2_switch_off(trans_buffer_io_enq_bits_dec_uops_2_switch_off),
    .io_enq_bits_dec_uops_2_is_unicore(trans_buffer_io_enq_bits_dec_uops_2_is_unicore),
    .io_enq_bits_dec_uops_2_shift(trans_buffer_io_enq_bits_dec_uops_2_shift),
    .io_enq_bits_dec_uops_2_lrs3_rtype(trans_buffer_io_enq_bits_dec_uops_2_lrs3_rtype),
    .io_enq_bits_dec_uops_2_rflag(trans_buffer_io_enq_bits_dec_uops_2_rflag),
    .io_enq_bits_dec_uops_2_wflag(trans_buffer_io_enq_bits_dec_uops_2_wflag),
    .io_enq_bits_dec_uops_2_prflag(trans_buffer_io_enq_bits_dec_uops_2_prflag),
    .io_enq_bits_dec_uops_2_pwflag(trans_buffer_io_enq_bits_dec_uops_2_pwflag),
    .io_enq_bits_dec_uops_2_pflag_busy(trans_buffer_io_enq_bits_dec_uops_2_pflag_busy),
    .io_enq_bits_dec_uops_2_stale_pflag(trans_buffer_io_enq_bits_dec_uops_2_stale_pflag),
    .io_enq_bits_dec_uops_2_op1_sel(trans_buffer_io_enq_bits_dec_uops_2_op1_sel),
    .io_enq_bits_dec_uops_2_op2_sel(trans_buffer_io_enq_bits_dec_uops_2_op2_sel),
    .io_enq_bits_dec_uops_2_split_num(trans_buffer_io_enq_bits_dec_uops_2_split_num),
    .io_enq_bits_dec_uops_2_self_index(trans_buffer_io_enq_bits_dec_uops_2_self_index),
    .io_enq_bits_dec_uops_2_rob_inst_idx(trans_buffer_io_enq_bits_dec_uops_2_rob_inst_idx),
    .io_enq_bits_dec_uops_2_address_num(trans_buffer_io_enq_bits_dec_uops_2_address_num),
    .io_enq_bits_dec_uops_2_uopc(trans_buffer_io_enq_bits_dec_uops_2_uopc),
    .io_enq_bits_dec_uops_2_inst(trans_buffer_io_enq_bits_dec_uops_2_inst),
    .io_enq_bits_dec_uops_2_debug_inst(trans_buffer_io_enq_bits_dec_uops_2_debug_inst),
    .io_enq_bits_dec_uops_2_is_rvc(trans_buffer_io_enq_bits_dec_uops_2_is_rvc),
    .io_enq_bits_dec_uops_2_debug_pc(trans_buffer_io_enq_bits_dec_uops_2_debug_pc),
    .io_enq_bits_dec_uops_2_iq_type(trans_buffer_io_enq_bits_dec_uops_2_iq_type),
    .io_enq_bits_dec_uops_2_fu_code(trans_buffer_io_enq_bits_dec_uops_2_fu_code),
    .io_enq_bits_dec_uops_2_ctrl_br_type(trans_buffer_io_enq_bits_dec_uops_2_ctrl_br_type),
    .io_enq_bits_dec_uops_2_ctrl_op1_sel(trans_buffer_io_enq_bits_dec_uops_2_ctrl_op1_sel),
    .io_enq_bits_dec_uops_2_ctrl_op2_sel(trans_buffer_io_enq_bits_dec_uops_2_ctrl_op2_sel),
    .io_enq_bits_dec_uops_2_ctrl_imm_sel(trans_buffer_io_enq_bits_dec_uops_2_ctrl_imm_sel),
    .io_enq_bits_dec_uops_2_ctrl_op_fcn(trans_buffer_io_enq_bits_dec_uops_2_ctrl_op_fcn),
    .io_enq_bits_dec_uops_2_ctrl_fcn_dw(trans_buffer_io_enq_bits_dec_uops_2_ctrl_fcn_dw),
    .io_enq_bits_dec_uops_2_ctrl_csr_cmd(trans_buffer_io_enq_bits_dec_uops_2_ctrl_csr_cmd),
    .io_enq_bits_dec_uops_2_ctrl_is_load(trans_buffer_io_enq_bits_dec_uops_2_ctrl_is_load),
    .io_enq_bits_dec_uops_2_ctrl_is_sta(trans_buffer_io_enq_bits_dec_uops_2_ctrl_is_sta),
    .io_enq_bits_dec_uops_2_ctrl_is_std(trans_buffer_io_enq_bits_dec_uops_2_ctrl_is_std),
    .io_enq_bits_dec_uops_2_ctrl_op3_sel(trans_buffer_io_enq_bits_dec_uops_2_ctrl_op3_sel),
    .io_enq_bits_dec_uops_2_iw_state(trans_buffer_io_enq_bits_dec_uops_2_iw_state),
    .io_enq_bits_dec_uops_2_iw_p1_poisoned(trans_buffer_io_enq_bits_dec_uops_2_iw_p1_poisoned),
    .io_enq_bits_dec_uops_2_iw_p2_poisoned(trans_buffer_io_enq_bits_dec_uops_2_iw_p2_poisoned),
    .io_enq_bits_dec_uops_2_is_br(trans_buffer_io_enq_bits_dec_uops_2_is_br),
    .io_enq_bits_dec_uops_2_is_jalr(trans_buffer_io_enq_bits_dec_uops_2_is_jalr),
    .io_enq_bits_dec_uops_2_is_jal(trans_buffer_io_enq_bits_dec_uops_2_is_jal),
    .io_enq_bits_dec_uops_2_is_sfb(trans_buffer_io_enq_bits_dec_uops_2_is_sfb),
    .io_enq_bits_dec_uops_2_br_mask(trans_buffer_io_enq_bits_dec_uops_2_br_mask),
    .io_enq_bits_dec_uops_2_br_tag(trans_buffer_io_enq_bits_dec_uops_2_br_tag),
    .io_enq_bits_dec_uops_2_ftq_idx(trans_buffer_io_enq_bits_dec_uops_2_ftq_idx),
    .io_enq_bits_dec_uops_2_edge_inst(trans_buffer_io_enq_bits_dec_uops_2_edge_inst),
    .io_enq_bits_dec_uops_2_pc_lob(trans_buffer_io_enq_bits_dec_uops_2_pc_lob),
    .io_enq_bits_dec_uops_2_taken(trans_buffer_io_enq_bits_dec_uops_2_taken),
    .io_enq_bits_dec_uops_2_imm_packed(trans_buffer_io_enq_bits_dec_uops_2_imm_packed),
    .io_enq_bits_dec_uops_2_csr_addr(trans_buffer_io_enq_bits_dec_uops_2_csr_addr),
    .io_enq_bits_dec_uops_2_rob_idx(trans_buffer_io_enq_bits_dec_uops_2_rob_idx),
    .io_enq_bits_dec_uops_2_ldq_idx(trans_buffer_io_enq_bits_dec_uops_2_ldq_idx),
    .io_enq_bits_dec_uops_2_stq_idx(trans_buffer_io_enq_bits_dec_uops_2_stq_idx),
    .io_enq_bits_dec_uops_2_rxq_idx(trans_buffer_io_enq_bits_dec_uops_2_rxq_idx),
    .io_enq_bits_dec_uops_2_pdst(trans_buffer_io_enq_bits_dec_uops_2_pdst),
    .io_enq_bits_dec_uops_2_prs1(trans_buffer_io_enq_bits_dec_uops_2_prs1),
    .io_enq_bits_dec_uops_2_prs2(trans_buffer_io_enq_bits_dec_uops_2_prs2),
    .io_enq_bits_dec_uops_2_prs3(trans_buffer_io_enq_bits_dec_uops_2_prs3),
    .io_enq_bits_dec_uops_2_ppred(trans_buffer_io_enq_bits_dec_uops_2_ppred),
    .io_enq_bits_dec_uops_2_prs1_busy(trans_buffer_io_enq_bits_dec_uops_2_prs1_busy),
    .io_enq_bits_dec_uops_2_prs2_busy(trans_buffer_io_enq_bits_dec_uops_2_prs2_busy),
    .io_enq_bits_dec_uops_2_prs3_busy(trans_buffer_io_enq_bits_dec_uops_2_prs3_busy),
    .io_enq_bits_dec_uops_2_ppred_busy(trans_buffer_io_enq_bits_dec_uops_2_ppred_busy),
    .io_enq_bits_dec_uops_2_stale_pdst(trans_buffer_io_enq_bits_dec_uops_2_stale_pdst),
    .io_enq_bits_dec_uops_2_exception(trans_buffer_io_enq_bits_dec_uops_2_exception),
    .io_enq_bits_dec_uops_2_exc_cause(trans_buffer_io_enq_bits_dec_uops_2_exc_cause),
    .io_enq_bits_dec_uops_2_bypassable(trans_buffer_io_enq_bits_dec_uops_2_bypassable),
    .io_enq_bits_dec_uops_2_mem_cmd(trans_buffer_io_enq_bits_dec_uops_2_mem_cmd),
    .io_enq_bits_dec_uops_2_mem_size(trans_buffer_io_enq_bits_dec_uops_2_mem_size),
    .io_enq_bits_dec_uops_2_mem_signed(trans_buffer_io_enq_bits_dec_uops_2_mem_signed),
    .io_enq_bits_dec_uops_2_is_fence(trans_buffer_io_enq_bits_dec_uops_2_is_fence),
    .io_enq_bits_dec_uops_2_is_fencei(trans_buffer_io_enq_bits_dec_uops_2_is_fencei),
    .io_enq_bits_dec_uops_2_is_amo(trans_buffer_io_enq_bits_dec_uops_2_is_amo),
    .io_enq_bits_dec_uops_2_uses_ldq(trans_buffer_io_enq_bits_dec_uops_2_uses_ldq),
    .io_enq_bits_dec_uops_2_uses_stq(trans_buffer_io_enq_bits_dec_uops_2_uses_stq),
    .io_enq_bits_dec_uops_2_is_sys_pc2epc(trans_buffer_io_enq_bits_dec_uops_2_is_sys_pc2epc),
    .io_enq_bits_dec_uops_2_is_unique(trans_buffer_io_enq_bits_dec_uops_2_is_unique),
    .io_enq_bits_dec_uops_2_flush_on_commit(trans_buffer_io_enq_bits_dec_uops_2_flush_on_commit),
    .io_enq_bits_dec_uops_2_ldst_is_rs1(trans_buffer_io_enq_bits_dec_uops_2_ldst_is_rs1),
    .io_enq_bits_dec_uops_2_ldst(trans_buffer_io_enq_bits_dec_uops_2_ldst),
    .io_enq_bits_dec_uops_2_lrs1(trans_buffer_io_enq_bits_dec_uops_2_lrs1),
    .io_enq_bits_dec_uops_2_lrs2(trans_buffer_io_enq_bits_dec_uops_2_lrs2),
    .io_enq_bits_dec_uops_2_lrs3(trans_buffer_io_enq_bits_dec_uops_2_lrs3),
    .io_enq_bits_dec_uops_2_ldst_val(trans_buffer_io_enq_bits_dec_uops_2_ldst_val),
    .io_enq_bits_dec_uops_2_dst_rtype(trans_buffer_io_enq_bits_dec_uops_2_dst_rtype),
    .io_enq_bits_dec_uops_2_lrs1_rtype(trans_buffer_io_enq_bits_dec_uops_2_lrs1_rtype),
    .io_enq_bits_dec_uops_2_lrs2_rtype(trans_buffer_io_enq_bits_dec_uops_2_lrs2_rtype),
    .io_enq_bits_dec_uops_2_frs3_en(trans_buffer_io_enq_bits_dec_uops_2_frs3_en),
    .io_enq_bits_dec_uops_2_fp_val(trans_buffer_io_enq_bits_dec_uops_2_fp_val),
    .io_enq_bits_dec_uops_2_fp_single(trans_buffer_io_enq_bits_dec_uops_2_fp_single),
    .io_enq_bits_dec_uops_2_xcpt_pf_if(trans_buffer_io_enq_bits_dec_uops_2_xcpt_pf_if),
    .io_enq_bits_dec_uops_2_xcpt_ae_if(trans_buffer_io_enq_bits_dec_uops_2_xcpt_ae_if),
    .io_enq_bits_dec_uops_2_xcpt_ma_if(trans_buffer_io_enq_bits_dec_uops_2_xcpt_ma_if),
    .io_enq_bits_dec_uops_2_bp_debug_if(trans_buffer_io_enq_bits_dec_uops_2_bp_debug_if),
    .io_enq_bits_dec_uops_2_bp_xcpt_if(trans_buffer_io_enq_bits_dec_uops_2_bp_xcpt_if),
    .io_enq_bits_dec_uops_2_debug_fsrc(trans_buffer_io_enq_bits_dec_uops_2_debug_fsrc),
    .io_enq_bits_dec_uops_2_debug_tsrc(trans_buffer_io_enq_bits_dec_uops_2_debug_tsrc),
    .io_enq_bits_dec_uops_3_switch(trans_buffer_io_enq_bits_dec_uops_3_switch),
    .io_enq_bits_dec_uops_3_switch_off(trans_buffer_io_enq_bits_dec_uops_3_switch_off),
    .io_enq_bits_dec_uops_3_is_unicore(trans_buffer_io_enq_bits_dec_uops_3_is_unicore),
    .io_enq_bits_dec_uops_3_shift(trans_buffer_io_enq_bits_dec_uops_3_shift),
    .io_enq_bits_dec_uops_3_lrs3_rtype(trans_buffer_io_enq_bits_dec_uops_3_lrs3_rtype),
    .io_enq_bits_dec_uops_3_rflag(trans_buffer_io_enq_bits_dec_uops_3_rflag),
    .io_enq_bits_dec_uops_3_wflag(trans_buffer_io_enq_bits_dec_uops_3_wflag),
    .io_enq_bits_dec_uops_3_prflag(trans_buffer_io_enq_bits_dec_uops_3_prflag),
    .io_enq_bits_dec_uops_3_pwflag(trans_buffer_io_enq_bits_dec_uops_3_pwflag),
    .io_enq_bits_dec_uops_3_pflag_busy(trans_buffer_io_enq_bits_dec_uops_3_pflag_busy),
    .io_enq_bits_dec_uops_3_stale_pflag(trans_buffer_io_enq_bits_dec_uops_3_stale_pflag),
    .io_enq_bits_dec_uops_3_op1_sel(trans_buffer_io_enq_bits_dec_uops_3_op1_sel),
    .io_enq_bits_dec_uops_3_op2_sel(trans_buffer_io_enq_bits_dec_uops_3_op2_sel),
    .io_enq_bits_dec_uops_3_split_num(trans_buffer_io_enq_bits_dec_uops_3_split_num),
    .io_enq_bits_dec_uops_3_self_index(trans_buffer_io_enq_bits_dec_uops_3_self_index),
    .io_enq_bits_dec_uops_3_rob_inst_idx(trans_buffer_io_enq_bits_dec_uops_3_rob_inst_idx),
    .io_enq_bits_dec_uops_3_address_num(trans_buffer_io_enq_bits_dec_uops_3_address_num),
    .io_enq_bits_dec_uops_3_uopc(trans_buffer_io_enq_bits_dec_uops_3_uopc),
    .io_enq_bits_dec_uops_3_inst(trans_buffer_io_enq_bits_dec_uops_3_inst),
    .io_enq_bits_dec_uops_3_debug_inst(trans_buffer_io_enq_bits_dec_uops_3_debug_inst),
    .io_enq_bits_dec_uops_3_is_rvc(trans_buffer_io_enq_bits_dec_uops_3_is_rvc),
    .io_enq_bits_dec_uops_3_debug_pc(trans_buffer_io_enq_bits_dec_uops_3_debug_pc),
    .io_enq_bits_dec_uops_3_iq_type(trans_buffer_io_enq_bits_dec_uops_3_iq_type),
    .io_enq_bits_dec_uops_3_fu_code(trans_buffer_io_enq_bits_dec_uops_3_fu_code),
    .io_enq_bits_dec_uops_3_ctrl_br_type(trans_buffer_io_enq_bits_dec_uops_3_ctrl_br_type),
    .io_enq_bits_dec_uops_3_ctrl_op1_sel(trans_buffer_io_enq_bits_dec_uops_3_ctrl_op1_sel),
    .io_enq_bits_dec_uops_3_ctrl_op2_sel(trans_buffer_io_enq_bits_dec_uops_3_ctrl_op2_sel),
    .io_enq_bits_dec_uops_3_ctrl_imm_sel(trans_buffer_io_enq_bits_dec_uops_3_ctrl_imm_sel),
    .io_enq_bits_dec_uops_3_ctrl_op_fcn(trans_buffer_io_enq_bits_dec_uops_3_ctrl_op_fcn),
    .io_enq_bits_dec_uops_3_ctrl_fcn_dw(trans_buffer_io_enq_bits_dec_uops_3_ctrl_fcn_dw),
    .io_enq_bits_dec_uops_3_ctrl_csr_cmd(trans_buffer_io_enq_bits_dec_uops_3_ctrl_csr_cmd),
    .io_enq_bits_dec_uops_3_ctrl_is_load(trans_buffer_io_enq_bits_dec_uops_3_ctrl_is_load),
    .io_enq_bits_dec_uops_3_ctrl_is_sta(trans_buffer_io_enq_bits_dec_uops_3_ctrl_is_sta),
    .io_enq_bits_dec_uops_3_ctrl_is_std(trans_buffer_io_enq_bits_dec_uops_3_ctrl_is_std),
    .io_enq_bits_dec_uops_3_ctrl_op3_sel(trans_buffer_io_enq_bits_dec_uops_3_ctrl_op3_sel),
    .io_enq_bits_dec_uops_3_iw_state(trans_buffer_io_enq_bits_dec_uops_3_iw_state),
    .io_enq_bits_dec_uops_3_iw_p1_poisoned(trans_buffer_io_enq_bits_dec_uops_3_iw_p1_poisoned),
    .io_enq_bits_dec_uops_3_iw_p2_poisoned(trans_buffer_io_enq_bits_dec_uops_3_iw_p2_poisoned),
    .io_enq_bits_dec_uops_3_is_br(trans_buffer_io_enq_bits_dec_uops_3_is_br),
    .io_enq_bits_dec_uops_3_is_jalr(trans_buffer_io_enq_bits_dec_uops_3_is_jalr),
    .io_enq_bits_dec_uops_3_is_jal(trans_buffer_io_enq_bits_dec_uops_3_is_jal),
    .io_enq_bits_dec_uops_3_is_sfb(trans_buffer_io_enq_bits_dec_uops_3_is_sfb),
    .io_enq_bits_dec_uops_3_br_mask(trans_buffer_io_enq_bits_dec_uops_3_br_mask),
    .io_enq_bits_dec_uops_3_br_tag(trans_buffer_io_enq_bits_dec_uops_3_br_tag),
    .io_enq_bits_dec_uops_3_ftq_idx(trans_buffer_io_enq_bits_dec_uops_3_ftq_idx),
    .io_enq_bits_dec_uops_3_edge_inst(trans_buffer_io_enq_bits_dec_uops_3_edge_inst),
    .io_enq_bits_dec_uops_3_pc_lob(trans_buffer_io_enq_bits_dec_uops_3_pc_lob),
    .io_enq_bits_dec_uops_3_taken(trans_buffer_io_enq_bits_dec_uops_3_taken),
    .io_enq_bits_dec_uops_3_imm_packed(trans_buffer_io_enq_bits_dec_uops_3_imm_packed),
    .io_enq_bits_dec_uops_3_csr_addr(trans_buffer_io_enq_bits_dec_uops_3_csr_addr),
    .io_enq_bits_dec_uops_3_rob_idx(trans_buffer_io_enq_bits_dec_uops_3_rob_idx),
    .io_enq_bits_dec_uops_3_ldq_idx(trans_buffer_io_enq_bits_dec_uops_3_ldq_idx),
    .io_enq_bits_dec_uops_3_stq_idx(trans_buffer_io_enq_bits_dec_uops_3_stq_idx),
    .io_enq_bits_dec_uops_3_rxq_idx(trans_buffer_io_enq_bits_dec_uops_3_rxq_idx),
    .io_enq_bits_dec_uops_3_pdst(trans_buffer_io_enq_bits_dec_uops_3_pdst),
    .io_enq_bits_dec_uops_3_prs1(trans_buffer_io_enq_bits_dec_uops_3_prs1),
    .io_enq_bits_dec_uops_3_prs2(trans_buffer_io_enq_bits_dec_uops_3_prs2),
    .io_enq_bits_dec_uops_3_prs3(trans_buffer_io_enq_bits_dec_uops_3_prs3),
    .io_enq_bits_dec_uops_3_ppred(trans_buffer_io_enq_bits_dec_uops_3_ppred),
    .io_enq_bits_dec_uops_3_prs1_busy(trans_buffer_io_enq_bits_dec_uops_3_prs1_busy),
    .io_enq_bits_dec_uops_3_prs2_busy(trans_buffer_io_enq_bits_dec_uops_3_prs2_busy),
    .io_enq_bits_dec_uops_3_prs3_busy(trans_buffer_io_enq_bits_dec_uops_3_prs3_busy),
    .io_enq_bits_dec_uops_3_ppred_busy(trans_buffer_io_enq_bits_dec_uops_3_ppred_busy),
    .io_enq_bits_dec_uops_3_stale_pdst(trans_buffer_io_enq_bits_dec_uops_3_stale_pdst),
    .io_enq_bits_dec_uops_3_exception(trans_buffer_io_enq_bits_dec_uops_3_exception),
    .io_enq_bits_dec_uops_3_exc_cause(trans_buffer_io_enq_bits_dec_uops_3_exc_cause),
    .io_enq_bits_dec_uops_3_bypassable(trans_buffer_io_enq_bits_dec_uops_3_bypassable),
    .io_enq_bits_dec_uops_3_mem_cmd(trans_buffer_io_enq_bits_dec_uops_3_mem_cmd),
    .io_enq_bits_dec_uops_3_mem_size(trans_buffer_io_enq_bits_dec_uops_3_mem_size),
    .io_enq_bits_dec_uops_3_mem_signed(trans_buffer_io_enq_bits_dec_uops_3_mem_signed),
    .io_enq_bits_dec_uops_3_is_fence(trans_buffer_io_enq_bits_dec_uops_3_is_fence),
    .io_enq_bits_dec_uops_3_is_fencei(trans_buffer_io_enq_bits_dec_uops_3_is_fencei),
    .io_enq_bits_dec_uops_3_is_amo(trans_buffer_io_enq_bits_dec_uops_3_is_amo),
    .io_enq_bits_dec_uops_3_uses_ldq(trans_buffer_io_enq_bits_dec_uops_3_uses_ldq),
    .io_enq_bits_dec_uops_3_uses_stq(trans_buffer_io_enq_bits_dec_uops_3_uses_stq),
    .io_enq_bits_dec_uops_3_is_sys_pc2epc(trans_buffer_io_enq_bits_dec_uops_3_is_sys_pc2epc),
    .io_enq_bits_dec_uops_3_is_unique(trans_buffer_io_enq_bits_dec_uops_3_is_unique),
    .io_enq_bits_dec_uops_3_flush_on_commit(trans_buffer_io_enq_bits_dec_uops_3_flush_on_commit),
    .io_enq_bits_dec_uops_3_ldst_is_rs1(trans_buffer_io_enq_bits_dec_uops_3_ldst_is_rs1),
    .io_enq_bits_dec_uops_3_ldst(trans_buffer_io_enq_bits_dec_uops_3_ldst),
    .io_enq_bits_dec_uops_3_lrs1(trans_buffer_io_enq_bits_dec_uops_3_lrs1),
    .io_enq_bits_dec_uops_3_lrs2(trans_buffer_io_enq_bits_dec_uops_3_lrs2),
    .io_enq_bits_dec_uops_3_lrs3(trans_buffer_io_enq_bits_dec_uops_3_lrs3),
    .io_enq_bits_dec_uops_3_ldst_val(trans_buffer_io_enq_bits_dec_uops_3_ldst_val),
    .io_enq_bits_dec_uops_3_dst_rtype(trans_buffer_io_enq_bits_dec_uops_3_dst_rtype),
    .io_enq_bits_dec_uops_3_lrs1_rtype(trans_buffer_io_enq_bits_dec_uops_3_lrs1_rtype),
    .io_enq_bits_dec_uops_3_lrs2_rtype(trans_buffer_io_enq_bits_dec_uops_3_lrs2_rtype),
    .io_enq_bits_dec_uops_3_frs3_en(trans_buffer_io_enq_bits_dec_uops_3_frs3_en),
    .io_enq_bits_dec_uops_3_fp_val(trans_buffer_io_enq_bits_dec_uops_3_fp_val),
    .io_enq_bits_dec_uops_3_fp_single(trans_buffer_io_enq_bits_dec_uops_3_fp_single),
    .io_enq_bits_dec_uops_3_xcpt_pf_if(trans_buffer_io_enq_bits_dec_uops_3_xcpt_pf_if),
    .io_enq_bits_dec_uops_3_xcpt_ae_if(trans_buffer_io_enq_bits_dec_uops_3_xcpt_ae_if),
    .io_enq_bits_dec_uops_3_xcpt_ma_if(trans_buffer_io_enq_bits_dec_uops_3_xcpt_ma_if),
    .io_enq_bits_dec_uops_3_bp_debug_if(trans_buffer_io_enq_bits_dec_uops_3_bp_debug_if),
    .io_enq_bits_dec_uops_3_bp_xcpt_if(trans_buffer_io_enq_bits_dec_uops_3_bp_xcpt_if),
    .io_enq_bits_dec_uops_3_debug_fsrc(trans_buffer_io_enq_bits_dec_uops_3_debug_fsrc),
    .io_enq_bits_dec_uops_3_debug_tsrc(trans_buffer_io_enq_bits_dec_uops_3_debug_tsrc),
    .io_enq_bits_val_mask_0(trans_buffer_io_enq_bits_val_mask_0),
    .io_enq_bits_val_mask_1(trans_buffer_io_enq_bits_val_mask_1),
    .io_enq_bits_val_mask_2(trans_buffer_io_enq_bits_val_mask_2),
    .io_enq_bits_val_mask_3(trans_buffer_io_enq_bits_val_mask_3),
    .io_deq_ready(trans_buffer_io_deq_ready),
    .io_deq_valid(trans_buffer_io_deq_valid),
    .io_deq_bits_tran_uops_0_switch(trans_buffer_io_deq_bits_tran_uops_0_switch),
    .io_deq_bits_tran_uops_0_switch_off(trans_buffer_io_deq_bits_tran_uops_0_switch_off),
    .io_deq_bits_tran_uops_0_is_unicore(trans_buffer_io_deq_bits_tran_uops_0_is_unicore),
    .io_deq_bits_tran_uops_0_shift(trans_buffer_io_deq_bits_tran_uops_0_shift),
    .io_deq_bits_tran_uops_0_lrs3_rtype(trans_buffer_io_deq_bits_tran_uops_0_lrs3_rtype),
    .io_deq_bits_tran_uops_0_rflag(trans_buffer_io_deq_bits_tran_uops_0_rflag),
    .io_deq_bits_tran_uops_0_wflag(trans_buffer_io_deq_bits_tran_uops_0_wflag),
    .io_deq_bits_tran_uops_0_prflag(trans_buffer_io_deq_bits_tran_uops_0_prflag),
    .io_deq_bits_tran_uops_0_pwflag(trans_buffer_io_deq_bits_tran_uops_0_pwflag),
    .io_deq_bits_tran_uops_0_pflag_busy(trans_buffer_io_deq_bits_tran_uops_0_pflag_busy),
    .io_deq_bits_tran_uops_0_stale_pflag(trans_buffer_io_deq_bits_tran_uops_0_stale_pflag),
    .io_deq_bits_tran_uops_0_op1_sel(trans_buffer_io_deq_bits_tran_uops_0_op1_sel),
    .io_deq_bits_tran_uops_0_op2_sel(trans_buffer_io_deq_bits_tran_uops_0_op2_sel),
    .io_deq_bits_tran_uops_0_split_num(trans_buffer_io_deq_bits_tran_uops_0_split_num),
    .io_deq_bits_tran_uops_0_self_index(trans_buffer_io_deq_bits_tran_uops_0_self_index),
    .io_deq_bits_tran_uops_0_rob_inst_idx(trans_buffer_io_deq_bits_tran_uops_0_rob_inst_idx),
    .io_deq_bits_tran_uops_0_address_num(trans_buffer_io_deq_bits_tran_uops_0_address_num),
    .io_deq_bits_tran_uops_0_uopc(trans_buffer_io_deq_bits_tran_uops_0_uopc),
    .io_deq_bits_tran_uops_0_inst(trans_buffer_io_deq_bits_tran_uops_0_inst),
    .io_deq_bits_tran_uops_0_debug_inst(trans_buffer_io_deq_bits_tran_uops_0_debug_inst),
    .io_deq_bits_tran_uops_0_is_rvc(trans_buffer_io_deq_bits_tran_uops_0_is_rvc),
    .io_deq_bits_tran_uops_0_debug_pc(trans_buffer_io_deq_bits_tran_uops_0_debug_pc),
    .io_deq_bits_tran_uops_0_iq_type(trans_buffer_io_deq_bits_tran_uops_0_iq_type),
    .io_deq_bits_tran_uops_0_fu_code(trans_buffer_io_deq_bits_tran_uops_0_fu_code),
    .io_deq_bits_tran_uops_0_ctrl_br_type(trans_buffer_io_deq_bits_tran_uops_0_ctrl_br_type),
    .io_deq_bits_tran_uops_0_ctrl_op1_sel(trans_buffer_io_deq_bits_tran_uops_0_ctrl_op1_sel),
    .io_deq_bits_tran_uops_0_ctrl_op2_sel(trans_buffer_io_deq_bits_tran_uops_0_ctrl_op2_sel),
    .io_deq_bits_tran_uops_0_ctrl_imm_sel(trans_buffer_io_deq_bits_tran_uops_0_ctrl_imm_sel),
    .io_deq_bits_tran_uops_0_ctrl_op_fcn(trans_buffer_io_deq_bits_tran_uops_0_ctrl_op_fcn),
    .io_deq_bits_tran_uops_0_ctrl_fcn_dw(trans_buffer_io_deq_bits_tran_uops_0_ctrl_fcn_dw),
    .io_deq_bits_tran_uops_0_ctrl_csr_cmd(trans_buffer_io_deq_bits_tran_uops_0_ctrl_csr_cmd),
    .io_deq_bits_tran_uops_0_ctrl_is_load(trans_buffer_io_deq_bits_tran_uops_0_ctrl_is_load),
    .io_deq_bits_tran_uops_0_ctrl_is_sta(trans_buffer_io_deq_bits_tran_uops_0_ctrl_is_sta),
    .io_deq_bits_tran_uops_0_ctrl_is_std(trans_buffer_io_deq_bits_tran_uops_0_ctrl_is_std),
    .io_deq_bits_tran_uops_0_ctrl_op3_sel(trans_buffer_io_deq_bits_tran_uops_0_ctrl_op3_sel),
    .io_deq_bits_tran_uops_0_iw_state(trans_buffer_io_deq_bits_tran_uops_0_iw_state),
    .io_deq_bits_tran_uops_0_iw_p1_poisoned(trans_buffer_io_deq_bits_tran_uops_0_iw_p1_poisoned),
    .io_deq_bits_tran_uops_0_iw_p2_poisoned(trans_buffer_io_deq_bits_tran_uops_0_iw_p2_poisoned),
    .io_deq_bits_tran_uops_0_is_br(trans_buffer_io_deq_bits_tran_uops_0_is_br),
    .io_deq_bits_tran_uops_0_is_jalr(trans_buffer_io_deq_bits_tran_uops_0_is_jalr),
    .io_deq_bits_tran_uops_0_is_jal(trans_buffer_io_deq_bits_tran_uops_0_is_jal),
    .io_deq_bits_tran_uops_0_is_sfb(trans_buffer_io_deq_bits_tran_uops_0_is_sfb),
    .io_deq_bits_tran_uops_0_br_mask(trans_buffer_io_deq_bits_tran_uops_0_br_mask),
    .io_deq_bits_tran_uops_0_br_tag(trans_buffer_io_deq_bits_tran_uops_0_br_tag),
    .io_deq_bits_tran_uops_0_ftq_idx(trans_buffer_io_deq_bits_tran_uops_0_ftq_idx),
    .io_deq_bits_tran_uops_0_edge_inst(trans_buffer_io_deq_bits_tran_uops_0_edge_inst),
    .io_deq_bits_tran_uops_0_pc_lob(trans_buffer_io_deq_bits_tran_uops_0_pc_lob),
    .io_deq_bits_tran_uops_0_taken(trans_buffer_io_deq_bits_tran_uops_0_taken),
    .io_deq_bits_tran_uops_0_imm_packed(trans_buffer_io_deq_bits_tran_uops_0_imm_packed),
    .io_deq_bits_tran_uops_0_csr_addr(trans_buffer_io_deq_bits_tran_uops_0_csr_addr),
    .io_deq_bits_tran_uops_0_rob_idx(trans_buffer_io_deq_bits_tran_uops_0_rob_idx),
    .io_deq_bits_tran_uops_0_ldq_idx(trans_buffer_io_deq_bits_tran_uops_0_ldq_idx),
    .io_deq_bits_tran_uops_0_stq_idx(trans_buffer_io_deq_bits_tran_uops_0_stq_idx),
    .io_deq_bits_tran_uops_0_rxq_idx(trans_buffer_io_deq_bits_tran_uops_0_rxq_idx),
    .io_deq_bits_tran_uops_0_pdst(trans_buffer_io_deq_bits_tran_uops_0_pdst),
    .io_deq_bits_tran_uops_0_prs1(trans_buffer_io_deq_bits_tran_uops_0_prs1),
    .io_deq_bits_tran_uops_0_prs2(trans_buffer_io_deq_bits_tran_uops_0_prs2),
    .io_deq_bits_tran_uops_0_prs3(trans_buffer_io_deq_bits_tran_uops_0_prs3),
    .io_deq_bits_tran_uops_0_ppred(trans_buffer_io_deq_bits_tran_uops_0_ppred),
    .io_deq_bits_tran_uops_0_prs1_busy(trans_buffer_io_deq_bits_tran_uops_0_prs1_busy),
    .io_deq_bits_tran_uops_0_prs2_busy(trans_buffer_io_deq_bits_tran_uops_0_prs2_busy),
    .io_deq_bits_tran_uops_0_prs3_busy(trans_buffer_io_deq_bits_tran_uops_0_prs3_busy),
    .io_deq_bits_tran_uops_0_ppred_busy(trans_buffer_io_deq_bits_tran_uops_0_ppred_busy),
    .io_deq_bits_tran_uops_0_stale_pdst(trans_buffer_io_deq_bits_tran_uops_0_stale_pdst),
    .io_deq_bits_tran_uops_0_exception(trans_buffer_io_deq_bits_tran_uops_0_exception),
    .io_deq_bits_tran_uops_0_exc_cause(trans_buffer_io_deq_bits_tran_uops_0_exc_cause),
    .io_deq_bits_tran_uops_0_bypassable(trans_buffer_io_deq_bits_tran_uops_0_bypassable),
    .io_deq_bits_tran_uops_0_mem_cmd(trans_buffer_io_deq_bits_tran_uops_0_mem_cmd),
    .io_deq_bits_tran_uops_0_mem_size(trans_buffer_io_deq_bits_tran_uops_0_mem_size),
    .io_deq_bits_tran_uops_0_mem_signed(trans_buffer_io_deq_bits_tran_uops_0_mem_signed),
    .io_deq_bits_tran_uops_0_is_fence(trans_buffer_io_deq_bits_tran_uops_0_is_fence),
    .io_deq_bits_tran_uops_0_is_fencei(trans_buffer_io_deq_bits_tran_uops_0_is_fencei),
    .io_deq_bits_tran_uops_0_is_amo(trans_buffer_io_deq_bits_tran_uops_0_is_amo),
    .io_deq_bits_tran_uops_0_uses_ldq(trans_buffer_io_deq_bits_tran_uops_0_uses_ldq),
    .io_deq_bits_tran_uops_0_uses_stq(trans_buffer_io_deq_bits_tran_uops_0_uses_stq),
    .io_deq_bits_tran_uops_0_is_sys_pc2epc(trans_buffer_io_deq_bits_tran_uops_0_is_sys_pc2epc),
    .io_deq_bits_tran_uops_0_is_unique(trans_buffer_io_deq_bits_tran_uops_0_is_unique),
    .io_deq_bits_tran_uops_0_flush_on_commit(trans_buffer_io_deq_bits_tran_uops_0_flush_on_commit),
    .io_deq_bits_tran_uops_0_ldst_is_rs1(trans_buffer_io_deq_bits_tran_uops_0_ldst_is_rs1),
    .io_deq_bits_tran_uops_0_ldst(trans_buffer_io_deq_bits_tran_uops_0_ldst),
    .io_deq_bits_tran_uops_0_lrs1(trans_buffer_io_deq_bits_tran_uops_0_lrs1),
    .io_deq_bits_tran_uops_0_lrs2(trans_buffer_io_deq_bits_tran_uops_0_lrs2),
    .io_deq_bits_tran_uops_0_lrs3(trans_buffer_io_deq_bits_tran_uops_0_lrs3),
    .io_deq_bits_tran_uops_0_ldst_val(trans_buffer_io_deq_bits_tran_uops_0_ldst_val),
    .io_deq_bits_tran_uops_0_dst_rtype(trans_buffer_io_deq_bits_tran_uops_0_dst_rtype),
    .io_deq_bits_tran_uops_0_lrs1_rtype(trans_buffer_io_deq_bits_tran_uops_0_lrs1_rtype),
    .io_deq_bits_tran_uops_0_lrs2_rtype(trans_buffer_io_deq_bits_tran_uops_0_lrs2_rtype),
    .io_deq_bits_tran_uops_0_frs3_en(trans_buffer_io_deq_bits_tran_uops_0_frs3_en),
    .io_deq_bits_tran_uops_0_fp_val(trans_buffer_io_deq_bits_tran_uops_0_fp_val),
    .io_deq_bits_tran_uops_0_fp_single(trans_buffer_io_deq_bits_tran_uops_0_fp_single),
    .io_deq_bits_tran_uops_0_xcpt_pf_if(trans_buffer_io_deq_bits_tran_uops_0_xcpt_pf_if),
    .io_deq_bits_tran_uops_0_xcpt_ae_if(trans_buffer_io_deq_bits_tran_uops_0_xcpt_ae_if),
    .io_deq_bits_tran_uops_0_xcpt_ma_if(trans_buffer_io_deq_bits_tran_uops_0_xcpt_ma_if),
    .io_deq_bits_tran_uops_0_bp_debug_if(trans_buffer_io_deq_bits_tran_uops_0_bp_debug_if),
    .io_deq_bits_tran_uops_0_bp_xcpt_if(trans_buffer_io_deq_bits_tran_uops_0_bp_xcpt_if),
    .io_deq_bits_tran_uops_0_debug_fsrc(trans_buffer_io_deq_bits_tran_uops_0_debug_fsrc),
    .io_deq_bits_tran_uops_0_debug_tsrc(trans_buffer_io_deq_bits_tran_uops_0_debug_tsrc),
    .io_deq_bits_tran_uops_1_switch(trans_buffer_io_deq_bits_tran_uops_1_switch),
    .io_deq_bits_tran_uops_1_switch_off(trans_buffer_io_deq_bits_tran_uops_1_switch_off),
    .io_deq_bits_tran_uops_1_is_unicore(trans_buffer_io_deq_bits_tran_uops_1_is_unicore),
    .io_deq_bits_tran_uops_1_shift(trans_buffer_io_deq_bits_tran_uops_1_shift),
    .io_deq_bits_tran_uops_1_lrs3_rtype(trans_buffer_io_deq_bits_tran_uops_1_lrs3_rtype),
    .io_deq_bits_tran_uops_1_rflag(trans_buffer_io_deq_bits_tran_uops_1_rflag),
    .io_deq_bits_tran_uops_1_wflag(trans_buffer_io_deq_bits_tran_uops_1_wflag),
    .io_deq_bits_tran_uops_1_prflag(trans_buffer_io_deq_bits_tran_uops_1_prflag),
    .io_deq_bits_tran_uops_1_pwflag(trans_buffer_io_deq_bits_tran_uops_1_pwflag),
    .io_deq_bits_tran_uops_1_pflag_busy(trans_buffer_io_deq_bits_tran_uops_1_pflag_busy),
    .io_deq_bits_tran_uops_1_stale_pflag(trans_buffer_io_deq_bits_tran_uops_1_stale_pflag),
    .io_deq_bits_tran_uops_1_op1_sel(trans_buffer_io_deq_bits_tran_uops_1_op1_sel),
    .io_deq_bits_tran_uops_1_op2_sel(trans_buffer_io_deq_bits_tran_uops_1_op2_sel),
    .io_deq_bits_tran_uops_1_split_num(trans_buffer_io_deq_bits_tran_uops_1_split_num),
    .io_deq_bits_tran_uops_1_self_index(trans_buffer_io_deq_bits_tran_uops_1_self_index),
    .io_deq_bits_tran_uops_1_rob_inst_idx(trans_buffer_io_deq_bits_tran_uops_1_rob_inst_idx),
    .io_deq_bits_tran_uops_1_address_num(trans_buffer_io_deq_bits_tran_uops_1_address_num),
    .io_deq_bits_tran_uops_1_uopc(trans_buffer_io_deq_bits_tran_uops_1_uopc),
    .io_deq_bits_tran_uops_1_inst(trans_buffer_io_deq_bits_tran_uops_1_inst),
    .io_deq_bits_tran_uops_1_debug_inst(trans_buffer_io_deq_bits_tran_uops_1_debug_inst),
    .io_deq_bits_tran_uops_1_is_rvc(trans_buffer_io_deq_bits_tran_uops_1_is_rvc),
    .io_deq_bits_tran_uops_1_debug_pc(trans_buffer_io_deq_bits_tran_uops_1_debug_pc),
    .io_deq_bits_tran_uops_1_iq_type(trans_buffer_io_deq_bits_tran_uops_1_iq_type),
    .io_deq_bits_tran_uops_1_fu_code(trans_buffer_io_deq_bits_tran_uops_1_fu_code),
    .io_deq_bits_tran_uops_1_ctrl_br_type(trans_buffer_io_deq_bits_tran_uops_1_ctrl_br_type),
    .io_deq_bits_tran_uops_1_ctrl_op1_sel(trans_buffer_io_deq_bits_tran_uops_1_ctrl_op1_sel),
    .io_deq_bits_tran_uops_1_ctrl_op2_sel(trans_buffer_io_deq_bits_tran_uops_1_ctrl_op2_sel),
    .io_deq_bits_tran_uops_1_ctrl_imm_sel(trans_buffer_io_deq_bits_tran_uops_1_ctrl_imm_sel),
    .io_deq_bits_tran_uops_1_ctrl_op_fcn(trans_buffer_io_deq_bits_tran_uops_1_ctrl_op_fcn),
    .io_deq_bits_tran_uops_1_ctrl_fcn_dw(trans_buffer_io_deq_bits_tran_uops_1_ctrl_fcn_dw),
    .io_deq_bits_tran_uops_1_ctrl_csr_cmd(trans_buffer_io_deq_bits_tran_uops_1_ctrl_csr_cmd),
    .io_deq_bits_tran_uops_1_ctrl_is_load(trans_buffer_io_deq_bits_tran_uops_1_ctrl_is_load),
    .io_deq_bits_tran_uops_1_ctrl_is_sta(trans_buffer_io_deq_bits_tran_uops_1_ctrl_is_sta),
    .io_deq_bits_tran_uops_1_ctrl_is_std(trans_buffer_io_deq_bits_tran_uops_1_ctrl_is_std),
    .io_deq_bits_tran_uops_1_ctrl_op3_sel(trans_buffer_io_deq_bits_tran_uops_1_ctrl_op3_sel),
    .io_deq_bits_tran_uops_1_iw_state(trans_buffer_io_deq_bits_tran_uops_1_iw_state),
    .io_deq_bits_tran_uops_1_iw_p1_poisoned(trans_buffer_io_deq_bits_tran_uops_1_iw_p1_poisoned),
    .io_deq_bits_tran_uops_1_iw_p2_poisoned(trans_buffer_io_deq_bits_tran_uops_1_iw_p2_poisoned),
    .io_deq_bits_tran_uops_1_is_br(trans_buffer_io_deq_bits_tran_uops_1_is_br),
    .io_deq_bits_tran_uops_1_is_jalr(trans_buffer_io_deq_bits_tran_uops_1_is_jalr),
    .io_deq_bits_tran_uops_1_is_jal(trans_buffer_io_deq_bits_tran_uops_1_is_jal),
    .io_deq_bits_tran_uops_1_is_sfb(trans_buffer_io_deq_bits_tran_uops_1_is_sfb),
    .io_deq_bits_tran_uops_1_br_mask(trans_buffer_io_deq_bits_tran_uops_1_br_mask),
    .io_deq_bits_tran_uops_1_br_tag(trans_buffer_io_deq_bits_tran_uops_1_br_tag),
    .io_deq_bits_tran_uops_1_ftq_idx(trans_buffer_io_deq_bits_tran_uops_1_ftq_idx),
    .io_deq_bits_tran_uops_1_edge_inst(trans_buffer_io_deq_bits_tran_uops_1_edge_inst),
    .io_deq_bits_tran_uops_1_pc_lob(trans_buffer_io_deq_bits_tran_uops_1_pc_lob),
    .io_deq_bits_tran_uops_1_taken(trans_buffer_io_deq_bits_tran_uops_1_taken),
    .io_deq_bits_tran_uops_1_imm_packed(trans_buffer_io_deq_bits_tran_uops_1_imm_packed),
    .io_deq_bits_tran_uops_1_csr_addr(trans_buffer_io_deq_bits_tran_uops_1_csr_addr),
    .io_deq_bits_tran_uops_1_rob_idx(trans_buffer_io_deq_bits_tran_uops_1_rob_idx),
    .io_deq_bits_tran_uops_1_ldq_idx(trans_buffer_io_deq_bits_tran_uops_1_ldq_idx),
    .io_deq_bits_tran_uops_1_stq_idx(trans_buffer_io_deq_bits_tran_uops_1_stq_idx),
    .io_deq_bits_tran_uops_1_rxq_idx(trans_buffer_io_deq_bits_tran_uops_1_rxq_idx),
    .io_deq_bits_tran_uops_1_pdst(trans_buffer_io_deq_bits_tran_uops_1_pdst),
    .io_deq_bits_tran_uops_1_prs1(trans_buffer_io_deq_bits_tran_uops_1_prs1),
    .io_deq_bits_tran_uops_1_prs2(trans_buffer_io_deq_bits_tran_uops_1_prs2),
    .io_deq_bits_tran_uops_1_prs3(trans_buffer_io_deq_bits_tran_uops_1_prs3),
    .io_deq_bits_tran_uops_1_ppred(trans_buffer_io_deq_bits_tran_uops_1_ppred),
    .io_deq_bits_tran_uops_1_prs1_busy(trans_buffer_io_deq_bits_tran_uops_1_prs1_busy),
    .io_deq_bits_tran_uops_1_prs2_busy(trans_buffer_io_deq_bits_tran_uops_1_prs2_busy),
    .io_deq_bits_tran_uops_1_prs3_busy(trans_buffer_io_deq_bits_tran_uops_1_prs3_busy),
    .io_deq_bits_tran_uops_1_ppred_busy(trans_buffer_io_deq_bits_tran_uops_1_ppred_busy),
    .io_deq_bits_tran_uops_1_stale_pdst(trans_buffer_io_deq_bits_tran_uops_1_stale_pdst),
    .io_deq_bits_tran_uops_1_exception(trans_buffer_io_deq_bits_tran_uops_1_exception),
    .io_deq_bits_tran_uops_1_exc_cause(trans_buffer_io_deq_bits_tran_uops_1_exc_cause),
    .io_deq_bits_tran_uops_1_bypassable(trans_buffer_io_deq_bits_tran_uops_1_bypassable),
    .io_deq_bits_tran_uops_1_mem_cmd(trans_buffer_io_deq_bits_tran_uops_1_mem_cmd),
    .io_deq_bits_tran_uops_1_mem_size(trans_buffer_io_deq_bits_tran_uops_1_mem_size),
    .io_deq_bits_tran_uops_1_mem_signed(trans_buffer_io_deq_bits_tran_uops_1_mem_signed),
    .io_deq_bits_tran_uops_1_is_fence(trans_buffer_io_deq_bits_tran_uops_1_is_fence),
    .io_deq_bits_tran_uops_1_is_fencei(trans_buffer_io_deq_bits_tran_uops_1_is_fencei),
    .io_deq_bits_tran_uops_1_is_amo(trans_buffer_io_deq_bits_tran_uops_1_is_amo),
    .io_deq_bits_tran_uops_1_uses_ldq(trans_buffer_io_deq_bits_tran_uops_1_uses_ldq),
    .io_deq_bits_tran_uops_1_uses_stq(trans_buffer_io_deq_bits_tran_uops_1_uses_stq),
    .io_deq_bits_tran_uops_1_is_sys_pc2epc(trans_buffer_io_deq_bits_tran_uops_1_is_sys_pc2epc),
    .io_deq_bits_tran_uops_1_is_unique(trans_buffer_io_deq_bits_tran_uops_1_is_unique),
    .io_deq_bits_tran_uops_1_flush_on_commit(trans_buffer_io_deq_bits_tran_uops_1_flush_on_commit),
    .io_deq_bits_tran_uops_1_ldst_is_rs1(trans_buffer_io_deq_bits_tran_uops_1_ldst_is_rs1),
    .io_deq_bits_tran_uops_1_ldst(trans_buffer_io_deq_bits_tran_uops_1_ldst),
    .io_deq_bits_tran_uops_1_lrs1(trans_buffer_io_deq_bits_tran_uops_1_lrs1),
    .io_deq_bits_tran_uops_1_lrs2(trans_buffer_io_deq_bits_tran_uops_1_lrs2),
    .io_deq_bits_tran_uops_1_lrs3(trans_buffer_io_deq_bits_tran_uops_1_lrs3),
    .io_deq_bits_tran_uops_1_ldst_val(trans_buffer_io_deq_bits_tran_uops_1_ldst_val),
    .io_deq_bits_tran_uops_1_dst_rtype(trans_buffer_io_deq_bits_tran_uops_1_dst_rtype),
    .io_deq_bits_tran_uops_1_lrs1_rtype(trans_buffer_io_deq_bits_tran_uops_1_lrs1_rtype),
    .io_deq_bits_tran_uops_1_lrs2_rtype(trans_buffer_io_deq_bits_tran_uops_1_lrs2_rtype),
    .io_deq_bits_tran_uops_1_frs3_en(trans_buffer_io_deq_bits_tran_uops_1_frs3_en),
    .io_deq_bits_tran_uops_1_fp_val(trans_buffer_io_deq_bits_tran_uops_1_fp_val),
    .io_deq_bits_tran_uops_1_fp_single(trans_buffer_io_deq_bits_tran_uops_1_fp_single),
    .io_deq_bits_tran_uops_1_xcpt_pf_if(trans_buffer_io_deq_bits_tran_uops_1_xcpt_pf_if),
    .io_deq_bits_tran_uops_1_xcpt_ae_if(trans_buffer_io_deq_bits_tran_uops_1_xcpt_ae_if),
    .io_deq_bits_tran_uops_1_xcpt_ma_if(trans_buffer_io_deq_bits_tran_uops_1_xcpt_ma_if),
    .io_deq_bits_tran_uops_1_bp_debug_if(trans_buffer_io_deq_bits_tran_uops_1_bp_debug_if),
    .io_deq_bits_tran_uops_1_bp_xcpt_if(trans_buffer_io_deq_bits_tran_uops_1_bp_xcpt_if),
    .io_deq_bits_tran_uops_1_debug_fsrc(trans_buffer_io_deq_bits_tran_uops_1_debug_fsrc),
    .io_deq_bits_tran_uops_1_debug_tsrc(trans_buffer_io_deq_bits_tran_uops_1_debug_tsrc),
    .io_deq_bits_tran_valids_0(trans_buffer_io_deq_bits_tran_valids_0),
    .io_deq_bits_tran_valids_1(trans_buffer_io_deq_bits_tran_valids_1),
    .io_clear(trans_buffer_io_clear),
    .io_isUnicoreMode(trans_buffer_io_isUnicoreMode)
  );
  assign io_enq_ready = io_clear | REG & trans_buffer_io_enq_ready; // @[enq_transBuff.scala 81:30]
  assign io_deq_tran_uops_0_switch = trans_buffer_io_deq_bits_tran_uops_0_switch; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_switch_off = trans_buffer_io_deq_bits_tran_uops_0_switch_off; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_is_unicore = trans_buffer_io_deq_bits_tran_uops_0_is_unicore; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_shift = trans_buffer_io_deq_bits_tran_uops_0_shift; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_lrs3_rtype = trans_buffer_io_deq_bits_tran_uops_0_lrs3_rtype; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_rflag = trans_buffer_io_deq_bits_tran_uops_0_rflag; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_wflag = trans_buffer_io_deq_bits_tran_uops_0_wflag; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_prflag = trans_buffer_io_deq_bits_tran_uops_0_prflag; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_pwflag = trans_buffer_io_deq_bits_tran_uops_0_pwflag; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_pflag_busy = trans_buffer_io_deq_bits_tran_uops_0_pflag_busy; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_stale_pflag = trans_buffer_io_deq_bits_tran_uops_0_stale_pflag; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_op1_sel = trans_buffer_io_deq_bits_tran_uops_0_op1_sel; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_op2_sel = trans_buffer_io_deq_bits_tran_uops_0_op2_sel; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_split_num = trans_buffer_io_deq_bits_tran_uops_0_split_num; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_self_index = trans_buffer_io_deq_bits_tran_uops_0_self_index; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_rob_inst_idx = trans_buffer_io_deq_bits_tran_uops_0_rob_inst_idx; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_address_num = trans_buffer_io_deq_bits_tran_uops_0_address_num; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_uopc = trans_buffer_io_deq_bits_tran_uops_0_uopc; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_inst = trans_buffer_io_deq_bits_tran_uops_0_inst; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_debug_inst = trans_buffer_io_deq_bits_tran_uops_0_debug_inst; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_is_rvc = trans_buffer_io_deq_bits_tran_uops_0_is_rvc; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_debug_pc = trans_buffer_io_deq_bits_tran_uops_0_debug_pc; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_iq_type = trans_buffer_io_deq_bits_tran_uops_0_iq_type; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_fu_code = trans_buffer_io_deq_bits_tran_uops_0_fu_code; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_ctrl_br_type = trans_buffer_io_deq_bits_tran_uops_0_ctrl_br_type; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_ctrl_op1_sel = trans_buffer_io_deq_bits_tran_uops_0_ctrl_op1_sel; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_ctrl_op2_sel = trans_buffer_io_deq_bits_tran_uops_0_ctrl_op2_sel; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_ctrl_imm_sel = trans_buffer_io_deq_bits_tran_uops_0_ctrl_imm_sel; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_ctrl_op_fcn = trans_buffer_io_deq_bits_tran_uops_0_ctrl_op_fcn; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_ctrl_fcn_dw = trans_buffer_io_deq_bits_tran_uops_0_ctrl_fcn_dw; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_ctrl_csr_cmd = trans_buffer_io_deq_bits_tran_uops_0_ctrl_csr_cmd; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_ctrl_is_load = trans_buffer_io_deq_bits_tran_uops_0_ctrl_is_load; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_ctrl_is_sta = trans_buffer_io_deq_bits_tran_uops_0_ctrl_is_sta; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_ctrl_is_std = trans_buffer_io_deq_bits_tran_uops_0_ctrl_is_std; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_ctrl_op3_sel = trans_buffer_io_deq_bits_tran_uops_0_ctrl_op3_sel; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_iw_state = trans_buffer_io_deq_bits_tran_uops_0_iw_state; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_iw_p1_poisoned = trans_buffer_io_deq_bits_tran_uops_0_iw_p1_poisoned; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_iw_p2_poisoned = trans_buffer_io_deq_bits_tran_uops_0_iw_p2_poisoned; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_is_br = trans_buffer_io_deq_bits_tran_uops_0_is_br; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_is_jalr = trans_buffer_io_deq_bits_tran_uops_0_is_jalr; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_is_jal = trans_buffer_io_deq_bits_tran_uops_0_is_jal; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_is_sfb = trans_buffer_io_deq_bits_tran_uops_0_is_sfb; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_br_mask = trans_buffer_io_deq_bits_tran_uops_0_br_mask; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_br_tag = trans_buffer_io_deq_bits_tran_uops_0_br_tag; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_ftq_idx = trans_buffer_io_deq_bits_tran_uops_0_ftq_idx; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_edge_inst = trans_buffer_io_deq_bits_tran_uops_0_edge_inst; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_pc_lob = trans_buffer_io_deq_bits_tran_uops_0_pc_lob; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_taken = trans_buffer_io_deq_bits_tran_uops_0_taken; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_imm_packed = trans_buffer_io_deq_bits_tran_uops_0_imm_packed; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_csr_addr = trans_buffer_io_deq_bits_tran_uops_0_csr_addr; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_rob_idx = trans_buffer_io_deq_bits_tran_uops_0_rob_idx; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_ldq_idx = trans_buffer_io_deq_bits_tran_uops_0_ldq_idx; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_stq_idx = trans_buffer_io_deq_bits_tran_uops_0_stq_idx; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_rxq_idx = trans_buffer_io_deq_bits_tran_uops_0_rxq_idx; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_pdst = trans_buffer_io_deq_bits_tran_uops_0_pdst; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_prs1 = trans_buffer_io_deq_bits_tran_uops_0_prs1; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_prs2 = trans_buffer_io_deq_bits_tran_uops_0_prs2; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_prs3 = trans_buffer_io_deq_bits_tran_uops_0_prs3; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_ppred = trans_buffer_io_deq_bits_tran_uops_0_ppred; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_prs1_busy = trans_buffer_io_deq_bits_tran_uops_0_prs1_busy; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_prs2_busy = trans_buffer_io_deq_bits_tran_uops_0_prs2_busy; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_prs3_busy = trans_buffer_io_deq_bits_tran_uops_0_prs3_busy; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_ppred_busy = trans_buffer_io_deq_bits_tran_uops_0_ppred_busy; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_stale_pdst = trans_buffer_io_deq_bits_tran_uops_0_stale_pdst; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_exception = trans_buffer_io_deq_bits_tran_uops_0_exception; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_exc_cause = trans_buffer_io_deq_bits_tran_uops_0_exc_cause; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_bypassable = trans_buffer_io_deq_bits_tran_uops_0_bypassable; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_mem_cmd = trans_buffer_io_deq_bits_tran_uops_0_mem_cmd; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_mem_size = trans_buffer_io_deq_bits_tran_uops_0_mem_size; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_mem_signed = trans_buffer_io_deq_bits_tran_uops_0_mem_signed; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_is_fence = trans_buffer_io_deq_bits_tran_uops_0_is_fence; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_is_fencei = trans_buffer_io_deq_bits_tran_uops_0_is_fencei; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_is_amo = trans_buffer_io_deq_bits_tran_uops_0_is_amo; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_uses_ldq = trans_buffer_io_deq_bits_tran_uops_0_uses_ldq; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_uses_stq = trans_buffer_io_deq_bits_tran_uops_0_uses_stq; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_is_sys_pc2epc = trans_buffer_io_deq_bits_tran_uops_0_is_sys_pc2epc; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_is_unique = trans_buffer_io_deq_bits_tran_uops_0_is_unique; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_flush_on_commit = trans_buffer_io_deq_bits_tran_uops_0_flush_on_commit; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_ldst_is_rs1 = trans_buffer_io_deq_bits_tran_uops_0_ldst_is_rs1; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_ldst = trans_buffer_io_deq_bits_tran_uops_0_ldst; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_lrs1 = trans_buffer_io_deq_bits_tran_uops_0_lrs1; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_lrs2 = trans_buffer_io_deq_bits_tran_uops_0_lrs2; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_lrs3 = trans_buffer_io_deq_bits_tran_uops_0_lrs3; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_ldst_val = trans_buffer_io_deq_bits_tran_uops_0_ldst_val; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_dst_rtype = trans_buffer_io_deq_bits_tran_uops_0_dst_rtype; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_lrs1_rtype = trans_buffer_io_deq_bits_tran_uops_0_lrs1_rtype; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_lrs2_rtype = trans_buffer_io_deq_bits_tran_uops_0_lrs2_rtype; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_frs3_en = trans_buffer_io_deq_bits_tran_uops_0_frs3_en; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_fp_val = trans_buffer_io_deq_bits_tran_uops_0_fp_val; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_fp_single = trans_buffer_io_deq_bits_tran_uops_0_fp_single; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_xcpt_pf_if = trans_buffer_io_deq_bits_tran_uops_0_xcpt_pf_if; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_xcpt_ae_if = trans_buffer_io_deq_bits_tran_uops_0_xcpt_ae_if; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_xcpt_ma_if = trans_buffer_io_deq_bits_tran_uops_0_xcpt_ma_if; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_bp_debug_if = trans_buffer_io_deq_bits_tran_uops_0_bp_debug_if; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_bp_xcpt_if = trans_buffer_io_deq_bits_tran_uops_0_bp_xcpt_if; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_debug_fsrc = trans_buffer_io_deq_bits_tran_uops_0_debug_fsrc; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_0_debug_tsrc = trans_buffer_io_deq_bits_tran_uops_0_debug_tsrc; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_switch = trans_buffer_io_deq_bits_tran_uops_1_switch; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_switch_off = trans_buffer_io_deq_bits_tran_uops_1_switch_off; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_is_unicore = trans_buffer_io_deq_bits_tran_uops_1_is_unicore; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_shift = trans_buffer_io_deq_bits_tran_uops_1_shift; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_lrs3_rtype = trans_buffer_io_deq_bits_tran_uops_1_lrs3_rtype; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_rflag = trans_buffer_io_deq_bits_tran_uops_1_rflag; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_wflag = trans_buffer_io_deq_bits_tran_uops_1_wflag; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_prflag = trans_buffer_io_deq_bits_tran_uops_1_prflag; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_pwflag = trans_buffer_io_deq_bits_tran_uops_1_pwflag; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_pflag_busy = trans_buffer_io_deq_bits_tran_uops_1_pflag_busy; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_stale_pflag = trans_buffer_io_deq_bits_tran_uops_1_stale_pflag; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_op1_sel = trans_buffer_io_deq_bits_tran_uops_1_op1_sel; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_op2_sel = trans_buffer_io_deq_bits_tran_uops_1_op2_sel; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_split_num = trans_buffer_io_deq_bits_tran_uops_1_split_num; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_self_index = trans_buffer_io_deq_bits_tran_uops_1_self_index; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_rob_inst_idx = trans_buffer_io_deq_bits_tran_uops_1_rob_inst_idx; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_address_num = trans_buffer_io_deq_bits_tran_uops_1_address_num; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_uopc = trans_buffer_io_deq_bits_tran_uops_1_uopc; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_inst = trans_buffer_io_deq_bits_tran_uops_1_inst; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_debug_inst = trans_buffer_io_deq_bits_tran_uops_1_debug_inst; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_is_rvc = trans_buffer_io_deq_bits_tran_uops_1_is_rvc; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_debug_pc = trans_buffer_io_deq_bits_tran_uops_1_debug_pc; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_iq_type = trans_buffer_io_deq_bits_tran_uops_1_iq_type; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_fu_code = trans_buffer_io_deq_bits_tran_uops_1_fu_code; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_ctrl_br_type = trans_buffer_io_deq_bits_tran_uops_1_ctrl_br_type; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_ctrl_op1_sel = trans_buffer_io_deq_bits_tran_uops_1_ctrl_op1_sel; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_ctrl_op2_sel = trans_buffer_io_deq_bits_tran_uops_1_ctrl_op2_sel; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_ctrl_imm_sel = trans_buffer_io_deq_bits_tran_uops_1_ctrl_imm_sel; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_ctrl_op_fcn = trans_buffer_io_deq_bits_tran_uops_1_ctrl_op_fcn; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_ctrl_fcn_dw = trans_buffer_io_deq_bits_tran_uops_1_ctrl_fcn_dw; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_ctrl_csr_cmd = trans_buffer_io_deq_bits_tran_uops_1_ctrl_csr_cmd; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_ctrl_is_load = trans_buffer_io_deq_bits_tran_uops_1_ctrl_is_load; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_ctrl_is_sta = trans_buffer_io_deq_bits_tran_uops_1_ctrl_is_sta; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_ctrl_is_std = trans_buffer_io_deq_bits_tran_uops_1_ctrl_is_std; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_ctrl_op3_sel = trans_buffer_io_deq_bits_tran_uops_1_ctrl_op3_sel; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_iw_state = trans_buffer_io_deq_bits_tran_uops_1_iw_state; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_iw_p1_poisoned = trans_buffer_io_deq_bits_tran_uops_1_iw_p1_poisoned; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_iw_p2_poisoned = trans_buffer_io_deq_bits_tran_uops_1_iw_p2_poisoned; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_is_br = trans_buffer_io_deq_bits_tran_uops_1_is_br; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_is_jalr = trans_buffer_io_deq_bits_tran_uops_1_is_jalr; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_is_jal = trans_buffer_io_deq_bits_tran_uops_1_is_jal; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_is_sfb = trans_buffer_io_deq_bits_tran_uops_1_is_sfb; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_br_mask = trans_buffer_io_deq_bits_tran_uops_1_br_mask; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_br_tag = trans_buffer_io_deq_bits_tran_uops_1_br_tag; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_ftq_idx = trans_buffer_io_deq_bits_tran_uops_1_ftq_idx; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_edge_inst = trans_buffer_io_deq_bits_tran_uops_1_edge_inst; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_pc_lob = trans_buffer_io_deq_bits_tran_uops_1_pc_lob; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_taken = trans_buffer_io_deq_bits_tran_uops_1_taken; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_imm_packed = trans_buffer_io_deq_bits_tran_uops_1_imm_packed; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_csr_addr = trans_buffer_io_deq_bits_tran_uops_1_csr_addr; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_rob_idx = trans_buffer_io_deq_bits_tran_uops_1_rob_idx; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_ldq_idx = trans_buffer_io_deq_bits_tran_uops_1_ldq_idx; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_stq_idx = trans_buffer_io_deq_bits_tran_uops_1_stq_idx; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_rxq_idx = trans_buffer_io_deq_bits_tran_uops_1_rxq_idx; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_pdst = trans_buffer_io_deq_bits_tran_uops_1_pdst; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_prs1 = trans_buffer_io_deq_bits_tran_uops_1_prs1; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_prs2 = trans_buffer_io_deq_bits_tran_uops_1_prs2; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_prs3 = trans_buffer_io_deq_bits_tran_uops_1_prs3; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_ppred = trans_buffer_io_deq_bits_tran_uops_1_ppred; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_prs1_busy = trans_buffer_io_deq_bits_tran_uops_1_prs1_busy; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_prs2_busy = trans_buffer_io_deq_bits_tran_uops_1_prs2_busy; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_prs3_busy = trans_buffer_io_deq_bits_tran_uops_1_prs3_busy; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_ppred_busy = trans_buffer_io_deq_bits_tran_uops_1_ppred_busy; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_stale_pdst = trans_buffer_io_deq_bits_tran_uops_1_stale_pdst; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_exception = trans_buffer_io_deq_bits_tran_uops_1_exception; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_exc_cause = trans_buffer_io_deq_bits_tran_uops_1_exc_cause; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_bypassable = trans_buffer_io_deq_bits_tran_uops_1_bypassable; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_mem_cmd = trans_buffer_io_deq_bits_tran_uops_1_mem_cmd; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_mem_size = trans_buffer_io_deq_bits_tran_uops_1_mem_size; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_mem_signed = trans_buffer_io_deq_bits_tran_uops_1_mem_signed; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_is_fence = trans_buffer_io_deq_bits_tran_uops_1_is_fence; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_is_fencei = trans_buffer_io_deq_bits_tran_uops_1_is_fencei; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_is_amo = trans_buffer_io_deq_bits_tran_uops_1_is_amo; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_uses_ldq = trans_buffer_io_deq_bits_tran_uops_1_uses_ldq; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_uses_stq = trans_buffer_io_deq_bits_tran_uops_1_uses_stq; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_is_sys_pc2epc = trans_buffer_io_deq_bits_tran_uops_1_is_sys_pc2epc; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_is_unique = trans_buffer_io_deq_bits_tran_uops_1_is_unique; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_flush_on_commit = trans_buffer_io_deq_bits_tran_uops_1_flush_on_commit; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_ldst_is_rs1 = trans_buffer_io_deq_bits_tran_uops_1_ldst_is_rs1; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_ldst = trans_buffer_io_deq_bits_tran_uops_1_ldst; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_lrs1 = trans_buffer_io_deq_bits_tran_uops_1_lrs1; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_lrs2 = trans_buffer_io_deq_bits_tran_uops_1_lrs2; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_lrs3 = trans_buffer_io_deq_bits_tran_uops_1_lrs3; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_ldst_val = trans_buffer_io_deq_bits_tran_uops_1_ldst_val; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_dst_rtype = trans_buffer_io_deq_bits_tran_uops_1_dst_rtype; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_lrs1_rtype = trans_buffer_io_deq_bits_tran_uops_1_lrs1_rtype; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_lrs2_rtype = trans_buffer_io_deq_bits_tran_uops_1_lrs2_rtype; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_frs3_en = trans_buffer_io_deq_bits_tran_uops_1_frs3_en; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_fp_val = trans_buffer_io_deq_bits_tran_uops_1_fp_val; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_fp_single = trans_buffer_io_deq_bits_tran_uops_1_fp_single; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_xcpt_pf_if = trans_buffer_io_deq_bits_tran_uops_1_xcpt_pf_if; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_xcpt_ae_if = trans_buffer_io_deq_bits_tran_uops_1_xcpt_ae_if; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_xcpt_ma_if = trans_buffer_io_deq_bits_tran_uops_1_xcpt_ma_if; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_bp_debug_if = trans_buffer_io_deq_bits_tran_uops_1_bp_debug_if; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_bp_xcpt_if = trans_buffer_io_deq_bits_tran_uops_1_bp_xcpt_if; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_debug_fsrc = trans_buffer_io_deq_bits_tran_uops_1_debug_fsrc; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_uops_1_debug_tsrc = trans_buffer_io_deq_bits_tran_uops_1_debug_tsrc; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_valids_0 = trans_buffer_io_deq_bits_tran_valids_0; // @[enq_transBuff.scala 46:12]
  assign io_deq_tran_valids_1 = trans_buffer_io_deq_bits_tran_valids_1; // @[enq_transBuff.scala 46:12]
  assign io_deq_valid = trans_buffer_io_deq_valid; // @[enq_transBuff.scala 45:18]
  assign trans_buffer_clock = clock;
  assign trans_buffer_reset = reset;
  assign trans_buffer_io_enq_valid = _T ? io_enq_valid : enq_valid; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 127:35 enq_transBuff.scala 131:35]
  assign trans_buffer_io_enq_bits_dec_uops_0_switch = _T ? io_enq_0_dec_uops_0_switch : _GEN_3950; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_switch_off = _T ? io_enq_0_dec_uops_0_switch_off : _GEN_3942; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_is_unicore = _T ? io_enq_0_dec_uops_0_is_unicore : _GEN_3934; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_shift = _T ? io_enq_0_dec_uops_0_shift : _GEN_3926; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_lrs3_rtype = _T ? io_enq_0_dec_uops_0_lrs3_rtype : _GEN_3918; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_rflag = _T ? io_enq_0_dec_uops_0_rflag : _GEN_3910; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_wflag = _T ? io_enq_0_dec_uops_0_wflag : _GEN_3902; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_prflag = _T ? io_enq_0_dec_uops_0_prflag : _GEN_3894; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_pwflag = _T ? io_enq_0_dec_uops_0_pwflag : _GEN_3886; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_pflag_busy = _T ? io_enq_0_dec_uops_0_pflag_busy : _GEN_3878; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_stale_pflag = _T ? io_enq_0_dec_uops_0_stale_pflag : _GEN_3870; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_op1_sel = _T ? io_enq_0_dec_uops_0_op1_sel : _GEN_3862; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_op2_sel = _T ? io_enq_0_dec_uops_0_op2_sel : _GEN_3854; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_split_num = _T ? io_enq_0_dec_uops_0_split_num : _GEN_3846; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_self_index = _T ? io_enq_0_dec_uops_0_self_index : _GEN_3838; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_rob_inst_idx = _T ? io_enq_0_dec_uops_0_rob_inst_idx : _GEN_3830; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_address_num = _T ? io_enq_0_dec_uops_0_address_num : _GEN_3822; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_uopc = _T ? io_enq_0_dec_uops_0_uopc : _GEN_3814; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_inst = _T ? io_enq_0_dec_uops_0_inst : _GEN_3806; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_debug_inst = _T ? io_enq_0_dec_uops_0_debug_inst : _GEN_3798; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_is_rvc = _T ? io_enq_0_dec_uops_0_is_rvc : _GEN_3790; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_debug_pc = _T ? io_enq_0_dec_uops_0_debug_pc : _GEN_3782; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_iq_type = _T ? io_enq_0_dec_uops_0_iq_type : _GEN_3774; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_fu_code = _T ? io_enq_0_dec_uops_0_fu_code : _GEN_3766; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_ctrl_br_type = _T ? io_enq_0_dec_uops_0_ctrl_br_type : _GEN_3758; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_ctrl_op1_sel = _T ? io_enq_0_dec_uops_0_ctrl_op1_sel : _GEN_3750; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_ctrl_op2_sel = _T ? io_enq_0_dec_uops_0_ctrl_op2_sel : _GEN_3742; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_ctrl_imm_sel = _T ? io_enq_0_dec_uops_0_ctrl_imm_sel : _GEN_3734; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_ctrl_op_fcn = _T ? io_enq_0_dec_uops_0_ctrl_op_fcn : _GEN_3726; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_ctrl_fcn_dw = _T ? io_enq_0_dec_uops_0_ctrl_fcn_dw : _GEN_3718; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_ctrl_csr_cmd = _T ? io_enq_0_dec_uops_0_ctrl_csr_cmd : _GEN_3710; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_ctrl_is_load = _T ? io_enq_0_dec_uops_0_ctrl_is_load : _GEN_3702; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_ctrl_is_sta = _T ? io_enq_0_dec_uops_0_ctrl_is_sta : _GEN_3694; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_ctrl_is_std = _T ? io_enq_0_dec_uops_0_ctrl_is_std : _GEN_3686; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_ctrl_op3_sel = _T ? io_enq_0_dec_uops_0_ctrl_op3_sel : _GEN_3678; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_iw_state = _T ? io_enq_0_dec_uops_0_iw_state : _GEN_3670; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_iw_p1_poisoned = _T ? io_enq_0_dec_uops_0_iw_p1_poisoned : _GEN_3662; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_iw_p2_poisoned = _T ? io_enq_0_dec_uops_0_iw_p2_poisoned : _GEN_3654; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_is_br = _T ? io_enq_0_dec_uops_0_is_br : _GEN_3646; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_is_jalr = _T ? io_enq_0_dec_uops_0_is_jalr : _GEN_3638; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_is_jal = _T ? io_enq_0_dec_uops_0_is_jal : _GEN_3630; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_is_sfb = _T ? io_enq_0_dec_uops_0_is_sfb : _GEN_3622; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_br_mask = _T ? io_enq_0_dec_uops_0_br_mask : _GEN_3614; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_br_tag = _T ? io_enq_0_dec_uops_0_br_tag : _GEN_3606; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_ftq_idx = _T ? io_enq_0_dec_uops_0_ftq_idx : _GEN_3598; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_edge_inst = _T ? io_enq_0_dec_uops_0_edge_inst : _GEN_3590; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_pc_lob = _T ? io_enq_0_dec_uops_0_pc_lob : _GEN_3582; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_taken = _T ? io_enq_0_dec_uops_0_taken : _GEN_3574; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_imm_packed = _T ? io_enq_0_dec_uops_0_imm_packed : _GEN_3566; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_csr_addr = _T ? io_enq_0_dec_uops_0_csr_addr : _GEN_3558; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_rob_idx = _T ? io_enq_0_dec_uops_0_rob_idx : _GEN_3550; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_ldq_idx = _T ? io_enq_0_dec_uops_0_ldq_idx : _GEN_3542; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_stq_idx = _T ? io_enq_0_dec_uops_0_stq_idx : _GEN_3534; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_rxq_idx = _T ? io_enq_0_dec_uops_0_rxq_idx : _GEN_3526; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_pdst = _T ? io_enq_0_dec_uops_0_pdst : _GEN_3518; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_prs1 = _T ? io_enq_0_dec_uops_0_prs1 : _GEN_3510; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_prs2 = _T ? io_enq_0_dec_uops_0_prs2 : _GEN_3502; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_prs3 = _T ? io_enq_0_dec_uops_0_prs3 : _GEN_3494; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_ppred = _T ? io_enq_0_dec_uops_0_ppred : _GEN_3486; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_prs1_busy = _T ? io_enq_0_dec_uops_0_prs1_busy : _GEN_3478; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_prs2_busy = _T ? io_enq_0_dec_uops_0_prs2_busy : _GEN_3470; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_prs3_busy = _T ? io_enq_0_dec_uops_0_prs3_busy : _GEN_3462; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_ppred_busy = _T ? io_enq_0_dec_uops_0_ppred_busy : _GEN_3454; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_stale_pdst = _T ? io_enq_0_dec_uops_0_stale_pdst : _GEN_3446; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_exception = _T ? io_enq_0_dec_uops_0_exception : _GEN_3438; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_exc_cause = _T ? io_enq_0_dec_uops_0_exc_cause : _GEN_3430; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_bypassable = _T ? io_enq_0_dec_uops_0_bypassable : _GEN_3422; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_mem_cmd = _T ? io_enq_0_dec_uops_0_mem_cmd : _GEN_3414; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_mem_size = _T ? io_enq_0_dec_uops_0_mem_size : _GEN_3406; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_mem_signed = _T ? io_enq_0_dec_uops_0_mem_signed : _GEN_3398; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_is_fence = _T ? io_enq_0_dec_uops_0_is_fence : _GEN_3390; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_is_fencei = _T ? io_enq_0_dec_uops_0_is_fencei : _GEN_3382; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_is_amo = _T ? io_enq_0_dec_uops_0_is_amo : _GEN_3374; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_uses_ldq = _T ? io_enq_0_dec_uops_0_uses_ldq : _GEN_3366; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_uses_stq = _T ? io_enq_0_dec_uops_0_uses_stq : _GEN_3358; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_is_sys_pc2epc = _T ? io_enq_0_dec_uops_0_is_sys_pc2epc : _GEN_3350; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_is_unique = _T ? io_enq_0_dec_uops_0_is_unique : _GEN_3342; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_flush_on_commit = _T ? io_enq_0_dec_uops_0_flush_on_commit : _GEN_3334; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_ldst_is_rs1 = _T ? io_enq_0_dec_uops_0_ldst_is_rs1 : _GEN_3326; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_ldst = _T ? io_enq_0_dec_uops_0_ldst : _GEN_3318; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_lrs1 = _T ? io_enq_0_dec_uops_0_lrs1 : _GEN_3310; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_lrs2 = _T ? io_enq_0_dec_uops_0_lrs2 : _GEN_3302; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_lrs3 = _T ? io_enq_0_dec_uops_0_lrs3 : _GEN_3294; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_ldst_val = _T ? io_enq_0_dec_uops_0_ldst_val : _GEN_3286; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_dst_rtype = _T ? io_enq_0_dec_uops_0_dst_rtype : _GEN_3278; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_lrs1_rtype = _T ? io_enq_0_dec_uops_0_lrs1_rtype : _GEN_3270; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_lrs2_rtype = _T ? io_enq_0_dec_uops_0_lrs2_rtype : _GEN_3262; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_frs3_en = _T ? io_enq_0_dec_uops_0_frs3_en : _GEN_3254; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_fp_val = _T ? io_enq_0_dec_uops_0_fp_val : _GEN_3246; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_fp_single = _T ? io_enq_0_dec_uops_0_fp_single : _GEN_3238; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_xcpt_pf_if = _T ? io_enq_0_dec_uops_0_xcpt_pf_if : _GEN_3230; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_xcpt_ae_if = _T ? io_enq_0_dec_uops_0_xcpt_ae_if : _GEN_3222; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_xcpt_ma_if = _T ? io_enq_0_dec_uops_0_xcpt_ma_if : _GEN_3214; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_bp_debug_if = _T ? io_enq_0_dec_uops_0_bp_debug_if : _GEN_3206; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_bp_xcpt_if = _T ? io_enq_0_dec_uops_0_bp_xcpt_if : _GEN_3198; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_debug_fsrc = _T ? io_enq_0_dec_uops_0_debug_fsrc : _GEN_3190; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_0_debug_tsrc = _T ? io_enq_0_dec_uops_0_debug_tsrc : _GEN_3182; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_switch = _T ? io_enq_0_dec_uops_1_switch : _GEN_4726; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_switch_off = _T ? io_enq_0_dec_uops_1_switch_off : _GEN_4718; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_is_unicore = _T ? io_enq_0_dec_uops_1_is_unicore : _GEN_4710; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_shift = _T ? io_enq_0_dec_uops_1_shift : _GEN_4702; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_lrs3_rtype = _T ? io_enq_0_dec_uops_1_lrs3_rtype : _GEN_4694; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_rflag = _T ? io_enq_0_dec_uops_1_rflag : _GEN_4686; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_wflag = _T ? io_enq_0_dec_uops_1_wflag : _GEN_4678; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_prflag = _T ? io_enq_0_dec_uops_1_prflag : _GEN_4670; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_pwflag = _T ? io_enq_0_dec_uops_1_pwflag : _GEN_4662; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_pflag_busy = _T ? io_enq_0_dec_uops_1_pflag_busy : _GEN_4654; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_stale_pflag = _T ? io_enq_0_dec_uops_1_stale_pflag : _GEN_4646; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_op1_sel = _T ? io_enq_0_dec_uops_1_op1_sel : _GEN_4638; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_op2_sel = _T ? io_enq_0_dec_uops_1_op2_sel : _GEN_4630; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_split_num = _T ? io_enq_0_dec_uops_1_split_num : _GEN_4622; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_self_index = _T ? io_enq_0_dec_uops_1_self_index : _GEN_4614; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_rob_inst_idx = _T ? io_enq_0_dec_uops_1_rob_inst_idx : _GEN_4606; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_address_num = _T ? io_enq_0_dec_uops_1_address_num : _GEN_4598; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_uopc = _T ? io_enq_0_dec_uops_1_uopc : _GEN_4590; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_inst = _T ? io_enq_0_dec_uops_1_inst : _GEN_4582; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_debug_inst = _T ? io_enq_0_dec_uops_1_debug_inst : _GEN_4574; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_is_rvc = _T ? io_enq_0_dec_uops_1_is_rvc : _GEN_4566; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_debug_pc = _T ? io_enq_0_dec_uops_1_debug_pc : _GEN_4558; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_iq_type = _T ? io_enq_0_dec_uops_1_iq_type : _GEN_4550; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_fu_code = _T ? io_enq_0_dec_uops_1_fu_code : _GEN_4542; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_ctrl_br_type = _T ? io_enq_0_dec_uops_1_ctrl_br_type : _GEN_4534; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_ctrl_op1_sel = _T ? io_enq_0_dec_uops_1_ctrl_op1_sel : _GEN_4526; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_ctrl_op2_sel = _T ? io_enq_0_dec_uops_1_ctrl_op2_sel : _GEN_4518; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_ctrl_imm_sel = _T ? io_enq_0_dec_uops_1_ctrl_imm_sel : _GEN_4510; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_ctrl_op_fcn = _T ? io_enq_0_dec_uops_1_ctrl_op_fcn : _GEN_4502; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_ctrl_fcn_dw = _T ? io_enq_0_dec_uops_1_ctrl_fcn_dw : _GEN_4494; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_ctrl_csr_cmd = _T ? io_enq_0_dec_uops_1_ctrl_csr_cmd : _GEN_4486; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_ctrl_is_load = _T ? io_enq_0_dec_uops_1_ctrl_is_load : _GEN_4478; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_ctrl_is_sta = _T ? io_enq_0_dec_uops_1_ctrl_is_sta : _GEN_4470; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_ctrl_is_std = _T ? io_enq_0_dec_uops_1_ctrl_is_std : _GEN_4462; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_ctrl_op3_sel = _T ? io_enq_0_dec_uops_1_ctrl_op3_sel : _GEN_4454; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_iw_state = _T ? io_enq_0_dec_uops_1_iw_state : _GEN_4446; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_iw_p1_poisoned = _T ? io_enq_0_dec_uops_1_iw_p1_poisoned : _GEN_4438; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_iw_p2_poisoned = _T ? io_enq_0_dec_uops_1_iw_p2_poisoned : _GEN_4430; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_is_br = _T ? io_enq_0_dec_uops_1_is_br : _GEN_4422; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_is_jalr = _T ? io_enq_0_dec_uops_1_is_jalr : _GEN_4414; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_is_jal = _T ? io_enq_0_dec_uops_1_is_jal : _GEN_4406; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_is_sfb = _T ? io_enq_0_dec_uops_1_is_sfb : _GEN_4398; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_br_mask = _T ? io_enq_0_dec_uops_1_br_mask : _GEN_4390; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_br_tag = _T ? io_enq_0_dec_uops_1_br_tag : _GEN_4382; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_ftq_idx = _T ? io_enq_0_dec_uops_1_ftq_idx : _GEN_4374; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_edge_inst = _T ? io_enq_0_dec_uops_1_edge_inst : _GEN_4366; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_pc_lob = _T ? io_enq_0_dec_uops_1_pc_lob : _GEN_4358; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_taken = _T ? io_enq_0_dec_uops_1_taken : _GEN_4350; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_imm_packed = _T ? io_enq_0_dec_uops_1_imm_packed : _GEN_4342; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_csr_addr = _T ? io_enq_0_dec_uops_1_csr_addr : _GEN_4334; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_rob_idx = _T ? io_enq_0_dec_uops_1_rob_idx : _GEN_4326; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_ldq_idx = _T ? io_enq_0_dec_uops_1_ldq_idx : _GEN_4318; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_stq_idx = _T ? io_enq_0_dec_uops_1_stq_idx : _GEN_4310; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_rxq_idx = _T ? io_enq_0_dec_uops_1_rxq_idx : _GEN_4302; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_pdst = _T ? io_enq_0_dec_uops_1_pdst : _GEN_4294; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_prs1 = _T ? io_enq_0_dec_uops_1_prs1 : _GEN_4286; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_prs2 = _T ? io_enq_0_dec_uops_1_prs2 : _GEN_4278; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_prs3 = _T ? io_enq_0_dec_uops_1_prs3 : _GEN_4270; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_ppred = _T ? io_enq_0_dec_uops_1_ppred : _GEN_4262; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_prs1_busy = _T ? io_enq_0_dec_uops_1_prs1_busy : _GEN_4254; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_prs2_busy = _T ? io_enq_0_dec_uops_1_prs2_busy : _GEN_4246; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_prs3_busy = _T ? io_enq_0_dec_uops_1_prs3_busy : _GEN_4238; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_ppred_busy = _T ? io_enq_0_dec_uops_1_ppred_busy : _GEN_4230; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_stale_pdst = _T ? io_enq_0_dec_uops_1_stale_pdst : _GEN_4222; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_exception = _T ? io_enq_0_dec_uops_1_exception : _GEN_4214; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_exc_cause = _T ? io_enq_0_dec_uops_1_exc_cause : _GEN_4206; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_bypassable = _T ? io_enq_0_dec_uops_1_bypassable : _GEN_4198; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_mem_cmd = _T ? io_enq_0_dec_uops_1_mem_cmd : _GEN_4190; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_mem_size = _T ? io_enq_0_dec_uops_1_mem_size : _GEN_4182; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_mem_signed = _T ? io_enq_0_dec_uops_1_mem_signed : _GEN_4174; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_is_fence = _T ? io_enq_0_dec_uops_1_is_fence : _GEN_4166; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_is_fencei = _T ? io_enq_0_dec_uops_1_is_fencei : _GEN_4158; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_is_amo = _T ? io_enq_0_dec_uops_1_is_amo : _GEN_4150; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_uses_ldq = _T ? io_enq_0_dec_uops_1_uses_ldq : _GEN_4142; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_uses_stq = _T ? io_enq_0_dec_uops_1_uses_stq : _GEN_4134; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_is_sys_pc2epc = _T ? io_enq_0_dec_uops_1_is_sys_pc2epc : _GEN_4126; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_is_unique = _T ? io_enq_0_dec_uops_1_is_unique : _GEN_4118; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_flush_on_commit = _T ? io_enq_0_dec_uops_1_flush_on_commit : _GEN_4110; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_ldst_is_rs1 = _T ? io_enq_0_dec_uops_1_ldst_is_rs1 : _GEN_4102; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_ldst = _T ? io_enq_0_dec_uops_1_ldst : _GEN_4094; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_lrs1 = _T ? io_enq_0_dec_uops_1_lrs1 : _GEN_4086; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_lrs2 = _T ? io_enq_0_dec_uops_1_lrs2 : _GEN_4078; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_lrs3 = _T ? io_enq_0_dec_uops_1_lrs3 : _GEN_4070; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_ldst_val = _T ? io_enq_0_dec_uops_1_ldst_val : _GEN_4062; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_dst_rtype = _T ? io_enq_0_dec_uops_1_dst_rtype : _GEN_4054; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_lrs1_rtype = _T ? io_enq_0_dec_uops_1_lrs1_rtype : _GEN_4046; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_lrs2_rtype = _T ? io_enq_0_dec_uops_1_lrs2_rtype : _GEN_4038; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_frs3_en = _T ? io_enq_0_dec_uops_1_frs3_en : _GEN_4030; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_fp_val = _T ? io_enq_0_dec_uops_1_fp_val : _GEN_4022; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_fp_single = _T ? io_enq_0_dec_uops_1_fp_single : _GEN_4014; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_xcpt_pf_if = _T ? io_enq_0_dec_uops_1_xcpt_pf_if : _GEN_4006; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_xcpt_ae_if = _T ? io_enq_0_dec_uops_1_xcpt_ae_if : _GEN_3998; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_xcpt_ma_if = _T ? io_enq_0_dec_uops_1_xcpt_ma_if : _GEN_3990; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_bp_debug_if = _T ? io_enq_0_dec_uops_1_bp_debug_if : _GEN_3982; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_bp_xcpt_if = _T ? io_enq_0_dec_uops_1_bp_xcpt_if : _GEN_3974; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_debug_fsrc = _T ? io_enq_0_dec_uops_1_debug_fsrc : _GEN_3966; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_1_debug_tsrc = _T ? io_enq_0_dec_uops_1_debug_tsrc : _GEN_3958; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_switch = _T ? io_enq_0_dec_uops_2_switch : _GEN_5502; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_switch_off = _T ? io_enq_0_dec_uops_2_switch_off : _GEN_5494; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_is_unicore = _T ? io_enq_0_dec_uops_2_is_unicore : _GEN_5486; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_shift = _T ? io_enq_0_dec_uops_2_shift : _GEN_5478; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_lrs3_rtype = _T ? io_enq_0_dec_uops_2_lrs3_rtype : _GEN_5470; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_rflag = _T ? io_enq_0_dec_uops_2_rflag : _GEN_5462; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_wflag = _T ? io_enq_0_dec_uops_2_wflag : _GEN_5454; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_prflag = _T ? io_enq_0_dec_uops_2_prflag : _GEN_5446; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_pwflag = _T ? io_enq_0_dec_uops_2_pwflag : _GEN_5438; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_pflag_busy = _T ? io_enq_0_dec_uops_2_pflag_busy : _GEN_5430; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_stale_pflag = _T ? io_enq_0_dec_uops_2_stale_pflag : _GEN_5422; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_op1_sel = _T ? io_enq_0_dec_uops_2_op1_sel : _GEN_5414; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_op2_sel = _T ? io_enq_0_dec_uops_2_op2_sel : _GEN_5406; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_split_num = _T ? io_enq_0_dec_uops_2_split_num : _GEN_5398; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_self_index = _T ? io_enq_0_dec_uops_2_self_index : _GEN_5390; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_rob_inst_idx = _T ? io_enq_0_dec_uops_2_rob_inst_idx : _GEN_5382; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_address_num = _T ? io_enq_0_dec_uops_2_address_num : _GEN_5374; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_uopc = _T ? io_enq_0_dec_uops_2_uopc : _GEN_5366; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_inst = _T ? io_enq_0_dec_uops_2_inst : _GEN_5358; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_debug_inst = _T ? io_enq_0_dec_uops_2_debug_inst : _GEN_5350; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_is_rvc = _T ? io_enq_0_dec_uops_2_is_rvc : _GEN_5342; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_debug_pc = _T ? io_enq_0_dec_uops_2_debug_pc : _GEN_5334; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_iq_type = _T ? io_enq_0_dec_uops_2_iq_type : _GEN_5326; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_fu_code = _T ? io_enq_0_dec_uops_2_fu_code : _GEN_5318; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_ctrl_br_type = _T ? io_enq_0_dec_uops_2_ctrl_br_type : _GEN_5310; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_ctrl_op1_sel = _T ? io_enq_0_dec_uops_2_ctrl_op1_sel : _GEN_5302; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_ctrl_op2_sel = _T ? io_enq_0_dec_uops_2_ctrl_op2_sel : _GEN_5294; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_ctrl_imm_sel = _T ? io_enq_0_dec_uops_2_ctrl_imm_sel : _GEN_5286; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_ctrl_op_fcn = _T ? io_enq_0_dec_uops_2_ctrl_op_fcn : _GEN_5278; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_ctrl_fcn_dw = _T ? io_enq_0_dec_uops_2_ctrl_fcn_dw : _GEN_5270; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_ctrl_csr_cmd = _T ? io_enq_0_dec_uops_2_ctrl_csr_cmd : _GEN_5262; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_ctrl_is_load = _T ? io_enq_0_dec_uops_2_ctrl_is_load : _GEN_5254; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_ctrl_is_sta = _T ? io_enq_0_dec_uops_2_ctrl_is_sta : _GEN_5246; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_ctrl_is_std = _T ? io_enq_0_dec_uops_2_ctrl_is_std : _GEN_5238; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_ctrl_op3_sel = _T ? io_enq_0_dec_uops_2_ctrl_op3_sel : _GEN_5230; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_iw_state = _T ? io_enq_0_dec_uops_2_iw_state : _GEN_5222; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_iw_p1_poisoned = _T ? io_enq_0_dec_uops_2_iw_p1_poisoned : _GEN_5214; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_iw_p2_poisoned = _T ? io_enq_0_dec_uops_2_iw_p2_poisoned : _GEN_5206; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_is_br = _T ? io_enq_0_dec_uops_2_is_br : _GEN_5198; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_is_jalr = _T ? io_enq_0_dec_uops_2_is_jalr : _GEN_5190; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_is_jal = _T ? io_enq_0_dec_uops_2_is_jal : _GEN_5182; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_is_sfb = _T ? io_enq_0_dec_uops_2_is_sfb : _GEN_5174; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_br_mask = _T ? io_enq_0_dec_uops_2_br_mask : _GEN_5166; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_br_tag = _T ? io_enq_0_dec_uops_2_br_tag : _GEN_5158; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_ftq_idx = _T ? io_enq_0_dec_uops_2_ftq_idx : _GEN_5150; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_edge_inst = _T ? io_enq_0_dec_uops_2_edge_inst : _GEN_5142; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_pc_lob = _T ? io_enq_0_dec_uops_2_pc_lob : _GEN_5134; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_taken = _T ? io_enq_0_dec_uops_2_taken : _GEN_5126; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_imm_packed = _T ? io_enq_0_dec_uops_2_imm_packed : _GEN_5118; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_csr_addr = _T ? io_enq_0_dec_uops_2_csr_addr : _GEN_5110; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_rob_idx = _T ? io_enq_0_dec_uops_2_rob_idx : _GEN_5102; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_ldq_idx = _T ? io_enq_0_dec_uops_2_ldq_idx : _GEN_5094; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_stq_idx = _T ? io_enq_0_dec_uops_2_stq_idx : _GEN_5086; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_rxq_idx = _T ? io_enq_0_dec_uops_2_rxq_idx : _GEN_5078; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_pdst = _T ? io_enq_0_dec_uops_2_pdst : _GEN_5070; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_prs1 = _T ? io_enq_0_dec_uops_2_prs1 : _GEN_5062; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_prs2 = _T ? io_enq_0_dec_uops_2_prs2 : _GEN_5054; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_prs3 = _T ? io_enq_0_dec_uops_2_prs3 : _GEN_5046; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_ppred = _T ? io_enq_0_dec_uops_2_ppred : _GEN_5038; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_prs1_busy = _T ? io_enq_0_dec_uops_2_prs1_busy : _GEN_5030; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_prs2_busy = _T ? io_enq_0_dec_uops_2_prs2_busy : _GEN_5022; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_prs3_busy = _T ? io_enq_0_dec_uops_2_prs3_busy : _GEN_5014; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_ppred_busy = _T ? io_enq_0_dec_uops_2_ppred_busy : _GEN_5006; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_stale_pdst = _T ? io_enq_0_dec_uops_2_stale_pdst : _GEN_4998; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_exception = _T ? io_enq_0_dec_uops_2_exception : _GEN_4990; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_exc_cause = _T ? io_enq_0_dec_uops_2_exc_cause : _GEN_4982; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_bypassable = _T ? io_enq_0_dec_uops_2_bypassable : _GEN_4974; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_mem_cmd = _T ? io_enq_0_dec_uops_2_mem_cmd : _GEN_4966; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_mem_size = _T ? io_enq_0_dec_uops_2_mem_size : _GEN_4958; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_mem_signed = _T ? io_enq_0_dec_uops_2_mem_signed : _GEN_4950; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_is_fence = _T ? io_enq_0_dec_uops_2_is_fence : _GEN_4942; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_is_fencei = _T ? io_enq_0_dec_uops_2_is_fencei : _GEN_4934; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_is_amo = _T ? io_enq_0_dec_uops_2_is_amo : _GEN_4926; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_uses_ldq = _T ? io_enq_0_dec_uops_2_uses_ldq : _GEN_4918; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_uses_stq = _T ? io_enq_0_dec_uops_2_uses_stq : _GEN_4910; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_is_sys_pc2epc = _T ? io_enq_0_dec_uops_2_is_sys_pc2epc : _GEN_4902; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_is_unique = _T ? io_enq_0_dec_uops_2_is_unique : _GEN_4894; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_flush_on_commit = _T ? io_enq_0_dec_uops_2_flush_on_commit : _GEN_4886; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_ldst_is_rs1 = _T ? io_enq_0_dec_uops_2_ldst_is_rs1 : _GEN_4878; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_ldst = _T ? io_enq_0_dec_uops_2_ldst : _GEN_4870; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_lrs1 = _T ? io_enq_0_dec_uops_2_lrs1 : _GEN_4862; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_lrs2 = _T ? io_enq_0_dec_uops_2_lrs2 : _GEN_4854; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_lrs3 = _T ? io_enq_0_dec_uops_2_lrs3 : _GEN_4846; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_ldst_val = _T ? io_enq_0_dec_uops_2_ldst_val : _GEN_4838; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_dst_rtype = _T ? io_enq_0_dec_uops_2_dst_rtype : _GEN_4830; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_lrs1_rtype = _T ? io_enq_0_dec_uops_2_lrs1_rtype : _GEN_4822; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_lrs2_rtype = _T ? io_enq_0_dec_uops_2_lrs2_rtype : _GEN_4814; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_frs3_en = _T ? io_enq_0_dec_uops_2_frs3_en : _GEN_4806; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_fp_val = _T ? io_enq_0_dec_uops_2_fp_val : _GEN_4798; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_fp_single = _T ? io_enq_0_dec_uops_2_fp_single : _GEN_4790; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_xcpt_pf_if = _T ? io_enq_0_dec_uops_2_xcpt_pf_if : _GEN_4782; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_xcpt_ae_if = _T ? io_enq_0_dec_uops_2_xcpt_ae_if : _GEN_4774; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_xcpt_ma_if = _T ? io_enq_0_dec_uops_2_xcpt_ma_if : _GEN_4766; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_bp_debug_if = _T ? io_enq_0_dec_uops_2_bp_debug_if : _GEN_4758; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_bp_xcpt_if = _T ? io_enq_0_dec_uops_2_bp_xcpt_if : _GEN_4750; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_debug_fsrc = _T ? io_enq_0_dec_uops_2_debug_fsrc : _GEN_4742; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_2_debug_tsrc = _T ? io_enq_0_dec_uops_2_debug_tsrc : _GEN_4734; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_switch = _T ? io_enq_0_dec_uops_3_switch : _GEN_6278; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_switch_off = _T ? io_enq_0_dec_uops_3_switch_off : _GEN_6270; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_is_unicore = _T ? io_enq_0_dec_uops_3_is_unicore : _GEN_6262; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_shift = _T ? io_enq_0_dec_uops_3_shift : _GEN_6254; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_lrs3_rtype = _T ? io_enq_0_dec_uops_3_lrs3_rtype : _GEN_6246; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_rflag = _T ? io_enq_0_dec_uops_3_rflag : _GEN_6238; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_wflag = _T ? io_enq_0_dec_uops_3_wflag : _GEN_6230; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_prflag = _T ? io_enq_0_dec_uops_3_prflag : _GEN_6222; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_pwflag = _T ? io_enq_0_dec_uops_3_pwflag : _GEN_6214; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_pflag_busy = _T ? io_enq_0_dec_uops_3_pflag_busy : _GEN_6206; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_stale_pflag = _T ? io_enq_0_dec_uops_3_stale_pflag : _GEN_6198; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_op1_sel = _T ? io_enq_0_dec_uops_3_op1_sel : _GEN_6190; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_op2_sel = _T ? io_enq_0_dec_uops_3_op2_sel : _GEN_6182; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_split_num = _T ? io_enq_0_dec_uops_3_split_num : _GEN_6174; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_self_index = _T ? io_enq_0_dec_uops_3_self_index : _GEN_6166; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_rob_inst_idx = _T ? io_enq_0_dec_uops_3_rob_inst_idx : _GEN_6158; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_address_num = _T ? io_enq_0_dec_uops_3_address_num : _GEN_6150; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_uopc = _T ? io_enq_0_dec_uops_3_uopc : _GEN_6142; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_inst = _T ? io_enq_0_dec_uops_3_inst : _GEN_6134; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_debug_inst = _T ? io_enq_0_dec_uops_3_debug_inst : _GEN_6126; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_is_rvc = _T ? io_enq_0_dec_uops_3_is_rvc : _GEN_6118; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_debug_pc = _T ? io_enq_0_dec_uops_3_debug_pc : _GEN_6110; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_iq_type = _T ? io_enq_0_dec_uops_3_iq_type : _GEN_6102; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_fu_code = _T ? io_enq_0_dec_uops_3_fu_code : _GEN_6094; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_ctrl_br_type = _T ? io_enq_0_dec_uops_3_ctrl_br_type : _GEN_6086; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_ctrl_op1_sel = _T ? io_enq_0_dec_uops_3_ctrl_op1_sel : _GEN_6078; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_ctrl_op2_sel = _T ? io_enq_0_dec_uops_3_ctrl_op2_sel : _GEN_6070; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_ctrl_imm_sel = _T ? io_enq_0_dec_uops_3_ctrl_imm_sel : _GEN_6062; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_ctrl_op_fcn = _T ? io_enq_0_dec_uops_3_ctrl_op_fcn : _GEN_6054; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_ctrl_fcn_dw = _T ? io_enq_0_dec_uops_3_ctrl_fcn_dw : _GEN_6046; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_ctrl_csr_cmd = _T ? io_enq_0_dec_uops_3_ctrl_csr_cmd : _GEN_6038; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_ctrl_is_load = _T ? io_enq_0_dec_uops_3_ctrl_is_load : _GEN_6030; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_ctrl_is_sta = _T ? io_enq_0_dec_uops_3_ctrl_is_sta : _GEN_6022; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_ctrl_is_std = _T ? io_enq_0_dec_uops_3_ctrl_is_std : _GEN_6014; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_ctrl_op3_sel = _T ? io_enq_0_dec_uops_3_ctrl_op3_sel : _GEN_6006; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_iw_state = _T ? io_enq_0_dec_uops_3_iw_state : _GEN_5998; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_iw_p1_poisoned = _T ? io_enq_0_dec_uops_3_iw_p1_poisoned : _GEN_5990; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_iw_p2_poisoned = _T ? io_enq_0_dec_uops_3_iw_p2_poisoned : _GEN_5982; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_is_br = _T ? io_enq_0_dec_uops_3_is_br : _GEN_5974; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_is_jalr = _T ? io_enq_0_dec_uops_3_is_jalr : _GEN_5966; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_is_jal = _T ? io_enq_0_dec_uops_3_is_jal : _GEN_5958; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_is_sfb = _T ? io_enq_0_dec_uops_3_is_sfb : _GEN_5950; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_br_mask = _T ? io_enq_0_dec_uops_3_br_mask : _GEN_5942; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_br_tag = _T ? io_enq_0_dec_uops_3_br_tag : _GEN_5934; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_ftq_idx = _T ? io_enq_0_dec_uops_3_ftq_idx : _GEN_5926; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_edge_inst = _T ? io_enq_0_dec_uops_3_edge_inst : _GEN_5918; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_pc_lob = _T ? io_enq_0_dec_uops_3_pc_lob : _GEN_5910; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_taken = _T ? io_enq_0_dec_uops_3_taken : _GEN_5902; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_imm_packed = _T ? io_enq_0_dec_uops_3_imm_packed : _GEN_5894; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_csr_addr = _T ? io_enq_0_dec_uops_3_csr_addr : _GEN_5886; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_rob_idx = _T ? io_enq_0_dec_uops_3_rob_idx : _GEN_5878; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_ldq_idx = _T ? io_enq_0_dec_uops_3_ldq_idx : _GEN_5870; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_stq_idx = _T ? io_enq_0_dec_uops_3_stq_idx : _GEN_5862; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_rxq_idx = _T ? io_enq_0_dec_uops_3_rxq_idx : _GEN_5854; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_pdst = _T ? io_enq_0_dec_uops_3_pdst : _GEN_5846; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_prs1 = _T ? io_enq_0_dec_uops_3_prs1 : _GEN_5838; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_prs2 = _T ? io_enq_0_dec_uops_3_prs2 : _GEN_5830; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_prs3 = _T ? io_enq_0_dec_uops_3_prs3 : _GEN_5822; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_ppred = _T ? io_enq_0_dec_uops_3_ppred : _GEN_5814; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_prs1_busy = _T ? io_enq_0_dec_uops_3_prs1_busy : _GEN_5806; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_prs2_busy = _T ? io_enq_0_dec_uops_3_prs2_busy : _GEN_5798; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_prs3_busy = _T ? io_enq_0_dec_uops_3_prs3_busy : _GEN_5790; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_ppred_busy = _T ? io_enq_0_dec_uops_3_ppred_busy : _GEN_5782; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_stale_pdst = _T ? io_enq_0_dec_uops_3_stale_pdst : _GEN_5774; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_exception = _T ? io_enq_0_dec_uops_3_exception : _GEN_5766; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_exc_cause = _T ? io_enq_0_dec_uops_3_exc_cause : _GEN_5758; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_bypassable = _T ? io_enq_0_dec_uops_3_bypassable : _GEN_5750; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_mem_cmd = _T ? io_enq_0_dec_uops_3_mem_cmd : _GEN_5742; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_mem_size = _T ? io_enq_0_dec_uops_3_mem_size : _GEN_5734; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_mem_signed = _T ? io_enq_0_dec_uops_3_mem_signed : _GEN_5726; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_is_fence = _T ? io_enq_0_dec_uops_3_is_fence : _GEN_5718; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_is_fencei = _T ? io_enq_0_dec_uops_3_is_fencei : _GEN_5710; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_is_amo = _T ? io_enq_0_dec_uops_3_is_amo : _GEN_5702; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_uses_ldq = _T ? io_enq_0_dec_uops_3_uses_ldq : _GEN_5694; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_uses_stq = _T ? io_enq_0_dec_uops_3_uses_stq : _GEN_5686; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_is_sys_pc2epc = _T ? io_enq_0_dec_uops_3_is_sys_pc2epc : _GEN_5678; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_is_unique = _T ? io_enq_0_dec_uops_3_is_unique : _GEN_5670; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_flush_on_commit = _T ? io_enq_0_dec_uops_3_flush_on_commit : _GEN_5662; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_ldst_is_rs1 = _T ? io_enq_0_dec_uops_3_ldst_is_rs1 : _GEN_5654; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_ldst = _T ? io_enq_0_dec_uops_3_ldst : _GEN_5646; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_lrs1 = _T ? io_enq_0_dec_uops_3_lrs1 : _GEN_5638; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_lrs2 = _T ? io_enq_0_dec_uops_3_lrs2 : _GEN_5630; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_lrs3 = _T ? io_enq_0_dec_uops_3_lrs3 : _GEN_5622; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_ldst_val = _T ? io_enq_0_dec_uops_3_ldst_val : _GEN_5614; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_dst_rtype = _T ? io_enq_0_dec_uops_3_dst_rtype : _GEN_5606; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_lrs1_rtype = _T ? io_enq_0_dec_uops_3_lrs1_rtype : _GEN_5598; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_lrs2_rtype = _T ? io_enq_0_dec_uops_3_lrs2_rtype : _GEN_5590; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_frs3_en = _T ? io_enq_0_dec_uops_3_frs3_en : _GEN_5582; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_fp_val = _T ? io_enq_0_dec_uops_3_fp_val : _GEN_5574; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_fp_single = _T ? io_enq_0_dec_uops_3_fp_single : _GEN_5566; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_xcpt_pf_if = _T ? io_enq_0_dec_uops_3_xcpt_pf_if : _GEN_5558; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_xcpt_ae_if = _T ? io_enq_0_dec_uops_3_xcpt_ae_if : _GEN_5550; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_xcpt_ma_if = _T ? io_enq_0_dec_uops_3_xcpt_ma_if : _GEN_5542; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_bp_debug_if = _T ? io_enq_0_dec_uops_3_bp_debug_if : _GEN_5534; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_bp_xcpt_if = _T ? io_enq_0_dec_uops_3_bp_xcpt_if : _GEN_5526; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_debug_fsrc = _T ? io_enq_0_dec_uops_3_debug_fsrc : _GEN_5518; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_dec_uops_3_debug_tsrc = _T ? io_enq_0_dec_uops_3_debug_tsrc : _GEN_5510; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_val_mask_0 = _T ? io_enq_0_val_mask_0 : _GEN_3150; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_val_mask_1 = _T ? io_enq_0_val_mask_1 : _GEN_3158; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_val_mask_2 = _T ? io_enq_0_val_mask_2 : _GEN_3166; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_enq_bits_val_mask_3 = _T ? io_enq_0_val_mask_3 : _GEN_3174; // @[enq_transBuff.scala 125:26 enq_transBuff.scala 126:34 enq_transBuff.scala 130:34]
  assign trans_buffer_io_deq_ready = io_deq_ready; // @[enq_transBuff.scala 42:31]
  assign trans_buffer_io_clear = io_clear; // @[enq_transBuff.scala 40:27]
  assign trans_buffer_io_isUnicoreMode = io_isUnicoreMode; // @[enq_transBuff.scala 41:35]
  always @(posedge clock) begin
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_switch <= io_enq_0_dec_uops_0_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_switch_off <= io_enq_0_dec_uops_0_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_is_unicore <= io_enq_0_dec_uops_0_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_shift <= io_enq_0_dec_uops_0_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_lrs3_rtype <= io_enq_0_dec_uops_0_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_rflag <= io_enq_0_dec_uops_0_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_wflag <= io_enq_0_dec_uops_0_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_prflag <= io_enq_0_dec_uops_0_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_pwflag <= io_enq_0_dec_uops_0_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_pflag_busy <= io_enq_0_dec_uops_0_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_stale_pflag <= io_enq_0_dec_uops_0_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_op1_sel <= io_enq_0_dec_uops_0_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_op2_sel <= io_enq_0_dec_uops_0_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_split_num <= io_enq_0_dec_uops_0_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_self_index <= io_enq_0_dec_uops_0_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_rob_inst_idx <= io_enq_0_dec_uops_0_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_address_num <= io_enq_0_dec_uops_0_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_uopc <= io_enq_0_dec_uops_0_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_inst <= io_enq_0_dec_uops_0_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_debug_inst <= io_enq_0_dec_uops_0_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_is_rvc <= io_enq_0_dec_uops_0_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_debug_pc <= io_enq_0_dec_uops_0_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_iq_type <= io_enq_0_dec_uops_0_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_fu_code <= io_enq_0_dec_uops_0_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_ctrl_br_type <= io_enq_0_dec_uops_0_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_ctrl_op1_sel <= io_enq_0_dec_uops_0_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_ctrl_op2_sel <= io_enq_0_dec_uops_0_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_ctrl_imm_sel <= io_enq_0_dec_uops_0_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_ctrl_op_fcn <= io_enq_0_dec_uops_0_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_ctrl_fcn_dw <= io_enq_0_dec_uops_0_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_ctrl_csr_cmd <= io_enq_0_dec_uops_0_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_ctrl_is_load <= io_enq_0_dec_uops_0_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_ctrl_is_sta <= io_enq_0_dec_uops_0_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_ctrl_is_std <= io_enq_0_dec_uops_0_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_ctrl_op3_sel <= io_enq_0_dec_uops_0_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_iw_state <= io_enq_0_dec_uops_0_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_iw_p1_poisoned <= io_enq_0_dec_uops_0_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_iw_p2_poisoned <= io_enq_0_dec_uops_0_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_is_br <= io_enq_0_dec_uops_0_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_is_jalr <= io_enq_0_dec_uops_0_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_is_jal <= io_enq_0_dec_uops_0_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_is_sfb <= io_enq_0_dec_uops_0_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_br_mask <= io_enq_0_dec_uops_0_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_br_tag <= io_enq_0_dec_uops_0_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_ftq_idx <= io_enq_0_dec_uops_0_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_edge_inst <= io_enq_0_dec_uops_0_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_pc_lob <= io_enq_0_dec_uops_0_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_taken <= io_enq_0_dec_uops_0_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_imm_packed <= io_enq_0_dec_uops_0_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_csr_addr <= io_enq_0_dec_uops_0_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_rob_idx <= io_enq_0_dec_uops_0_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_ldq_idx <= io_enq_0_dec_uops_0_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_stq_idx <= io_enq_0_dec_uops_0_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_rxq_idx <= io_enq_0_dec_uops_0_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_pdst <= io_enq_0_dec_uops_0_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_prs1 <= io_enq_0_dec_uops_0_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_prs2 <= io_enq_0_dec_uops_0_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_prs3 <= io_enq_0_dec_uops_0_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_ppred <= io_enq_0_dec_uops_0_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_prs1_busy <= io_enq_0_dec_uops_0_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_prs2_busy <= io_enq_0_dec_uops_0_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_prs3_busy <= io_enq_0_dec_uops_0_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_ppred_busy <= io_enq_0_dec_uops_0_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_stale_pdst <= io_enq_0_dec_uops_0_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_exception <= io_enq_0_dec_uops_0_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_exc_cause <= io_enq_0_dec_uops_0_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_bypassable <= io_enq_0_dec_uops_0_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_mem_cmd <= io_enq_0_dec_uops_0_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_mem_size <= io_enq_0_dec_uops_0_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_mem_signed <= io_enq_0_dec_uops_0_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_is_fence <= io_enq_0_dec_uops_0_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_is_fencei <= io_enq_0_dec_uops_0_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_is_amo <= io_enq_0_dec_uops_0_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_uses_ldq <= io_enq_0_dec_uops_0_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_uses_stq <= io_enq_0_dec_uops_0_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_is_sys_pc2epc <= io_enq_0_dec_uops_0_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_is_unique <= io_enq_0_dec_uops_0_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_flush_on_commit <= io_enq_0_dec_uops_0_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_ldst_is_rs1 <= io_enq_0_dec_uops_0_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_ldst <= io_enq_0_dec_uops_0_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_lrs1 <= io_enq_0_dec_uops_0_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_lrs2 <= io_enq_0_dec_uops_0_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_lrs3 <= io_enq_0_dec_uops_0_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_ldst_val <= io_enq_0_dec_uops_0_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_dst_rtype <= io_enq_0_dec_uops_0_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_lrs1_rtype <= io_enq_0_dec_uops_0_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_lrs2_rtype <= io_enq_0_dec_uops_0_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_frs3_en <= io_enq_0_dec_uops_0_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_fp_val <= io_enq_0_dec_uops_0_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_fp_single <= io_enq_0_dec_uops_0_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_xcpt_pf_if <= io_enq_0_dec_uops_0_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_xcpt_ae_if <= io_enq_0_dec_uops_0_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_xcpt_ma_if <= io_enq_0_dec_uops_0_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_bp_debug_if <= io_enq_0_dec_uops_0_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_bp_xcpt_if <= io_enq_0_dec_uops_0_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_debug_fsrc <= io_enq_0_dec_uops_0_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_0_debug_tsrc <= io_enq_0_dec_uops_0_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_switch <= io_enq_0_dec_uops_1_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_switch_off <= io_enq_0_dec_uops_1_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_is_unicore <= io_enq_0_dec_uops_1_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_shift <= io_enq_0_dec_uops_1_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_lrs3_rtype <= io_enq_0_dec_uops_1_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_rflag <= io_enq_0_dec_uops_1_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_wflag <= io_enq_0_dec_uops_1_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_prflag <= io_enq_0_dec_uops_1_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_pwflag <= io_enq_0_dec_uops_1_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_pflag_busy <= io_enq_0_dec_uops_1_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_stale_pflag <= io_enq_0_dec_uops_1_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_op1_sel <= io_enq_0_dec_uops_1_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_op2_sel <= io_enq_0_dec_uops_1_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_split_num <= io_enq_0_dec_uops_1_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_self_index <= io_enq_0_dec_uops_1_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_rob_inst_idx <= io_enq_0_dec_uops_1_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_address_num <= io_enq_0_dec_uops_1_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_uopc <= io_enq_0_dec_uops_1_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_inst <= io_enq_0_dec_uops_1_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_debug_inst <= io_enq_0_dec_uops_1_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_is_rvc <= io_enq_0_dec_uops_1_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_debug_pc <= io_enq_0_dec_uops_1_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_iq_type <= io_enq_0_dec_uops_1_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_fu_code <= io_enq_0_dec_uops_1_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_ctrl_br_type <= io_enq_0_dec_uops_1_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_ctrl_op1_sel <= io_enq_0_dec_uops_1_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_ctrl_op2_sel <= io_enq_0_dec_uops_1_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_ctrl_imm_sel <= io_enq_0_dec_uops_1_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_ctrl_op_fcn <= io_enq_0_dec_uops_1_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_ctrl_fcn_dw <= io_enq_0_dec_uops_1_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_ctrl_csr_cmd <= io_enq_0_dec_uops_1_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_ctrl_is_load <= io_enq_0_dec_uops_1_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_ctrl_is_sta <= io_enq_0_dec_uops_1_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_ctrl_is_std <= io_enq_0_dec_uops_1_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_ctrl_op3_sel <= io_enq_0_dec_uops_1_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_iw_state <= io_enq_0_dec_uops_1_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_iw_p1_poisoned <= io_enq_0_dec_uops_1_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_iw_p2_poisoned <= io_enq_0_dec_uops_1_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_is_br <= io_enq_0_dec_uops_1_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_is_jalr <= io_enq_0_dec_uops_1_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_is_jal <= io_enq_0_dec_uops_1_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_is_sfb <= io_enq_0_dec_uops_1_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_br_mask <= io_enq_0_dec_uops_1_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_br_tag <= io_enq_0_dec_uops_1_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_ftq_idx <= io_enq_0_dec_uops_1_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_edge_inst <= io_enq_0_dec_uops_1_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_pc_lob <= io_enq_0_dec_uops_1_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_taken <= io_enq_0_dec_uops_1_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_imm_packed <= io_enq_0_dec_uops_1_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_csr_addr <= io_enq_0_dec_uops_1_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_rob_idx <= io_enq_0_dec_uops_1_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_ldq_idx <= io_enq_0_dec_uops_1_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_stq_idx <= io_enq_0_dec_uops_1_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_rxq_idx <= io_enq_0_dec_uops_1_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_pdst <= io_enq_0_dec_uops_1_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_prs1 <= io_enq_0_dec_uops_1_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_prs2 <= io_enq_0_dec_uops_1_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_prs3 <= io_enq_0_dec_uops_1_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_ppred <= io_enq_0_dec_uops_1_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_prs1_busy <= io_enq_0_dec_uops_1_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_prs2_busy <= io_enq_0_dec_uops_1_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_prs3_busy <= io_enq_0_dec_uops_1_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_ppred_busy <= io_enq_0_dec_uops_1_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_stale_pdst <= io_enq_0_dec_uops_1_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_exception <= io_enq_0_dec_uops_1_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_exc_cause <= io_enq_0_dec_uops_1_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_bypassable <= io_enq_0_dec_uops_1_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_mem_cmd <= io_enq_0_dec_uops_1_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_mem_size <= io_enq_0_dec_uops_1_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_mem_signed <= io_enq_0_dec_uops_1_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_is_fence <= io_enq_0_dec_uops_1_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_is_fencei <= io_enq_0_dec_uops_1_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_is_amo <= io_enq_0_dec_uops_1_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_uses_ldq <= io_enq_0_dec_uops_1_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_uses_stq <= io_enq_0_dec_uops_1_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_is_sys_pc2epc <= io_enq_0_dec_uops_1_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_is_unique <= io_enq_0_dec_uops_1_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_flush_on_commit <= io_enq_0_dec_uops_1_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_ldst_is_rs1 <= io_enq_0_dec_uops_1_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_ldst <= io_enq_0_dec_uops_1_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_lrs1 <= io_enq_0_dec_uops_1_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_lrs2 <= io_enq_0_dec_uops_1_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_lrs3 <= io_enq_0_dec_uops_1_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_ldst_val <= io_enq_0_dec_uops_1_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_dst_rtype <= io_enq_0_dec_uops_1_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_lrs1_rtype <= io_enq_0_dec_uops_1_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_lrs2_rtype <= io_enq_0_dec_uops_1_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_frs3_en <= io_enq_0_dec_uops_1_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_fp_val <= io_enq_0_dec_uops_1_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_fp_single <= io_enq_0_dec_uops_1_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_xcpt_pf_if <= io_enq_0_dec_uops_1_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_xcpt_ae_if <= io_enq_0_dec_uops_1_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_xcpt_ma_if <= io_enq_0_dec_uops_1_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_bp_debug_if <= io_enq_0_dec_uops_1_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_bp_xcpt_if <= io_enq_0_dec_uops_1_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_debug_fsrc <= io_enq_0_dec_uops_1_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_1_debug_tsrc <= io_enq_0_dec_uops_1_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_switch <= io_enq_0_dec_uops_2_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_switch_off <= io_enq_0_dec_uops_2_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_is_unicore <= io_enq_0_dec_uops_2_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_shift <= io_enq_0_dec_uops_2_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_lrs3_rtype <= io_enq_0_dec_uops_2_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_rflag <= io_enq_0_dec_uops_2_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_wflag <= io_enq_0_dec_uops_2_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_prflag <= io_enq_0_dec_uops_2_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_pwflag <= io_enq_0_dec_uops_2_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_pflag_busy <= io_enq_0_dec_uops_2_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_stale_pflag <= io_enq_0_dec_uops_2_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_op1_sel <= io_enq_0_dec_uops_2_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_op2_sel <= io_enq_0_dec_uops_2_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_split_num <= io_enq_0_dec_uops_2_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_self_index <= io_enq_0_dec_uops_2_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_rob_inst_idx <= io_enq_0_dec_uops_2_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_address_num <= io_enq_0_dec_uops_2_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_uopc <= io_enq_0_dec_uops_2_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_inst <= io_enq_0_dec_uops_2_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_debug_inst <= io_enq_0_dec_uops_2_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_is_rvc <= io_enq_0_dec_uops_2_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_debug_pc <= io_enq_0_dec_uops_2_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_iq_type <= io_enq_0_dec_uops_2_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_fu_code <= io_enq_0_dec_uops_2_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_ctrl_br_type <= io_enq_0_dec_uops_2_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_ctrl_op1_sel <= io_enq_0_dec_uops_2_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_ctrl_op2_sel <= io_enq_0_dec_uops_2_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_ctrl_imm_sel <= io_enq_0_dec_uops_2_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_ctrl_op_fcn <= io_enq_0_dec_uops_2_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_ctrl_fcn_dw <= io_enq_0_dec_uops_2_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_ctrl_csr_cmd <= io_enq_0_dec_uops_2_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_ctrl_is_load <= io_enq_0_dec_uops_2_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_ctrl_is_sta <= io_enq_0_dec_uops_2_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_ctrl_is_std <= io_enq_0_dec_uops_2_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_ctrl_op3_sel <= io_enq_0_dec_uops_2_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_iw_state <= io_enq_0_dec_uops_2_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_iw_p1_poisoned <= io_enq_0_dec_uops_2_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_iw_p2_poisoned <= io_enq_0_dec_uops_2_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_is_br <= io_enq_0_dec_uops_2_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_is_jalr <= io_enq_0_dec_uops_2_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_is_jal <= io_enq_0_dec_uops_2_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_is_sfb <= io_enq_0_dec_uops_2_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_br_mask <= io_enq_0_dec_uops_2_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_br_tag <= io_enq_0_dec_uops_2_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_ftq_idx <= io_enq_0_dec_uops_2_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_edge_inst <= io_enq_0_dec_uops_2_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_pc_lob <= io_enq_0_dec_uops_2_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_taken <= io_enq_0_dec_uops_2_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_imm_packed <= io_enq_0_dec_uops_2_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_csr_addr <= io_enq_0_dec_uops_2_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_rob_idx <= io_enq_0_dec_uops_2_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_ldq_idx <= io_enq_0_dec_uops_2_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_stq_idx <= io_enq_0_dec_uops_2_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_rxq_idx <= io_enq_0_dec_uops_2_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_pdst <= io_enq_0_dec_uops_2_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_prs1 <= io_enq_0_dec_uops_2_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_prs2 <= io_enq_0_dec_uops_2_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_prs3 <= io_enq_0_dec_uops_2_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_ppred <= io_enq_0_dec_uops_2_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_prs1_busy <= io_enq_0_dec_uops_2_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_prs2_busy <= io_enq_0_dec_uops_2_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_prs3_busy <= io_enq_0_dec_uops_2_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_ppred_busy <= io_enq_0_dec_uops_2_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_stale_pdst <= io_enq_0_dec_uops_2_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_exception <= io_enq_0_dec_uops_2_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_exc_cause <= io_enq_0_dec_uops_2_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_bypassable <= io_enq_0_dec_uops_2_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_mem_cmd <= io_enq_0_dec_uops_2_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_mem_size <= io_enq_0_dec_uops_2_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_mem_signed <= io_enq_0_dec_uops_2_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_is_fence <= io_enq_0_dec_uops_2_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_is_fencei <= io_enq_0_dec_uops_2_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_is_amo <= io_enq_0_dec_uops_2_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_uses_ldq <= io_enq_0_dec_uops_2_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_uses_stq <= io_enq_0_dec_uops_2_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_is_sys_pc2epc <= io_enq_0_dec_uops_2_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_is_unique <= io_enq_0_dec_uops_2_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_flush_on_commit <= io_enq_0_dec_uops_2_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_ldst_is_rs1 <= io_enq_0_dec_uops_2_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_ldst <= io_enq_0_dec_uops_2_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_lrs1 <= io_enq_0_dec_uops_2_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_lrs2 <= io_enq_0_dec_uops_2_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_lrs3 <= io_enq_0_dec_uops_2_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_ldst_val <= io_enq_0_dec_uops_2_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_dst_rtype <= io_enq_0_dec_uops_2_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_lrs1_rtype <= io_enq_0_dec_uops_2_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_lrs2_rtype <= io_enq_0_dec_uops_2_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_frs3_en <= io_enq_0_dec_uops_2_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_fp_val <= io_enq_0_dec_uops_2_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_fp_single <= io_enq_0_dec_uops_2_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_xcpt_pf_if <= io_enq_0_dec_uops_2_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_xcpt_ae_if <= io_enq_0_dec_uops_2_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_xcpt_ma_if <= io_enq_0_dec_uops_2_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_bp_debug_if <= io_enq_0_dec_uops_2_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_bp_xcpt_if <= io_enq_0_dec_uops_2_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_debug_fsrc <= io_enq_0_dec_uops_2_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_2_debug_tsrc <= io_enq_0_dec_uops_2_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_switch <= io_enq_0_dec_uops_3_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_switch_off <= io_enq_0_dec_uops_3_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_is_unicore <= io_enq_0_dec_uops_3_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_shift <= io_enq_0_dec_uops_3_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_lrs3_rtype <= io_enq_0_dec_uops_3_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_rflag <= io_enq_0_dec_uops_3_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_wflag <= io_enq_0_dec_uops_3_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_prflag <= io_enq_0_dec_uops_3_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_pwflag <= io_enq_0_dec_uops_3_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_pflag_busy <= io_enq_0_dec_uops_3_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_stale_pflag <= io_enq_0_dec_uops_3_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_op1_sel <= io_enq_0_dec_uops_3_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_op2_sel <= io_enq_0_dec_uops_3_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_split_num <= io_enq_0_dec_uops_3_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_self_index <= io_enq_0_dec_uops_3_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_rob_inst_idx <= io_enq_0_dec_uops_3_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_address_num <= io_enq_0_dec_uops_3_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_uopc <= io_enq_0_dec_uops_3_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_inst <= io_enq_0_dec_uops_3_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_debug_inst <= io_enq_0_dec_uops_3_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_is_rvc <= io_enq_0_dec_uops_3_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_debug_pc <= io_enq_0_dec_uops_3_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_iq_type <= io_enq_0_dec_uops_3_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_fu_code <= io_enq_0_dec_uops_3_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_ctrl_br_type <= io_enq_0_dec_uops_3_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_ctrl_op1_sel <= io_enq_0_dec_uops_3_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_ctrl_op2_sel <= io_enq_0_dec_uops_3_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_ctrl_imm_sel <= io_enq_0_dec_uops_3_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_ctrl_op_fcn <= io_enq_0_dec_uops_3_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_ctrl_fcn_dw <= io_enq_0_dec_uops_3_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_ctrl_csr_cmd <= io_enq_0_dec_uops_3_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_ctrl_is_load <= io_enq_0_dec_uops_3_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_ctrl_is_sta <= io_enq_0_dec_uops_3_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_ctrl_is_std <= io_enq_0_dec_uops_3_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_ctrl_op3_sel <= io_enq_0_dec_uops_3_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_iw_state <= io_enq_0_dec_uops_3_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_iw_p1_poisoned <= io_enq_0_dec_uops_3_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_iw_p2_poisoned <= io_enq_0_dec_uops_3_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_is_br <= io_enq_0_dec_uops_3_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_is_jalr <= io_enq_0_dec_uops_3_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_is_jal <= io_enq_0_dec_uops_3_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_is_sfb <= io_enq_0_dec_uops_3_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_br_mask <= io_enq_0_dec_uops_3_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_br_tag <= io_enq_0_dec_uops_3_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_ftq_idx <= io_enq_0_dec_uops_3_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_edge_inst <= io_enq_0_dec_uops_3_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_pc_lob <= io_enq_0_dec_uops_3_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_taken <= io_enq_0_dec_uops_3_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_imm_packed <= io_enq_0_dec_uops_3_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_csr_addr <= io_enq_0_dec_uops_3_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_rob_idx <= io_enq_0_dec_uops_3_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_ldq_idx <= io_enq_0_dec_uops_3_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_stq_idx <= io_enq_0_dec_uops_3_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_rxq_idx <= io_enq_0_dec_uops_3_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_pdst <= io_enq_0_dec_uops_3_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_prs1 <= io_enq_0_dec_uops_3_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_prs2 <= io_enq_0_dec_uops_3_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_prs3 <= io_enq_0_dec_uops_3_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_ppred <= io_enq_0_dec_uops_3_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_prs1_busy <= io_enq_0_dec_uops_3_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_prs2_busy <= io_enq_0_dec_uops_3_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_prs3_busy <= io_enq_0_dec_uops_3_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_ppred_busy <= io_enq_0_dec_uops_3_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_stale_pdst <= io_enq_0_dec_uops_3_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_exception <= io_enq_0_dec_uops_3_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_exc_cause <= io_enq_0_dec_uops_3_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_bypassable <= io_enq_0_dec_uops_3_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_mem_cmd <= io_enq_0_dec_uops_3_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_mem_size <= io_enq_0_dec_uops_3_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_mem_signed <= io_enq_0_dec_uops_3_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_is_fence <= io_enq_0_dec_uops_3_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_is_fencei <= io_enq_0_dec_uops_3_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_is_amo <= io_enq_0_dec_uops_3_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_uses_ldq <= io_enq_0_dec_uops_3_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_uses_stq <= io_enq_0_dec_uops_3_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_is_sys_pc2epc <= io_enq_0_dec_uops_3_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_is_unique <= io_enq_0_dec_uops_3_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_flush_on_commit <= io_enq_0_dec_uops_3_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_ldst_is_rs1 <= io_enq_0_dec_uops_3_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_ldst <= io_enq_0_dec_uops_3_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_lrs1 <= io_enq_0_dec_uops_3_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_lrs2 <= io_enq_0_dec_uops_3_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_lrs3 <= io_enq_0_dec_uops_3_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_ldst_val <= io_enq_0_dec_uops_3_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_dst_rtype <= io_enq_0_dec_uops_3_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_lrs1_rtype <= io_enq_0_dec_uops_3_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_lrs2_rtype <= io_enq_0_dec_uops_3_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_frs3_en <= io_enq_0_dec_uops_3_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_fp_val <= io_enq_0_dec_uops_3_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_fp_single <= io_enq_0_dec_uops_3_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_xcpt_pf_if <= io_enq_0_dec_uops_3_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_xcpt_ae_if <= io_enq_0_dec_uops_3_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_xcpt_ma_if <= io_enq_0_dec_uops_3_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_bp_debug_if <= io_enq_0_dec_uops_3_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_bp_xcpt_if <= io_enq_0_dec_uops_3_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_debug_fsrc <= io_enq_0_dec_uops_3_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_dec_uops_3_debug_tsrc <= io_enq_0_dec_uops_3_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_0_val_mask_0 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_val_mask_0 <= io_enq_0_val_mask_0; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_0_val_mask_1 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_val_mask_1 <= io_enq_0_val_mask_1; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_0_val_mask_2 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_val_mask_2 <= io_enq_0_val_mask_2; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_0_val_mask_3 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_0_val_mask_3 <= io_enq_0_val_mask_3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_switch <= io_enq_1_dec_uops_0_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_switch_off <= io_enq_1_dec_uops_0_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_is_unicore <= io_enq_1_dec_uops_0_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_shift <= io_enq_1_dec_uops_0_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_lrs3_rtype <= io_enq_1_dec_uops_0_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_rflag <= io_enq_1_dec_uops_0_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_wflag <= io_enq_1_dec_uops_0_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_prflag <= io_enq_1_dec_uops_0_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_pwflag <= io_enq_1_dec_uops_0_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_pflag_busy <= io_enq_1_dec_uops_0_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_stale_pflag <= io_enq_1_dec_uops_0_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_op1_sel <= io_enq_1_dec_uops_0_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_op2_sel <= io_enq_1_dec_uops_0_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_split_num <= io_enq_1_dec_uops_0_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_self_index <= io_enq_1_dec_uops_0_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_rob_inst_idx <= io_enq_1_dec_uops_0_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_address_num <= io_enq_1_dec_uops_0_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_uopc <= io_enq_1_dec_uops_0_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_inst <= io_enq_1_dec_uops_0_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_debug_inst <= io_enq_1_dec_uops_0_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_is_rvc <= io_enq_1_dec_uops_0_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_debug_pc <= io_enq_1_dec_uops_0_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_iq_type <= io_enq_1_dec_uops_0_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_fu_code <= io_enq_1_dec_uops_0_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_ctrl_br_type <= io_enq_1_dec_uops_0_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_ctrl_op1_sel <= io_enq_1_dec_uops_0_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_ctrl_op2_sel <= io_enq_1_dec_uops_0_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_ctrl_imm_sel <= io_enq_1_dec_uops_0_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_ctrl_op_fcn <= io_enq_1_dec_uops_0_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_ctrl_fcn_dw <= io_enq_1_dec_uops_0_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_ctrl_csr_cmd <= io_enq_1_dec_uops_0_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_ctrl_is_load <= io_enq_1_dec_uops_0_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_ctrl_is_sta <= io_enq_1_dec_uops_0_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_ctrl_is_std <= io_enq_1_dec_uops_0_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_ctrl_op3_sel <= io_enq_1_dec_uops_0_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_iw_state <= io_enq_1_dec_uops_0_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_iw_p1_poisoned <= io_enq_1_dec_uops_0_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_iw_p2_poisoned <= io_enq_1_dec_uops_0_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_is_br <= io_enq_1_dec_uops_0_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_is_jalr <= io_enq_1_dec_uops_0_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_is_jal <= io_enq_1_dec_uops_0_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_is_sfb <= io_enq_1_dec_uops_0_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_br_mask <= io_enq_1_dec_uops_0_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_br_tag <= io_enq_1_dec_uops_0_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_ftq_idx <= io_enq_1_dec_uops_0_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_edge_inst <= io_enq_1_dec_uops_0_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_pc_lob <= io_enq_1_dec_uops_0_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_taken <= io_enq_1_dec_uops_0_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_imm_packed <= io_enq_1_dec_uops_0_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_csr_addr <= io_enq_1_dec_uops_0_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_rob_idx <= io_enq_1_dec_uops_0_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_ldq_idx <= io_enq_1_dec_uops_0_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_stq_idx <= io_enq_1_dec_uops_0_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_rxq_idx <= io_enq_1_dec_uops_0_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_pdst <= io_enq_1_dec_uops_0_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_prs1 <= io_enq_1_dec_uops_0_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_prs2 <= io_enq_1_dec_uops_0_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_prs3 <= io_enq_1_dec_uops_0_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_ppred <= io_enq_1_dec_uops_0_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_prs1_busy <= io_enq_1_dec_uops_0_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_prs2_busy <= io_enq_1_dec_uops_0_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_prs3_busy <= io_enq_1_dec_uops_0_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_ppred_busy <= io_enq_1_dec_uops_0_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_stale_pdst <= io_enq_1_dec_uops_0_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_exception <= io_enq_1_dec_uops_0_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_exc_cause <= io_enq_1_dec_uops_0_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_bypassable <= io_enq_1_dec_uops_0_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_mem_cmd <= io_enq_1_dec_uops_0_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_mem_size <= io_enq_1_dec_uops_0_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_mem_signed <= io_enq_1_dec_uops_0_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_is_fence <= io_enq_1_dec_uops_0_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_is_fencei <= io_enq_1_dec_uops_0_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_is_amo <= io_enq_1_dec_uops_0_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_uses_ldq <= io_enq_1_dec_uops_0_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_uses_stq <= io_enq_1_dec_uops_0_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_is_sys_pc2epc <= io_enq_1_dec_uops_0_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_is_unique <= io_enq_1_dec_uops_0_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_flush_on_commit <= io_enq_1_dec_uops_0_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_ldst_is_rs1 <= io_enq_1_dec_uops_0_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_ldst <= io_enq_1_dec_uops_0_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_lrs1 <= io_enq_1_dec_uops_0_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_lrs2 <= io_enq_1_dec_uops_0_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_lrs3 <= io_enq_1_dec_uops_0_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_ldst_val <= io_enq_1_dec_uops_0_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_dst_rtype <= io_enq_1_dec_uops_0_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_lrs1_rtype <= io_enq_1_dec_uops_0_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_lrs2_rtype <= io_enq_1_dec_uops_0_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_frs3_en <= io_enq_1_dec_uops_0_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_fp_val <= io_enq_1_dec_uops_0_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_fp_single <= io_enq_1_dec_uops_0_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_xcpt_pf_if <= io_enq_1_dec_uops_0_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_xcpt_ae_if <= io_enq_1_dec_uops_0_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_xcpt_ma_if <= io_enq_1_dec_uops_0_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_bp_debug_if <= io_enq_1_dec_uops_0_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_bp_xcpt_if <= io_enq_1_dec_uops_0_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_debug_fsrc <= io_enq_1_dec_uops_0_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_0_debug_tsrc <= io_enq_1_dec_uops_0_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_switch <= io_enq_1_dec_uops_1_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_switch_off <= io_enq_1_dec_uops_1_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_is_unicore <= io_enq_1_dec_uops_1_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_shift <= io_enq_1_dec_uops_1_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_lrs3_rtype <= io_enq_1_dec_uops_1_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_rflag <= io_enq_1_dec_uops_1_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_wflag <= io_enq_1_dec_uops_1_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_prflag <= io_enq_1_dec_uops_1_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_pwflag <= io_enq_1_dec_uops_1_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_pflag_busy <= io_enq_1_dec_uops_1_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_stale_pflag <= io_enq_1_dec_uops_1_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_op1_sel <= io_enq_1_dec_uops_1_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_op2_sel <= io_enq_1_dec_uops_1_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_split_num <= io_enq_1_dec_uops_1_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_self_index <= io_enq_1_dec_uops_1_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_rob_inst_idx <= io_enq_1_dec_uops_1_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_address_num <= io_enq_1_dec_uops_1_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_uopc <= io_enq_1_dec_uops_1_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_inst <= io_enq_1_dec_uops_1_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_debug_inst <= io_enq_1_dec_uops_1_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_is_rvc <= io_enq_1_dec_uops_1_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_debug_pc <= io_enq_1_dec_uops_1_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_iq_type <= io_enq_1_dec_uops_1_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_fu_code <= io_enq_1_dec_uops_1_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_ctrl_br_type <= io_enq_1_dec_uops_1_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_ctrl_op1_sel <= io_enq_1_dec_uops_1_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_ctrl_op2_sel <= io_enq_1_dec_uops_1_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_ctrl_imm_sel <= io_enq_1_dec_uops_1_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_ctrl_op_fcn <= io_enq_1_dec_uops_1_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_ctrl_fcn_dw <= io_enq_1_dec_uops_1_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_ctrl_csr_cmd <= io_enq_1_dec_uops_1_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_ctrl_is_load <= io_enq_1_dec_uops_1_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_ctrl_is_sta <= io_enq_1_dec_uops_1_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_ctrl_is_std <= io_enq_1_dec_uops_1_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_ctrl_op3_sel <= io_enq_1_dec_uops_1_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_iw_state <= io_enq_1_dec_uops_1_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_iw_p1_poisoned <= io_enq_1_dec_uops_1_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_iw_p2_poisoned <= io_enq_1_dec_uops_1_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_is_br <= io_enq_1_dec_uops_1_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_is_jalr <= io_enq_1_dec_uops_1_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_is_jal <= io_enq_1_dec_uops_1_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_is_sfb <= io_enq_1_dec_uops_1_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_br_mask <= io_enq_1_dec_uops_1_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_br_tag <= io_enq_1_dec_uops_1_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_ftq_idx <= io_enq_1_dec_uops_1_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_edge_inst <= io_enq_1_dec_uops_1_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_pc_lob <= io_enq_1_dec_uops_1_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_taken <= io_enq_1_dec_uops_1_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_imm_packed <= io_enq_1_dec_uops_1_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_csr_addr <= io_enq_1_dec_uops_1_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_rob_idx <= io_enq_1_dec_uops_1_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_ldq_idx <= io_enq_1_dec_uops_1_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_stq_idx <= io_enq_1_dec_uops_1_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_rxq_idx <= io_enq_1_dec_uops_1_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_pdst <= io_enq_1_dec_uops_1_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_prs1 <= io_enq_1_dec_uops_1_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_prs2 <= io_enq_1_dec_uops_1_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_prs3 <= io_enq_1_dec_uops_1_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_ppred <= io_enq_1_dec_uops_1_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_prs1_busy <= io_enq_1_dec_uops_1_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_prs2_busy <= io_enq_1_dec_uops_1_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_prs3_busy <= io_enq_1_dec_uops_1_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_ppred_busy <= io_enq_1_dec_uops_1_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_stale_pdst <= io_enq_1_dec_uops_1_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_exception <= io_enq_1_dec_uops_1_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_exc_cause <= io_enq_1_dec_uops_1_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_bypassable <= io_enq_1_dec_uops_1_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_mem_cmd <= io_enq_1_dec_uops_1_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_mem_size <= io_enq_1_dec_uops_1_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_mem_signed <= io_enq_1_dec_uops_1_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_is_fence <= io_enq_1_dec_uops_1_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_is_fencei <= io_enq_1_dec_uops_1_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_is_amo <= io_enq_1_dec_uops_1_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_uses_ldq <= io_enq_1_dec_uops_1_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_uses_stq <= io_enq_1_dec_uops_1_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_is_sys_pc2epc <= io_enq_1_dec_uops_1_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_is_unique <= io_enq_1_dec_uops_1_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_flush_on_commit <= io_enq_1_dec_uops_1_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_ldst_is_rs1 <= io_enq_1_dec_uops_1_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_ldst <= io_enq_1_dec_uops_1_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_lrs1 <= io_enq_1_dec_uops_1_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_lrs2 <= io_enq_1_dec_uops_1_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_lrs3 <= io_enq_1_dec_uops_1_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_ldst_val <= io_enq_1_dec_uops_1_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_dst_rtype <= io_enq_1_dec_uops_1_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_lrs1_rtype <= io_enq_1_dec_uops_1_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_lrs2_rtype <= io_enq_1_dec_uops_1_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_frs3_en <= io_enq_1_dec_uops_1_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_fp_val <= io_enq_1_dec_uops_1_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_fp_single <= io_enq_1_dec_uops_1_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_xcpt_pf_if <= io_enq_1_dec_uops_1_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_xcpt_ae_if <= io_enq_1_dec_uops_1_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_xcpt_ma_if <= io_enq_1_dec_uops_1_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_bp_debug_if <= io_enq_1_dec_uops_1_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_bp_xcpt_if <= io_enq_1_dec_uops_1_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_debug_fsrc <= io_enq_1_dec_uops_1_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_1_debug_tsrc <= io_enq_1_dec_uops_1_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_switch <= io_enq_1_dec_uops_2_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_switch_off <= io_enq_1_dec_uops_2_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_is_unicore <= io_enq_1_dec_uops_2_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_shift <= io_enq_1_dec_uops_2_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_lrs3_rtype <= io_enq_1_dec_uops_2_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_rflag <= io_enq_1_dec_uops_2_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_wflag <= io_enq_1_dec_uops_2_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_prflag <= io_enq_1_dec_uops_2_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_pwflag <= io_enq_1_dec_uops_2_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_pflag_busy <= io_enq_1_dec_uops_2_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_stale_pflag <= io_enq_1_dec_uops_2_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_op1_sel <= io_enq_1_dec_uops_2_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_op2_sel <= io_enq_1_dec_uops_2_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_split_num <= io_enq_1_dec_uops_2_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_self_index <= io_enq_1_dec_uops_2_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_rob_inst_idx <= io_enq_1_dec_uops_2_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_address_num <= io_enq_1_dec_uops_2_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_uopc <= io_enq_1_dec_uops_2_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_inst <= io_enq_1_dec_uops_2_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_debug_inst <= io_enq_1_dec_uops_2_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_is_rvc <= io_enq_1_dec_uops_2_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_debug_pc <= io_enq_1_dec_uops_2_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_iq_type <= io_enq_1_dec_uops_2_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_fu_code <= io_enq_1_dec_uops_2_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_ctrl_br_type <= io_enq_1_dec_uops_2_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_ctrl_op1_sel <= io_enq_1_dec_uops_2_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_ctrl_op2_sel <= io_enq_1_dec_uops_2_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_ctrl_imm_sel <= io_enq_1_dec_uops_2_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_ctrl_op_fcn <= io_enq_1_dec_uops_2_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_ctrl_fcn_dw <= io_enq_1_dec_uops_2_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_ctrl_csr_cmd <= io_enq_1_dec_uops_2_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_ctrl_is_load <= io_enq_1_dec_uops_2_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_ctrl_is_sta <= io_enq_1_dec_uops_2_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_ctrl_is_std <= io_enq_1_dec_uops_2_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_ctrl_op3_sel <= io_enq_1_dec_uops_2_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_iw_state <= io_enq_1_dec_uops_2_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_iw_p1_poisoned <= io_enq_1_dec_uops_2_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_iw_p2_poisoned <= io_enq_1_dec_uops_2_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_is_br <= io_enq_1_dec_uops_2_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_is_jalr <= io_enq_1_dec_uops_2_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_is_jal <= io_enq_1_dec_uops_2_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_is_sfb <= io_enq_1_dec_uops_2_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_br_mask <= io_enq_1_dec_uops_2_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_br_tag <= io_enq_1_dec_uops_2_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_ftq_idx <= io_enq_1_dec_uops_2_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_edge_inst <= io_enq_1_dec_uops_2_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_pc_lob <= io_enq_1_dec_uops_2_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_taken <= io_enq_1_dec_uops_2_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_imm_packed <= io_enq_1_dec_uops_2_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_csr_addr <= io_enq_1_dec_uops_2_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_rob_idx <= io_enq_1_dec_uops_2_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_ldq_idx <= io_enq_1_dec_uops_2_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_stq_idx <= io_enq_1_dec_uops_2_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_rxq_idx <= io_enq_1_dec_uops_2_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_pdst <= io_enq_1_dec_uops_2_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_prs1 <= io_enq_1_dec_uops_2_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_prs2 <= io_enq_1_dec_uops_2_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_prs3 <= io_enq_1_dec_uops_2_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_ppred <= io_enq_1_dec_uops_2_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_prs1_busy <= io_enq_1_dec_uops_2_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_prs2_busy <= io_enq_1_dec_uops_2_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_prs3_busy <= io_enq_1_dec_uops_2_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_ppred_busy <= io_enq_1_dec_uops_2_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_stale_pdst <= io_enq_1_dec_uops_2_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_exception <= io_enq_1_dec_uops_2_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_exc_cause <= io_enq_1_dec_uops_2_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_bypassable <= io_enq_1_dec_uops_2_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_mem_cmd <= io_enq_1_dec_uops_2_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_mem_size <= io_enq_1_dec_uops_2_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_mem_signed <= io_enq_1_dec_uops_2_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_is_fence <= io_enq_1_dec_uops_2_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_is_fencei <= io_enq_1_dec_uops_2_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_is_amo <= io_enq_1_dec_uops_2_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_uses_ldq <= io_enq_1_dec_uops_2_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_uses_stq <= io_enq_1_dec_uops_2_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_is_sys_pc2epc <= io_enq_1_dec_uops_2_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_is_unique <= io_enq_1_dec_uops_2_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_flush_on_commit <= io_enq_1_dec_uops_2_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_ldst_is_rs1 <= io_enq_1_dec_uops_2_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_ldst <= io_enq_1_dec_uops_2_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_lrs1 <= io_enq_1_dec_uops_2_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_lrs2 <= io_enq_1_dec_uops_2_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_lrs3 <= io_enq_1_dec_uops_2_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_ldst_val <= io_enq_1_dec_uops_2_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_dst_rtype <= io_enq_1_dec_uops_2_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_lrs1_rtype <= io_enq_1_dec_uops_2_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_lrs2_rtype <= io_enq_1_dec_uops_2_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_frs3_en <= io_enq_1_dec_uops_2_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_fp_val <= io_enq_1_dec_uops_2_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_fp_single <= io_enq_1_dec_uops_2_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_xcpt_pf_if <= io_enq_1_dec_uops_2_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_xcpt_ae_if <= io_enq_1_dec_uops_2_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_xcpt_ma_if <= io_enq_1_dec_uops_2_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_bp_debug_if <= io_enq_1_dec_uops_2_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_bp_xcpt_if <= io_enq_1_dec_uops_2_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_debug_fsrc <= io_enq_1_dec_uops_2_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_2_debug_tsrc <= io_enq_1_dec_uops_2_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_switch <= io_enq_1_dec_uops_3_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_switch_off <= io_enq_1_dec_uops_3_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_is_unicore <= io_enq_1_dec_uops_3_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_shift <= io_enq_1_dec_uops_3_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_lrs3_rtype <= io_enq_1_dec_uops_3_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_rflag <= io_enq_1_dec_uops_3_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_wflag <= io_enq_1_dec_uops_3_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_prflag <= io_enq_1_dec_uops_3_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_pwflag <= io_enq_1_dec_uops_3_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_pflag_busy <= io_enq_1_dec_uops_3_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_stale_pflag <= io_enq_1_dec_uops_3_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_op1_sel <= io_enq_1_dec_uops_3_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_op2_sel <= io_enq_1_dec_uops_3_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_split_num <= io_enq_1_dec_uops_3_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_self_index <= io_enq_1_dec_uops_3_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_rob_inst_idx <= io_enq_1_dec_uops_3_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_address_num <= io_enq_1_dec_uops_3_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_uopc <= io_enq_1_dec_uops_3_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_inst <= io_enq_1_dec_uops_3_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_debug_inst <= io_enq_1_dec_uops_3_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_is_rvc <= io_enq_1_dec_uops_3_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_debug_pc <= io_enq_1_dec_uops_3_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_iq_type <= io_enq_1_dec_uops_3_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_fu_code <= io_enq_1_dec_uops_3_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_ctrl_br_type <= io_enq_1_dec_uops_3_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_ctrl_op1_sel <= io_enq_1_dec_uops_3_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_ctrl_op2_sel <= io_enq_1_dec_uops_3_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_ctrl_imm_sel <= io_enq_1_dec_uops_3_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_ctrl_op_fcn <= io_enq_1_dec_uops_3_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_ctrl_fcn_dw <= io_enq_1_dec_uops_3_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_ctrl_csr_cmd <= io_enq_1_dec_uops_3_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_ctrl_is_load <= io_enq_1_dec_uops_3_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_ctrl_is_sta <= io_enq_1_dec_uops_3_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_ctrl_is_std <= io_enq_1_dec_uops_3_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_ctrl_op3_sel <= io_enq_1_dec_uops_3_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_iw_state <= io_enq_1_dec_uops_3_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_iw_p1_poisoned <= io_enq_1_dec_uops_3_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_iw_p2_poisoned <= io_enq_1_dec_uops_3_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_is_br <= io_enq_1_dec_uops_3_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_is_jalr <= io_enq_1_dec_uops_3_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_is_jal <= io_enq_1_dec_uops_3_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_is_sfb <= io_enq_1_dec_uops_3_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_br_mask <= io_enq_1_dec_uops_3_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_br_tag <= io_enq_1_dec_uops_3_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_ftq_idx <= io_enq_1_dec_uops_3_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_edge_inst <= io_enq_1_dec_uops_3_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_pc_lob <= io_enq_1_dec_uops_3_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_taken <= io_enq_1_dec_uops_3_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_imm_packed <= io_enq_1_dec_uops_3_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_csr_addr <= io_enq_1_dec_uops_3_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_rob_idx <= io_enq_1_dec_uops_3_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_ldq_idx <= io_enq_1_dec_uops_3_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_stq_idx <= io_enq_1_dec_uops_3_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_rxq_idx <= io_enq_1_dec_uops_3_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_pdst <= io_enq_1_dec_uops_3_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_prs1 <= io_enq_1_dec_uops_3_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_prs2 <= io_enq_1_dec_uops_3_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_prs3 <= io_enq_1_dec_uops_3_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_ppred <= io_enq_1_dec_uops_3_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_prs1_busy <= io_enq_1_dec_uops_3_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_prs2_busy <= io_enq_1_dec_uops_3_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_prs3_busy <= io_enq_1_dec_uops_3_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_ppred_busy <= io_enq_1_dec_uops_3_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_stale_pdst <= io_enq_1_dec_uops_3_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_exception <= io_enq_1_dec_uops_3_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_exc_cause <= io_enq_1_dec_uops_3_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_bypassable <= io_enq_1_dec_uops_3_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_mem_cmd <= io_enq_1_dec_uops_3_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_mem_size <= io_enq_1_dec_uops_3_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_mem_signed <= io_enq_1_dec_uops_3_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_is_fence <= io_enq_1_dec_uops_3_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_is_fencei <= io_enq_1_dec_uops_3_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_is_amo <= io_enq_1_dec_uops_3_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_uses_ldq <= io_enq_1_dec_uops_3_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_uses_stq <= io_enq_1_dec_uops_3_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_is_sys_pc2epc <= io_enq_1_dec_uops_3_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_is_unique <= io_enq_1_dec_uops_3_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_flush_on_commit <= io_enq_1_dec_uops_3_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_ldst_is_rs1 <= io_enq_1_dec_uops_3_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_ldst <= io_enq_1_dec_uops_3_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_lrs1 <= io_enq_1_dec_uops_3_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_lrs2 <= io_enq_1_dec_uops_3_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_lrs3 <= io_enq_1_dec_uops_3_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_ldst_val <= io_enq_1_dec_uops_3_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_dst_rtype <= io_enq_1_dec_uops_3_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_lrs1_rtype <= io_enq_1_dec_uops_3_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_lrs2_rtype <= io_enq_1_dec_uops_3_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_frs3_en <= io_enq_1_dec_uops_3_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_fp_val <= io_enq_1_dec_uops_3_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_fp_single <= io_enq_1_dec_uops_3_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_xcpt_pf_if <= io_enq_1_dec_uops_3_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_xcpt_ae_if <= io_enq_1_dec_uops_3_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_xcpt_ma_if <= io_enq_1_dec_uops_3_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_bp_debug_if <= io_enq_1_dec_uops_3_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_bp_xcpt_if <= io_enq_1_dec_uops_3_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_debug_fsrc <= io_enq_1_dec_uops_3_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_dec_uops_3_debug_tsrc <= io_enq_1_dec_uops_3_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_1_val_mask_0 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_val_mask_0 <= io_enq_1_val_mask_0; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_1_val_mask_1 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_val_mask_1 <= io_enq_1_val_mask_1; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_1_val_mask_2 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_val_mask_2 <= io_enq_1_val_mask_2; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_1_val_mask_3 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_1_val_mask_3 <= io_enq_1_val_mask_3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_switch <= io_enq_2_dec_uops_0_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_switch_off <= io_enq_2_dec_uops_0_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_is_unicore <= io_enq_2_dec_uops_0_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_shift <= io_enq_2_dec_uops_0_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_lrs3_rtype <= io_enq_2_dec_uops_0_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_rflag <= io_enq_2_dec_uops_0_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_wflag <= io_enq_2_dec_uops_0_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_prflag <= io_enq_2_dec_uops_0_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_pwflag <= io_enq_2_dec_uops_0_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_pflag_busy <= io_enq_2_dec_uops_0_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_stale_pflag <= io_enq_2_dec_uops_0_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_op1_sel <= io_enq_2_dec_uops_0_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_op2_sel <= io_enq_2_dec_uops_0_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_split_num <= io_enq_2_dec_uops_0_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_self_index <= io_enq_2_dec_uops_0_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_rob_inst_idx <= io_enq_2_dec_uops_0_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_address_num <= io_enq_2_dec_uops_0_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_uopc <= io_enq_2_dec_uops_0_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_inst <= io_enq_2_dec_uops_0_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_debug_inst <= io_enq_2_dec_uops_0_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_is_rvc <= io_enq_2_dec_uops_0_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_debug_pc <= io_enq_2_dec_uops_0_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_iq_type <= io_enq_2_dec_uops_0_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_fu_code <= io_enq_2_dec_uops_0_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_ctrl_br_type <= io_enq_2_dec_uops_0_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_ctrl_op1_sel <= io_enq_2_dec_uops_0_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_ctrl_op2_sel <= io_enq_2_dec_uops_0_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_ctrl_imm_sel <= io_enq_2_dec_uops_0_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_ctrl_op_fcn <= io_enq_2_dec_uops_0_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_ctrl_fcn_dw <= io_enq_2_dec_uops_0_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_ctrl_csr_cmd <= io_enq_2_dec_uops_0_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_ctrl_is_load <= io_enq_2_dec_uops_0_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_ctrl_is_sta <= io_enq_2_dec_uops_0_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_ctrl_is_std <= io_enq_2_dec_uops_0_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_ctrl_op3_sel <= io_enq_2_dec_uops_0_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_iw_state <= io_enq_2_dec_uops_0_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_iw_p1_poisoned <= io_enq_2_dec_uops_0_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_iw_p2_poisoned <= io_enq_2_dec_uops_0_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_is_br <= io_enq_2_dec_uops_0_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_is_jalr <= io_enq_2_dec_uops_0_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_is_jal <= io_enq_2_dec_uops_0_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_is_sfb <= io_enq_2_dec_uops_0_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_br_mask <= io_enq_2_dec_uops_0_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_br_tag <= io_enq_2_dec_uops_0_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_ftq_idx <= io_enq_2_dec_uops_0_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_edge_inst <= io_enq_2_dec_uops_0_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_pc_lob <= io_enq_2_dec_uops_0_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_taken <= io_enq_2_dec_uops_0_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_imm_packed <= io_enq_2_dec_uops_0_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_csr_addr <= io_enq_2_dec_uops_0_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_rob_idx <= io_enq_2_dec_uops_0_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_ldq_idx <= io_enq_2_dec_uops_0_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_stq_idx <= io_enq_2_dec_uops_0_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_rxq_idx <= io_enq_2_dec_uops_0_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_pdst <= io_enq_2_dec_uops_0_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_prs1 <= io_enq_2_dec_uops_0_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_prs2 <= io_enq_2_dec_uops_0_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_prs3 <= io_enq_2_dec_uops_0_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_ppred <= io_enq_2_dec_uops_0_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_prs1_busy <= io_enq_2_dec_uops_0_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_prs2_busy <= io_enq_2_dec_uops_0_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_prs3_busy <= io_enq_2_dec_uops_0_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_ppred_busy <= io_enq_2_dec_uops_0_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_stale_pdst <= io_enq_2_dec_uops_0_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_exception <= io_enq_2_dec_uops_0_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_exc_cause <= io_enq_2_dec_uops_0_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_bypassable <= io_enq_2_dec_uops_0_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_mem_cmd <= io_enq_2_dec_uops_0_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_mem_size <= io_enq_2_dec_uops_0_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_mem_signed <= io_enq_2_dec_uops_0_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_is_fence <= io_enq_2_dec_uops_0_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_is_fencei <= io_enq_2_dec_uops_0_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_is_amo <= io_enq_2_dec_uops_0_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_uses_ldq <= io_enq_2_dec_uops_0_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_uses_stq <= io_enq_2_dec_uops_0_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_is_sys_pc2epc <= io_enq_2_dec_uops_0_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_is_unique <= io_enq_2_dec_uops_0_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_flush_on_commit <= io_enq_2_dec_uops_0_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_ldst_is_rs1 <= io_enq_2_dec_uops_0_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_ldst <= io_enq_2_dec_uops_0_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_lrs1 <= io_enq_2_dec_uops_0_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_lrs2 <= io_enq_2_dec_uops_0_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_lrs3 <= io_enq_2_dec_uops_0_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_ldst_val <= io_enq_2_dec_uops_0_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_dst_rtype <= io_enq_2_dec_uops_0_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_lrs1_rtype <= io_enq_2_dec_uops_0_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_lrs2_rtype <= io_enq_2_dec_uops_0_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_frs3_en <= io_enq_2_dec_uops_0_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_fp_val <= io_enq_2_dec_uops_0_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_fp_single <= io_enq_2_dec_uops_0_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_xcpt_pf_if <= io_enq_2_dec_uops_0_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_xcpt_ae_if <= io_enq_2_dec_uops_0_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_xcpt_ma_if <= io_enq_2_dec_uops_0_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_bp_debug_if <= io_enq_2_dec_uops_0_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_bp_xcpt_if <= io_enq_2_dec_uops_0_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_debug_fsrc <= io_enq_2_dec_uops_0_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_0_debug_tsrc <= io_enq_2_dec_uops_0_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_switch <= io_enq_2_dec_uops_1_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_switch_off <= io_enq_2_dec_uops_1_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_is_unicore <= io_enq_2_dec_uops_1_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_shift <= io_enq_2_dec_uops_1_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_lrs3_rtype <= io_enq_2_dec_uops_1_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_rflag <= io_enq_2_dec_uops_1_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_wflag <= io_enq_2_dec_uops_1_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_prflag <= io_enq_2_dec_uops_1_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_pwflag <= io_enq_2_dec_uops_1_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_pflag_busy <= io_enq_2_dec_uops_1_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_stale_pflag <= io_enq_2_dec_uops_1_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_op1_sel <= io_enq_2_dec_uops_1_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_op2_sel <= io_enq_2_dec_uops_1_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_split_num <= io_enq_2_dec_uops_1_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_self_index <= io_enq_2_dec_uops_1_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_rob_inst_idx <= io_enq_2_dec_uops_1_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_address_num <= io_enq_2_dec_uops_1_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_uopc <= io_enq_2_dec_uops_1_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_inst <= io_enq_2_dec_uops_1_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_debug_inst <= io_enq_2_dec_uops_1_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_is_rvc <= io_enq_2_dec_uops_1_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_debug_pc <= io_enq_2_dec_uops_1_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_iq_type <= io_enq_2_dec_uops_1_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_fu_code <= io_enq_2_dec_uops_1_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_ctrl_br_type <= io_enq_2_dec_uops_1_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_ctrl_op1_sel <= io_enq_2_dec_uops_1_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_ctrl_op2_sel <= io_enq_2_dec_uops_1_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_ctrl_imm_sel <= io_enq_2_dec_uops_1_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_ctrl_op_fcn <= io_enq_2_dec_uops_1_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_ctrl_fcn_dw <= io_enq_2_dec_uops_1_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_ctrl_csr_cmd <= io_enq_2_dec_uops_1_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_ctrl_is_load <= io_enq_2_dec_uops_1_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_ctrl_is_sta <= io_enq_2_dec_uops_1_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_ctrl_is_std <= io_enq_2_dec_uops_1_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_ctrl_op3_sel <= io_enq_2_dec_uops_1_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_iw_state <= io_enq_2_dec_uops_1_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_iw_p1_poisoned <= io_enq_2_dec_uops_1_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_iw_p2_poisoned <= io_enq_2_dec_uops_1_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_is_br <= io_enq_2_dec_uops_1_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_is_jalr <= io_enq_2_dec_uops_1_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_is_jal <= io_enq_2_dec_uops_1_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_is_sfb <= io_enq_2_dec_uops_1_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_br_mask <= io_enq_2_dec_uops_1_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_br_tag <= io_enq_2_dec_uops_1_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_ftq_idx <= io_enq_2_dec_uops_1_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_edge_inst <= io_enq_2_dec_uops_1_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_pc_lob <= io_enq_2_dec_uops_1_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_taken <= io_enq_2_dec_uops_1_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_imm_packed <= io_enq_2_dec_uops_1_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_csr_addr <= io_enq_2_dec_uops_1_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_rob_idx <= io_enq_2_dec_uops_1_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_ldq_idx <= io_enq_2_dec_uops_1_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_stq_idx <= io_enq_2_dec_uops_1_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_rxq_idx <= io_enq_2_dec_uops_1_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_pdst <= io_enq_2_dec_uops_1_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_prs1 <= io_enq_2_dec_uops_1_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_prs2 <= io_enq_2_dec_uops_1_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_prs3 <= io_enq_2_dec_uops_1_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_ppred <= io_enq_2_dec_uops_1_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_prs1_busy <= io_enq_2_dec_uops_1_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_prs2_busy <= io_enq_2_dec_uops_1_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_prs3_busy <= io_enq_2_dec_uops_1_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_ppred_busy <= io_enq_2_dec_uops_1_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_stale_pdst <= io_enq_2_dec_uops_1_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_exception <= io_enq_2_dec_uops_1_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_exc_cause <= io_enq_2_dec_uops_1_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_bypassable <= io_enq_2_dec_uops_1_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_mem_cmd <= io_enq_2_dec_uops_1_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_mem_size <= io_enq_2_dec_uops_1_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_mem_signed <= io_enq_2_dec_uops_1_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_is_fence <= io_enq_2_dec_uops_1_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_is_fencei <= io_enq_2_dec_uops_1_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_is_amo <= io_enq_2_dec_uops_1_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_uses_ldq <= io_enq_2_dec_uops_1_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_uses_stq <= io_enq_2_dec_uops_1_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_is_sys_pc2epc <= io_enq_2_dec_uops_1_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_is_unique <= io_enq_2_dec_uops_1_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_flush_on_commit <= io_enq_2_dec_uops_1_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_ldst_is_rs1 <= io_enq_2_dec_uops_1_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_ldst <= io_enq_2_dec_uops_1_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_lrs1 <= io_enq_2_dec_uops_1_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_lrs2 <= io_enq_2_dec_uops_1_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_lrs3 <= io_enq_2_dec_uops_1_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_ldst_val <= io_enq_2_dec_uops_1_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_dst_rtype <= io_enq_2_dec_uops_1_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_lrs1_rtype <= io_enq_2_dec_uops_1_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_lrs2_rtype <= io_enq_2_dec_uops_1_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_frs3_en <= io_enq_2_dec_uops_1_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_fp_val <= io_enq_2_dec_uops_1_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_fp_single <= io_enq_2_dec_uops_1_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_xcpt_pf_if <= io_enq_2_dec_uops_1_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_xcpt_ae_if <= io_enq_2_dec_uops_1_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_xcpt_ma_if <= io_enq_2_dec_uops_1_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_bp_debug_if <= io_enq_2_dec_uops_1_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_bp_xcpt_if <= io_enq_2_dec_uops_1_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_debug_fsrc <= io_enq_2_dec_uops_1_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_1_debug_tsrc <= io_enq_2_dec_uops_1_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_switch <= io_enq_2_dec_uops_2_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_switch_off <= io_enq_2_dec_uops_2_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_is_unicore <= io_enq_2_dec_uops_2_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_shift <= io_enq_2_dec_uops_2_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_lrs3_rtype <= io_enq_2_dec_uops_2_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_rflag <= io_enq_2_dec_uops_2_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_wflag <= io_enq_2_dec_uops_2_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_prflag <= io_enq_2_dec_uops_2_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_pwflag <= io_enq_2_dec_uops_2_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_pflag_busy <= io_enq_2_dec_uops_2_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_stale_pflag <= io_enq_2_dec_uops_2_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_op1_sel <= io_enq_2_dec_uops_2_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_op2_sel <= io_enq_2_dec_uops_2_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_split_num <= io_enq_2_dec_uops_2_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_self_index <= io_enq_2_dec_uops_2_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_rob_inst_idx <= io_enq_2_dec_uops_2_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_address_num <= io_enq_2_dec_uops_2_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_uopc <= io_enq_2_dec_uops_2_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_inst <= io_enq_2_dec_uops_2_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_debug_inst <= io_enq_2_dec_uops_2_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_is_rvc <= io_enq_2_dec_uops_2_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_debug_pc <= io_enq_2_dec_uops_2_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_iq_type <= io_enq_2_dec_uops_2_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_fu_code <= io_enq_2_dec_uops_2_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_ctrl_br_type <= io_enq_2_dec_uops_2_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_ctrl_op1_sel <= io_enq_2_dec_uops_2_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_ctrl_op2_sel <= io_enq_2_dec_uops_2_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_ctrl_imm_sel <= io_enq_2_dec_uops_2_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_ctrl_op_fcn <= io_enq_2_dec_uops_2_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_ctrl_fcn_dw <= io_enq_2_dec_uops_2_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_ctrl_csr_cmd <= io_enq_2_dec_uops_2_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_ctrl_is_load <= io_enq_2_dec_uops_2_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_ctrl_is_sta <= io_enq_2_dec_uops_2_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_ctrl_is_std <= io_enq_2_dec_uops_2_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_ctrl_op3_sel <= io_enq_2_dec_uops_2_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_iw_state <= io_enq_2_dec_uops_2_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_iw_p1_poisoned <= io_enq_2_dec_uops_2_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_iw_p2_poisoned <= io_enq_2_dec_uops_2_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_is_br <= io_enq_2_dec_uops_2_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_is_jalr <= io_enq_2_dec_uops_2_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_is_jal <= io_enq_2_dec_uops_2_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_is_sfb <= io_enq_2_dec_uops_2_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_br_mask <= io_enq_2_dec_uops_2_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_br_tag <= io_enq_2_dec_uops_2_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_ftq_idx <= io_enq_2_dec_uops_2_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_edge_inst <= io_enq_2_dec_uops_2_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_pc_lob <= io_enq_2_dec_uops_2_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_taken <= io_enq_2_dec_uops_2_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_imm_packed <= io_enq_2_dec_uops_2_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_csr_addr <= io_enq_2_dec_uops_2_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_rob_idx <= io_enq_2_dec_uops_2_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_ldq_idx <= io_enq_2_dec_uops_2_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_stq_idx <= io_enq_2_dec_uops_2_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_rxq_idx <= io_enq_2_dec_uops_2_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_pdst <= io_enq_2_dec_uops_2_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_prs1 <= io_enq_2_dec_uops_2_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_prs2 <= io_enq_2_dec_uops_2_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_prs3 <= io_enq_2_dec_uops_2_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_ppred <= io_enq_2_dec_uops_2_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_prs1_busy <= io_enq_2_dec_uops_2_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_prs2_busy <= io_enq_2_dec_uops_2_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_prs3_busy <= io_enq_2_dec_uops_2_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_ppred_busy <= io_enq_2_dec_uops_2_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_stale_pdst <= io_enq_2_dec_uops_2_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_exception <= io_enq_2_dec_uops_2_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_exc_cause <= io_enq_2_dec_uops_2_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_bypassable <= io_enq_2_dec_uops_2_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_mem_cmd <= io_enq_2_dec_uops_2_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_mem_size <= io_enq_2_dec_uops_2_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_mem_signed <= io_enq_2_dec_uops_2_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_is_fence <= io_enq_2_dec_uops_2_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_is_fencei <= io_enq_2_dec_uops_2_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_is_amo <= io_enq_2_dec_uops_2_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_uses_ldq <= io_enq_2_dec_uops_2_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_uses_stq <= io_enq_2_dec_uops_2_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_is_sys_pc2epc <= io_enq_2_dec_uops_2_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_is_unique <= io_enq_2_dec_uops_2_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_flush_on_commit <= io_enq_2_dec_uops_2_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_ldst_is_rs1 <= io_enq_2_dec_uops_2_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_ldst <= io_enq_2_dec_uops_2_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_lrs1 <= io_enq_2_dec_uops_2_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_lrs2 <= io_enq_2_dec_uops_2_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_lrs3 <= io_enq_2_dec_uops_2_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_ldst_val <= io_enq_2_dec_uops_2_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_dst_rtype <= io_enq_2_dec_uops_2_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_lrs1_rtype <= io_enq_2_dec_uops_2_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_lrs2_rtype <= io_enq_2_dec_uops_2_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_frs3_en <= io_enq_2_dec_uops_2_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_fp_val <= io_enq_2_dec_uops_2_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_fp_single <= io_enq_2_dec_uops_2_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_xcpt_pf_if <= io_enq_2_dec_uops_2_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_xcpt_ae_if <= io_enq_2_dec_uops_2_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_xcpt_ma_if <= io_enq_2_dec_uops_2_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_bp_debug_if <= io_enq_2_dec_uops_2_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_bp_xcpt_if <= io_enq_2_dec_uops_2_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_debug_fsrc <= io_enq_2_dec_uops_2_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_2_debug_tsrc <= io_enq_2_dec_uops_2_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_switch <= io_enq_2_dec_uops_3_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_switch_off <= io_enq_2_dec_uops_3_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_is_unicore <= io_enq_2_dec_uops_3_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_shift <= io_enq_2_dec_uops_3_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_lrs3_rtype <= io_enq_2_dec_uops_3_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_rflag <= io_enq_2_dec_uops_3_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_wflag <= io_enq_2_dec_uops_3_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_prflag <= io_enq_2_dec_uops_3_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_pwflag <= io_enq_2_dec_uops_3_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_pflag_busy <= io_enq_2_dec_uops_3_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_stale_pflag <= io_enq_2_dec_uops_3_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_op1_sel <= io_enq_2_dec_uops_3_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_op2_sel <= io_enq_2_dec_uops_3_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_split_num <= io_enq_2_dec_uops_3_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_self_index <= io_enq_2_dec_uops_3_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_rob_inst_idx <= io_enq_2_dec_uops_3_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_address_num <= io_enq_2_dec_uops_3_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_uopc <= io_enq_2_dec_uops_3_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_inst <= io_enq_2_dec_uops_3_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_debug_inst <= io_enq_2_dec_uops_3_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_is_rvc <= io_enq_2_dec_uops_3_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_debug_pc <= io_enq_2_dec_uops_3_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_iq_type <= io_enq_2_dec_uops_3_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_fu_code <= io_enq_2_dec_uops_3_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_ctrl_br_type <= io_enq_2_dec_uops_3_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_ctrl_op1_sel <= io_enq_2_dec_uops_3_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_ctrl_op2_sel <= io_enq_2_dec_uops_3_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_ctrl_imm_sel <= io_enq_2_dec_uops_3_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_ctrl_op_fcn <= io_enq_2_dec_uops_3_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_ctrl_fcn_dw <= io_enq_2_dec_uops_3_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_ctrl_csr_cmd <= io_enq_2_dec_uops_3_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_ctrl_is_load <= io_enq_2_dec_uops_3_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_ctrl_is_sta <= io_enq_2_dec_uops_3_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_ctrl_is_std <= io_enq_2_dec_uops_3_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_ctrl_op3_sel <= io_enq_2_dec_uops_3_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_iw_state <= io_enq_2_dec_uops_3_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_iw_p1_poisoned <= io_enq_2_dec_uops_3_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_iw_p2_poisoned <= io_enq_2_dec_uops_3_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_is_br <= io_enq_2_dec_uops_3_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_is_jalr <= io_enq_2_dec_uops_3_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_is_jal <= io_enq_2_dec_uops_3_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_is_sfb <= io_enq_2_dec_uops_3_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_br_mask <= io_enq_2_dec_uops_3_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_br_tag <= io_enq_2_dec_uops_3_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_ftq_idx <= io_enq_2_dec_uops_3_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_edge_inst <= io_enq_2_dec_uops_3_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_pc_lob <= io_enq_2_dec_uops_3_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_taken <= io_enq_2_dec_uops_3_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_imm_packed <= io_enq_2_dec_uops_3_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_csr_addr <= io_enq_2_dec_uops_3_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_rob_idx <= io_enq_2_dec_uops_3_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_ldq_idx <= io_enq_2_dec_uops_3_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_stq_idx <= io_enq_2_dec_uops_3_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_rxq_idx <= io_enq_2_dec_uops_3_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_pdst <= io_enq_2_dec_uops_3_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_prs1 <= io_enq_2_dec_uops_3_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_prs2 <= io_enq_2_dec_uops_3_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_prs3 <= io_enq_2_dec_uops_3_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_ppred <= io_enq_2_dec_uops_3_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_prs1_busy <= io_enq_2_dec_uops_3_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_prs2_busy <= io_enq_2_dec_uops_3_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_prs3_busy <= io_enq_2_dec_uops_3_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_ppred_busy <= io_enq_2_dec_uops_3_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_stale_pdst <= io_enq_2_dec_uops_3_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_exception <= io_enq_2_dec_uops_3_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_exc_cause <= io_enq_2_dec_uops_3_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_bypassable <= io_enq_2_dec_uops_3_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_mem_cmd <= io_enq_2_dec_uops_3_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_mem_size <= io_enq_2_dec_uops_3_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_mem_signed <= io_enq_2_dec_uops_3_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_is_fence <= io_enq_2_dec_uops_3_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_is_fencei <= io_enq_2_dec_uops_3_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_is_amo <= io_enq_2_dec_uops_3_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_uses_ldq <= io_enq_2_dec_uops_3_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_uses_stq <= io_enq_2_dec_uops_3_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_is_sys_pc2epc <= io_enq_2_dec_uops_3_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_is_unique <= io_enq_2_dec_uops_3_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_flush_on_commit <= io_enq_2_dec_uops_3_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_ldst_is_rs1 <= io_enq_2_dec_uops_3_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_ldst <= io_enq_2_dec_uops_3_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_lrs1 <= io_enq_2_dec_uops_3_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_lrs2 <= io_enq_2_dec_uops_3_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_lrs3 <= io_enq_2_dec_uops_3_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_ldst_val <= io_enq_2_dec_uops_3_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_dst_rtype <= io_enq_2_dec_uops_3_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_lrs1_rtype <= io_enq_2_dec_uops_3_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_lrs2_rtype <= io_enq_2_dec_uops_3_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_frs3_en <= io_enq_2_dec_uops_3_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_fp_val <= io_enq_2_dec_uops_3_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_fp_single <= io_enq_2_dec_uops_3_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_xcpt_pf_if <= io_enq_2_dec_uops_3_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_xcpt_ae_if <= io_enq_2_dec_uops_3_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_xcpt_ma_if <= io_enq_2_dec_uops_3_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_bp_debug_if <= io_enq_2_dec_uops_3_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_bp_xcpt_if <= io_enq_2_dec_uops_3_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_debug_fsrc <= io_enq_2_dec_uops_3_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_dec_uops_3_debug_tsrc <= io_enq_2_dec_uops_3_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_2_val_mask_0 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_val_mask_0 <= io_enq_2_val_mask_0; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_2_val_mask_1 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_val_mask_1 <= io_enq_2_val_mask_1; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_2_val_mask_2 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_val_mask_2 <= io_enq_2_val_mask_2; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_2_val_mask_3 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_2_val_mask_3 <= io_enq_2_val_mask_3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_switch <= io_enq_3_dec_uops_0_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_switch_off <= io_enq_3_dec_uops_0_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_is_unicore <= io_enq_3_dec_uops_0_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_shift <= io_enq_3_dec_uops_0_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_lrs3_rtype <= io_enq_3_dec_uops_0_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_rflag <= io_enq_3_dec_uops_0_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_wflag <= io_enq_3_dec_uops_0_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_prflag <= io_enq_3_dec_uops_0_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_pwflag <= io_enq_3_dec_uops_0_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_pflag_busy <= io_enq_3_dec_uops_0_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_stale_pflag <= io_enq_3_dec_uops_0_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_op1_sel <= io_enq_3_dec_uops_0_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_op2_sel <= io_enq_3_dec_uops_0_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_split_num <= io_enq_3_dec_uops_0_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_self_index <= io_enq_3_dec_uops_0_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_rob_inst_idx <= io_enq_3_dec_uops_0_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_address_num <= io_enq_3_dec_uops_0_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_uopc <= io_enq_3_dec_uops_0_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_inst <= io_enq_3_dec_uops_0_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_debug_inst <= io_enq_3_dec_uops_0_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_is_rvc <= io_enq_3_dec_uops_0_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_debug_pc <= io_enq_3_dec_uops_0_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_iq_type <= io_enq_3_dec_uops_0_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_fu_code <= io_enq_3_dec_uops_0_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_ctrl_br_type <= io_enq_3_dec_uops_0_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_ctrl_op1_sel <= io_enq_3_dec_uops_0_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_ctrl_op2_sel <= io_enq_3_dec_uops_0_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_ctrl_imm_sel <= io_enq_3_dec_uops_0_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_ctrl_op_fcn <= io_enq_3_dec_uops_0_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_ctrl_fcn_dw <= io_enq_3_dec_uops_0_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_ctrl_csr_cmd <= io_enq_3_dec_uops_0_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_ctrl_is_load <= io_enq_3_dec_uops_0_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_ctrl_is_sta <= io_enq_3_dec_uops_0_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_ctrl_is_std <= io_enq_3_dec_uops_0_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_ctrl_op3_sel <= io_enq_3_dec_uops_0_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_iw_state <= io_enq_3_dec_uops_0_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_iw_p1_poisoned <= io_enq_3_dec_uops_0_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_iw_p2_poisoned <= io_enq_3_dec_uops_0_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_is_br <= io_enq_3_dec_uops_0_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_is_jalr <= io_enq_3_dec_uops_0_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_is_jal <= io_enq_3_dec_uops_0_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_is_sfb <= io_enq_3_dec_uops_0_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_br_mask <= io_enq_3_dec_uops_0_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_br_tag <= io_enq_3_dec_uops_0_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_ftq_idx <= io_enq_3_dec_uops_0_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_edge_inst <= io_enq_3_dec_uops_0_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_pc_lob <= io_enq_3_dec_uops_0_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_taken <= io_enq_3_dec_uops_0_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_imm_packed <= io_enq_3_dec_uops_0_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_csr_addr <= io_enq_3_dec_uops_0_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_rob_idx <= io_enq_3_dec_uops_0_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_ldq_idx <= io_enq_3_dec_uops_0_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_stq_idx <= io_enq_3_dec_uops_0_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_rxq_idx <= io_enq_3_dec_uops_0_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_pdst <= io_enq_3_dec_uops_0_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_prs1 <= io_enq_3_dec_uops_0_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_prs2 <= io_enq_3_dec_uops_0_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_prs3 <= io_enq_3_dec_uops_0_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_ppred <= io_enq_3_dec_uops_0_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_prs1_busy <= io_enq_3_dec_uops_0_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_prs2_busy <= io_enq_3_dec_uops_0_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_prs3_busy <= io_enq_3_dec_uops_0_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_ppred_busy <= io_enq_3_dec_uops_0_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_stale_pdst <= io_enq_3_dec_uops_0_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_exception <= io_enq_3_dec_uops_0_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_exc_cause <= io_enq_3_dec_uops_0_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_bypassable <= io_enq_3_dec_uops_0_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_mem_cmd <= io_enq_3_dec_uops_0_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_mem_size <= io_enq_3_dec_uops_0_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_mem_signed <= io_enq_3_dec_uops_0_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_is_fence <= io_enq_3_dec_uops_0_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_is_fencei <= io_enq_3_dec_uops_0_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_is_amo <= io_enq_3_dec_uops_0_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_uses_ldq <= io_enq_3_dec_uops_0_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_uses_stq <= io_enq_3_dec_uops_0_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_is_sys_pc2epc <= io_enq_3_dec_uops_0_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_is_unique <= io_enq_3_dec_uops_0_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_flush_on_commit <= io_enq_3_dec_uops_0_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_ldst_is_rs1 <= io_enq_3_dec_uops_0_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_ldst <= io_enq_3_dec_uops_0_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_lrs1 <= io_enq_3_dec_uops_0_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_lrs2 <= io_enq_3_dec_uops_0_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_lrs3 <= io_enq_3_dec_uops_0_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_ldst_val <= io_enq_3_dec_uops_0_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_dst_rtype <= io_enq_3_dec_uops_0_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_lrs1_rtype <= io_enq_3_dec_uops_0_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_lrs2_rtype <= io_enq_3_dec_uops_0_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_frs3_en <= io_enq_3_dec_uops_0_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_fp_val <= io_enq_3_dec_uops_0_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_fp_single <= io_enq_3_dec_uops_0_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_xcpt_pf_if <= io_enq_3_dec_uops_0_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_xcpt_ae_if <= io_enq_3_dec_uops_0_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_xcpt_ma_if <= io_enq_3_dec_uops_0_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_bp_debug_if <= io_enq_3_dec_uops_0_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_bp_xcpt_if <= io_enq_3_dec_uops_0_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_debug_fsrc <= io_enq_3_dec_uops_0_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_0_debug_tsrc <= io_enq_3_dec_uops_0_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_switch <= io_enq_3_dec_uops_1_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_switch_off <= io_enq_3_dec_uops_1_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_is_unicore <= io_enq_3_dec_uops_1_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_shift <= io_enq_3_dec_uops_1_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_lrs3_rtype <= io_enq_3_dec_uops_1_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_rflag <= io_enq_3_dec_uops_1_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_wflag <= io_enq_3_dec_uops_1_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_prflag <= io_enq_3_dec_uops_1_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_pwflag <= io_enq_3_dec_uops_1_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_pflag_busy <= io_enq_3_dec_uops_1_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_stale_pflag <= io_enq_3_dec_uops_1_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_op1_sel <= io_enq_3_dec_uops_1_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_op2_sel <= io_enq_3_dec_uops_1_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_split_num <= io_enq_3_dec_uops_1_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_self_index <= io_enq_3_dec_uops_1_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_rob_inst_idx <= io_enq_3_dec_uops_1_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_address_num <= io_enq_3_dec_uops_1_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_uopc <= io_enq_3_dec_uops_1_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_inst <= io_enq_3_dec_uops_1_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_debug_inst <= io_enq_3_dec_uops_1_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_is_rvc <= io_enq_3_dec_uops_1_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_debug_pc <= io_enq_3_dec_uops_1_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_iq_type <= io_enq_3_dec_uops_1_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_fu_code <= io_enq_3_dec_uops_1_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_ctrl_br_type <= io_enq_3_dec_uops_1_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_ctrl_op1_sel <= io_enq_3_dec_uops_1_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_ctrl_op2_sel <= io_enq_3_dec_uops_1_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_ctrl_imm_sel <= io_enq_3_dec_uops_1_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_ctrl_op_fcn <= io_enq_3_dec_uops_1_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_ctrl_fcn_dw <= io_enq_3_dec_uops_1_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_ctrl_csr_cmd <= io_enq_3_dec_uops_1_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_ctrl_is_load <= io_enq_3_dec_uops_1_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_ctrl_is_sta <= io_enq_3_dec_uops_1_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_ctrl_is_std <= io_enq_3_dec_uops_1_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_ctrl_op3_sel <= io_enq_3_dec_uops_1_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_iw_state <= io_enq_3_dec_uops_1_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_iw_p1_poisoned <= io_enq_3_dec_uops_1_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_iw_p2_poisoned <= io_enq_3_dec_uops_1_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_is_br <= io_enq_3_dec_uops_1_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_is_jalr <= io_enq_3_dec_uops_1_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_is_jal <= io_enq_3_dec_uops_1_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_is_sfb <= io_enq_3_dec_uops_1_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_br_mask <= io_enq_3_dec_uops_1_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_br_tag <= io_enq_3_dec_uops_1_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_ftq_idx <= io_enq_3_dec_uops_1_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_edge_inst <= io_enq_3_dec_uops_1_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_pc_lob <= io_enq_3_dec_uops_1_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_taken <= io_enq_3_dec_uops_1_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_imm_packed <= io_enq_3_dec_uops_1_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_csr_addr <= io_enq_3_dec_uops_1_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_rob_idx <= io_enq_3_dec_uops_1_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_ldq_idx <= io_enq_3_dec_uops_1_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_stq_idx <= io_enq_3_dec_uops_1_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_rxq_idx <= io_enq_3_dec_uops_1_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_pdst <= io_enq_3_dec_uops_1_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_prs1 <= io_enq_3_dec_uops_1_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_prs2 <= io_enq_3_dec_uops_1_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_prs3 <= io_enq_3_dec_uops_1_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_ppred <= io_enq_3_dec_uops_1_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_prs1_busy <= io_enq_3_dec_uops_1_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_prs2_busy <= io_enq_3_dec_uops_1_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_prs3_busy <= io_enq_3_dec_uops_1_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_ppred_busy <= io_enq_3_dec_uops_1_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_stale_pdst <= io_enq_3_dec_uops_1_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_exception <= io_enq_3_dec_uops_1_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_exc_cause <= io_enq_3_dec_uops_1_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_bypassable <= io_enq_3_dec_uops_1_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_mem_cmd <= io_enq_3_dec_uops_1_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_mem_size <= io_enq_3_dec_uops_1_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_mem_signed <= io_enq_3_dec_uops_1_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_is_fence <= io_enq_3_dec_uops_1_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_is_fencei <= io_enq_3_dec_uops_1_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_is_amo <= io_enq_3_dec_uops_1_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_uses_ldq <= io_enq_3_dec_uops_1_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_uses_stq <= io_enq_3_dec_uops_1_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_is_sys_pc2epc <= io_enq_3_dec_uops_1_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_is_unique <= io_enq_3_dec_uops_1_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_flush_on_commit <= io_enq_3_dec_uops_1_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_ldst_is_rs1 <= io_enq_3_dec_uops_1_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_ldst <= io_enq_3_dec_uops_1_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_lrs1 <= io_enq_3_dec_uops_1_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_lrs2 <= io_enq_3_dec_uops_1_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_lrs3 <= io_enq_3_dec_uops_1_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_ldst_val <= io_enq_3_dec_uops_1_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_dst_rtype <= io_enq_3_dec_uops_1_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_lrs1_rtype <= io_enq_3_dec_uops_1_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_lrs2_rtype <= io_enq_3_dec_uops_1_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_frs3_en <= io_enq_3_dec_uops_1_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_fp_val <= io_enq_3_dec_uops_1_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_fp_single <= io_enq_3_dec_uops_1_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_xcpt_pf_if <= io_enq_3_dec_uops_1_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_xcpt_ae_if <= io_enq_3_dec_uops_1_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_xcpt_ma_if <= io_enq_3_dec_uops_1_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_bp_debug_if <= io_enq_3_dec_uops_1_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_bp_xcpt_if <= io_enq_3_dec_uops_1_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_debug_fsrc <= io_enq_3_dec_uops_1_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_1_debug_tsrc <= io_enq_3_dec_uops_1_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_switch <= io_enq_3_dec_uops_2_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_switch_off <= io_enq_3_dec_uops_2_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_is_unicore <= io_enq_3_dec_uops_2_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_shift <= io_enq_3_dec_uops_2_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_lrs3_rtype <= io_enq_3_dec_uops_2_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_rflag <= io_enq_3_dec_uops_2_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_wflag <= io_enq_3_dec_uops_2_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_prflag <= io_enq_3_dec_uops_2_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_pwflag <= io_enq_3_dec_uops_2_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_pflag_busy <= io_enq_3_dec_uops_2_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_stale_pflag <= io_enq_3_dec_uops_2_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_op1_sel <= io_enq_3_dec_uops_2_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_op2_sel <= io_enq_3_dec_uops_2_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_split_num <= io_enq_3_dec_uops_2_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_self_index <= io_enq_3_dec_uops_2_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_rob_inst_idx <= io_enq_3_dec_uops_2_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_address_num <= io_enq_3_dec_uops_2_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_uopc <= io_enq_3_dec_uops_2_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_inst <= io_enq_3_dec_uops_2_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_debug_inst <= io_enq_3_dec_uops_2_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_is_rvc <= io_enq_3_dec_uops_2_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_debug_pc <= io_enq_3_dec_uops_2_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_iq_type <= io_enq_3_dec_uops_2_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_fu_code <= io_enq_3_dec_uops_2_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_ctrl_br_type <= io_enq_3_dec_uops_2_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_ctrl_op1_sel <= io_enq_3_dec_uops_2_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_ctrl_op2_sel <= io_enq_3_dec_uops_2_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_ctrl_imm_sel <= io_enq_3_dec_uops_2_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_ctrl_op_fcn <= io_enq_3_dec_uops_2_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_ctrl_fcn_dw <= io_enq_3_dec_uops_2_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_ctrl_csr_cmd <= io_enq_3_dec_uops_2_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_ctrl_is_load <= io_enq_3_dec_uops_2_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_ctrl_is_sta <= io_enq_3_dec_uops_2_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_ctrl_is_std <= io_enq_3_dec_uops_2_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_ctrl_op3_sel <= io_enq_3_dec_uops_2_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_iw_state <= io_enq_3_dec_uops_2_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_iw_p1_poisoned <= io_enq_3_dec_uops_2_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_iw_p2_poisoned <= io_enq_3_dec_uops_2_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_is_br <= io_enq_3_dec_uops_2_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_is_jalr <= io_enq_3_dec_uops_2_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_is_jal <= io_enq_3_dec_uops_2_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_is_sfb <= io_enq_3_dec_uops_2_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_br_mask <= io_enq_3_dec_uops_2_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_br_tag <= io_enq_3_dec_uops_2_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_ftq_idx <= io_enq_3_dec_uops_2_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_edge_inst <= io_enq_3_dec_uops_2_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_pc_lob <= io_enq_3_dec_uops_2_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_taken <= io_enq_3_dec_uops_2_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_imm_packed <= io_enq_3_dec_uops_2_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_csr_addr <= io_enq_3_dec_uops_2_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_rob_idx <= io_enq_3_dec_uops_2_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_ldq_idx <= io_enq_3_dec_uops_2_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_stq_idx <= io_enq_3_dec_uops_2_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_rxq_idx <= io_enq_3_dec_uops_2_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_pdst <= io_enq_3_dec_uops_2_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_prs1 <= io_enq_3_dec_uops_2_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_prs2 <= io_enq_3_dec_uops_2_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_prs3 <= io_enq_3_dec_uops_2_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_ppred <= io_enq_3_dec_uops_2_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_prs1_busy <= io_enq_3_dec_uops_2_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_prs2_busy <= io_enq_3_dec_uops_2_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_prs3_busy <= io_enq_3_dec_uops_2_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_ppred_busy <= io_enq_3_dec_uops_2_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_stale_pdst <= io_enq_3_dec_uops_2_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_exception <= io_enq_3_dec_uops_2_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_exc_cause <= io_enq_3_dec_uops_2_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_bypassable <= io_enq_3_dec_uops_2_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_mem_cmd <= io_enq_3_dec_uops_2_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_mem_size <= io_enq_3_dec_uops_2_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_mem_signed <= io_enq_3_dec_uops_2_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_is_fence <= io_enq_3_dec_uops_2_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_is_fencei <= io_enq_3_dec_uops_2_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_is_amo <= io_enq_3_dec_uops_2_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_uses_ldq <= io_enq_3_dec_uops_2_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_uses_stq <= io_enq_3_dec_uops_2_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_is_sys_pc2epc <= io_enq_3_dec_uops_2_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_is_unique <= io_enq_3_dec_uops_2_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_flush_on_commit <= io_enq_3_dec_uops_2_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_ldst_is_rs1 <= io_enq_3_dec_uops_2_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_ldst <= io_enq_3_dec_uops_2_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_lrs1 <= io_enq_3_dec_uops_2_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_lrs2 <= io_enq_3_dec_uops_2_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_lrs3 <= io_enq_3_dec_uops_2_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_ldst_val <= io_enq_3_dec_uops_2_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_dst_rtype <= io_enq_3_dec_uops_2_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_lrs1_rtype <= io_enq_3_dec_uops_2_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_lrs2_rtype <= io_enq_3_dec_uops_2_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_frs3_en <= io_enq_3_dec_uops_2_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_fp_val <= io_enq_3_dec_uops_2_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_fp_single <= io_enq_3_dec_uops_2_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_xcpt_pf_if <= io_enq_3_dec_uops_2_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_xcpt_ae_if <= io_enq_3_dec_uops_2_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_xcpt_ma_if <= io_enq_3_dec_uops_2_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_bp_debug_if <= io_enq_3_dec_uops_2_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_bp_xcpt_if <= io_enq_3_dec_uops_2_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_debug_fsrc <= io_enq_3_dec_uops_2_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_2_debug_tsrc <= io_enq_3_dec_uops_2_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_switch <= io_enq_3_dec_uops_3_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_switch_off <= io_enq_3_dec_uops_3_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_is_unicore <= io_enq_3_dec_uops_3_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_shift <= io_enq_3_dec_uops_3_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_lrs3_rtype <= io_enq_3_dec_uops_3_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_rflag <= io_enq_3_dec_uops_3_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_wflag <= io_enq_3_dec_uops_3_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_prflag <= io_enq_3_dec_uops_3_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_pwflag <= io_enq_3_dec_uops_3_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_pflag_busy <= io_enq_3_dec_uops_3_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_stale_pflag <= io_enq_3_dec_uops_3_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_op1_sel <= io_enq_3_dec_uops_3_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_op2_sel <= io_enq_3_dec_uops_3_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_split_num <= io_enq_3_dec_uops_3_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_self_index <= io_enq_3_dec_uops_3_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_rob_inst_idx <= io_enq_3_dec_uops_3_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_address_num <= io_enq_3_dec_uops_3_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_uopc <= io_enq_3_dec_uops_3_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_inst <= io_enq_3_dec_uops_3_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_debug_inst <= io_enq_3_dec_uops_3_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_is_rvc <= io_enq_3_dec_uops_3_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_debug_pc <= io_enq_3_dec_uops_3_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_iq_type <= io_enq_3_dec_uops_3_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_fu_code <= io_enq_3_dec_uops_3_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_ctrl_br_type <= io_enq_3_dec_uops_3_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_ctrl_op1_sel <= io_enq_3_dec_uops_3_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_ctrl_op2_sel <= io_enq_3_dec_uops_3_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_ctrl_imm_sel <= io_enq_3_dec_uops_3_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_ctrl_op_fcn <= io_enq_3_dec_uops_3_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_ctrl_fcn_dw <= io_enq_3_dec_uops_3_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_ctrl_csr_cmd <= io_enq_3_dec_uops_3_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_ctrl_is_load <= io_enq_3_dec_uops_3_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_ctrl_is_sta <= io_enq_3_dec_uops_3_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_ctrl_is_std <= io_enq_3_dec_uops_3_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_ctrl_op3_sel <= io_enq_3_dec_uops_3_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_iw_state <= io_enq_3_dec_uops_3_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_iw_p1_poisoned <= io_enq_3_dec_uops_3_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_iw_p2_poisoned <= io_enq_3_dec_uops_3_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_is_br <= io_enq_3_dec_uops_3_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_is_jalr <= io_enq_3_dec_uops_3_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_is_jal <= io_enq_3_dec_uops_3_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_is_sfb <= io_enq_3_dec_uops_3_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_br_mask <= io_enq_3_dec_uops_3_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_br_tag <= io_enq_3_dec_uops_3_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_ftq_idx <= io_enq_3_dec_uops_3_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_edge_inst <= io_enq_3_dec_uops_3_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_pc_lob <= io_enq_3_dec_uops_3_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_taken <= io_enq_3_dec_uops_3_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_imm_packed <= io_enq_3_dec_uops_3_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_csr_addr <= io_enq_3_dec_uops_3_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_rob_idx <= io_enq_3_dec_uops_3_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_ldq_idx <= io_enq_3_dec_uops_3_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_stq_idx <= io_enq_3_dec_uops_3_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_rxq_idx <= io_enq_3_dec_uops_3_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_pdst <= io_enq_3_dec_uops_3_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_prs1 <= io_enq_3_dec_uops_3_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_prs2 <= io_enq_3_dec_uops_3_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_prs3 <= io_enq_3_dec_uops_3_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_ppred <= io_enq_3_dec_uops_3_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_prs1_busy <= io_enq_3_dec_uops_3_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_prs2_busy <= io_enq_3_dec_uops_3_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_prs3_busy <= io_enq_3_dec_uops_3_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_ppred_busy <= io_enq_3_dec_uops_3_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_stale_pdst <= io_enq_3_dec_uops_3_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_exception <= io_enq_3_dec_uops_3_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_exc_cause <= io_enq_3_dec_uops_3_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_bypassable <= io_enq_3_dec_uops_3_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_mem_cmd <= io_enq_3_dec_uops_3_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_mem_size <= io_enq_3_dec_uops_3_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_mem_signed <= io_enq_3_dec_uops_3_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_is_fence <= io_enq_3_dec_uops_3_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_is_fencei <= io_enq_3_dec_uops_3_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_is_amo <= io_enq_3_dec_uops_3_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_uses_ldq <= io_enq_3_dec_uops_3_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_uses_stq <= io_enq_3_dec_uops_3_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_is_sys_pc2epc <= io_enq_3_dec_uops_3_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_is_unique <= io_enq_3_dec_uops_3_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_flush_on_commit <= io_enq_3_dec_uops_3_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_ldst_is_rs1 <= io_enq_3_dec_uops_3_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_ldst <= io_enq_3_dec_uops_3_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_lrs1 <= io_enq_3_dec_uops_3_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_lrs2 <= io_enq_3_dec_uops_3_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_lrs3 <= io_enq_3_dec_uops_3_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_ldst_val <= io_enq_3_dec_uops_3_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_dst_rtype <= io_enq_3_dec_uops_3_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_lrs1_rtype <= io_enq_3_dec_uops_3_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_lrs2_rtype <= io_enq_3_dec_uops_3_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_frs3_en <= io_enq_3_dec_uops_3_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_fp_val <= io_enq_3_dec_uops_3_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_fp_single <= io_enq_3_dec_uops_3_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_xcpt_pf_if <= io_enq_3_dec_uops_3_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_xcpt_ae_if <= io_enq_3_dec_uops_3_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_xcpt_ma_if <= io_enq_3_dec_uops_3_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_bp_debug_if <= io_enq_3_dec_uops_3_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_bp_xcpt_if <= io_enq_3_dec_uops_3_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_debug_fsrc <= io_enq_3_dec_uops_3_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_dec_uops_3_debug_tsrc <= io_enq_3_dec_uops_3_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_3_val_mask_0 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_val_mask_0 <= io_enq_3_val_mask_0; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_3_val_mask_1 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_val_mask_1 <= io_enq_3_val_mask_1; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_3_val_mask_2 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_val_mask_2 <= io_enq_3_val_mask_2; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_3_val_mask_3 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_3_val_mask_3 <= io_enq_3_val_mask_3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_switch <= io_enq_4_dec_uops_0_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_switch_off <= io_enq_4_dec_uops_0_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_is_unicore <= io_enq_4_dec_uops_0_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_shift <= io_enq_4_dec_uops_0_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_lrs3_rtype <= io_enq_4_dec_uops_0_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_rflag <= io_enq_4_dec_uops_0_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_wflag <= io_enq_4_dec_uops_0_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_prflag <= io_enq_4_dec_uops_0_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_pwflag <= io_enq_4_dec_uops_0_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_pflag_busy <= io_enq_4_dec_uops_0_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_stale_pflag <= io_enq_4_dec_uops_0_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_op1_sel <= io_enq_4_dec_uops_0_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_op2_sel <= io_enq_4_dec_uops_0_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_split_num <= io_enq_4_dec_uops_0_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_self_index <= io_enq_4_dec_uops_0_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_rob_inst_idx <= io_enq_4_dec_uops_0_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_address_num <= io_enq_4_dec_uops_0_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_uopc <= io_enq_4_dec_uops_0_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_inst <= io_enq_4_dec_uops_0_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_debug_inst <= io_enq_4_dec_uops_0_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_is_rvc <= io_enq_4_dec_uops_0_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_debug_pc <= io_enq_4_dec_uops_0_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_iq_type <= io_enq_4_dec_uops_0_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_fu_code <= io_enq_4_dec_uops_0_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_ctrl_br_type <= io_enq_4_dec_uops_0_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_ctrl_op1_sel <= io_enq_4_dec_uops_0_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_ctrl_op2_sel <= io_enq_4_dec_uops_0_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_ctrl_imm_sel <= io_enq_4_dec_uops_0_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_ctrl_op_fcn <= io_enq_4_dec_uops_0_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_ctrl_fcn_dw <= io_enq_4_dec_uops_0_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_ctrl_csr_cmd <= io_enq_4_dec_uops_0_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_ctrl_is_load <= io_enq_4_dec_uops_0_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_ctrl_is_sta <= io_enq_4_dec_uops_0_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_ctrl_is_std <= io_enq_4_dec_uops_0_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_ctrl_op3_sel <= io_enq_4_dec_uops_0_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_iw_state <= io_enq_4_dec_uops_0_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_iw_p1_poisoned <= io_enq_4_dec_uops_0_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_iw_p2_poisoned <= io_enq_4_dec_uops_0_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_is_br <= io_enq_4_dec_uops_0_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_is_jalr <= io_enq_4_dec_uops_0_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_is_jal <= io_enq_4_dec_uops_0_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_is_sfb <= io_enq_4_dec_uops_0_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_br_mask <= io_enq_4_dec_uops_0_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_br_tag <= io_enq_4_dec_uops_0_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_ftq_idx <= io_enq_4_dec_uops_0_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_edge_inst <= io_enq_4_dec_uops_0_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_pc_lob <= io_enq_4_dec_uops_0_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_taken <= io_enq_4_dec_uops_0_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_imm_packed <= io_enq_4_dec_uops_0_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_csr_addr <= io_enq_4_dec_uops_0_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_rob_idx <= io_enq_4_dec_uops_0_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_ldq_idx <= io_enq_4_dec_uops_0_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_stq_idx <= io_enq_4_dec_uops_0_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_rxq_idx <= io_enq_4_dec_uops_0_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_pdst <= io_enq_4_dec_uops_0_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_prs1 <= io_enq_4_dec_uops_0_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_prs2 <= io_enq_4_dec_uops_0_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_prs3 <= io_enq_4_dec_uops_0_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_ppred <= io_enq_4_dec_uops_0_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_prs1_busy <= io_enq_4_dec_uops_0_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_prs2_busy <= io_enq_4_dec_uops_0_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_prs3_busy <= io_enq_4_dec_uops_0_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_ppred_busy <= io_enq_4_dec_uops_0_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_stale_pdst <= io_enq_4_dec_uops_0_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_exception <= io_enq_4_dec_uops_0_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_exc_cause <= io_enq_4_dec_uops_0_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_bypassable <= io_enq_4_dec_uops_0_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_mem_cmd <= io_enq_4_dec_uops_0_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_mem_size <= io_enq_4_dec_uops_0_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_mem_signed <= io_enq_4_dec_uops_0_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_is_fence <= io_enq_4_dec_uops_0_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_is_fencei <= io_enq_4_dec_uops_0_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_is_amo <= io_enq_4_dec_uops_0_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_uses_ldq <= io_enq_4_dec_uops_0_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_uses_stq <= io_enq_4_dec_uops_0_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_is_sys_pc2epc <= io_enq_4_dec_uops_0_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_is_unique <= io_enq_4_dec_uops_0_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_flush_on_commit <= io_enq_4_dec_uops_0_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_ldst_is_rs1 <= io_enq_4_dec_uops_0_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_ldst <= io_enq_4_dec_uops_0_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_lrs1 <= io_enq_4_dec_uops_0_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_lrs2 <= io_enq_4_dec_uops_0_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_lrs3 <= io_enq_4_dec_uops_0_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_ldst_val <= io_enq_4_dec_uops_0_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_dst_rtype <= io_enq_4_dec_uops_0_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_lrs1_rtype <= io_enq_4_dec_uops_0_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_lrs2_rtype <= io_enq_4_dec_uops_0_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_frs3_en <= io_enq_4_dec_uops_0_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_fp_val <= io_enq_4_dec_uops_0_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_fp_single <= io_enq_4_dec_uops_0_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_xcpt_pf_if <= io_enq_4_dec_uops_0_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_xcpt_ae_if <= io_enq_4_dec_uops_0_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_xcpt_ma_if <= io_enq_4_dec_uops_0_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_bp_debug_if <= io_enq_4_dec_uops_0_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_bp_xcpt_if <= io_enq_4_dec_uops_0_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_debug_fsrc <= io_enq_4_dec_uops_0_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_0_debug_tsrc <= io_enq_4_dec_uops_0_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_switch <= io_enq_4_dec_uops_1_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_switch_off <= io_enq_4_dec_uops_1_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_is_unicore <= io_enq_4_dec_uops_1_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_shift <= io_enq_4_dec_uops_1_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_lrs3_rtype <= io_enq_4_dec_uops_1_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_rflag <= io_enq_4_dec_uops_1_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_wflag <= io_enq_4_dec_uops_1_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_prflag <= io_enq_4_dec_uops_1_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_pwflag <= io_enq_4_dec_uops_1_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_pflag_busy <= io_enq_4_dec_uops_1_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_stale_pflag <= io_enq_4_dec_uops_1_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_op1_sel <= io_enq_4_dec_uops_1_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_op2_sel <= io_enq_4_dec_uops_1_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_split_num <= io_enq_4_dec_uops_1_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_self_index <= io_enq_4_dec_uops_1_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_rob_inst_idx <= io_enq_4_dec_uops_1_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_address_num <= io_enq_4_dec_uops_1_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_uopc <= io_enq_4_dec_uops_1_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_inst <= io_enq_4_dec_uops_1_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_debug_inst <= io_enq_4_dec_uops_1_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_is_rvc <= io_enq_4_dec_uops_1_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_debug_pc <= io_enq_4_dec_uops_1_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_iq_type <= io_enq_4_dec_uops_1_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_fu_code <= io_enq_4_dec_uops_1_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_ctrl_br_type <= io_enq_4_dec_uops_1_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_ctrl_op1_sel <= io_enq_4_dec_uops_1_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_ctrl_op2_sel <= io_enq_4_dec_uops_1_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_ctrl_imm_sel <= io_enq_4_dec_uops_1_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_ctrl_op_fcn <= io_enq_4_dec_uops_1_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_ctrl_fcn_dw <= io_enq_4_dec_uops_1_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_ctrl_csr_cmd <= io_enq_4_dec_uops_1_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_ctrl_is_load <= io_enq_4_dec_uops_1_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_ctrl_is_sta <= io_enq_4_dec_uops_1_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_ctrl_is_std <= io_enq_4_dec_uops_1_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_ctrl_op3_sel <= io_enq_4_dec_uops_1_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_iw_state <= io_enq_4_dec_uops_1_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_iw_p1_poisoned <= io_enq_4_dec_uops_1_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_iw_p2_poisoned <= io_enq_4_dec_uops_1_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_is_br <= io_enq_4_dec_uops_1_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_is_jalr <= io_enq_4_dec_uops_1_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_is_jal <= io_enq_4_dec_uops_1_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_is_sfb <= io_enq_4_dec_uops_1_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_br_mask <= io_enq_4_dec_uops_1_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_br_tag <= io_enq_4_dec_uops_1_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_ftq_idx <= io_enq_4_dec_uops_1_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_edge_inst <= io_enq_4_dec_uops_1_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_pc_lob <= io_enq_4_dec_uops_1_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_taken <= io_enq_4_dec_uops_1_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_imm_packed <= io_enq_4_dec_uops_1_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_csr_addr <= io_enq_4_dec_uops_1_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_rob_idx <= io_enq_4_dec_uops_1_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_ldq_idx <= io_enq_4_dec_uops_1_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_stq_idx <= io_enq_4_dec_uops_1_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_rxq_idx <= io_enq_4_dec_uops_1_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_pdst <= io_enq_4_dec_uops_1_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_prs1 <= io_enq_4_dec_uops_1_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_prs2 <= io_enq_4_dec_uops_1_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_prs3 <= io_enq_4_dec_uops_1_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_ppred <= io_enq_4_dec_uops_1_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_prs1_busy <= io_enq_4_dec_uops_1_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_prs2_busy <= io_enq_4_dec_uops_1_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_prs3_busy <= io_enq_4_dec_uops_1_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_ppred_busy <= io_enq_4_dec_uops_1_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_stale_pdst <= io_enq_4_dec_uops_1_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_exception <= io_enq_4_dec_uops_1_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_exc_cause <= io_enq_4_dec_uops_1_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_bypassable <= io_enq_4_dec_uops_1_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_mem_cmd <= io_enq_4_dec_uops_1_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_mem_size <= io_enq_4_dec_uops_1_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_mem_signed <= io_enq_4_dec_uops_1_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_is_fence <= io_enq_4_dec_uops_1_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_is_fencei <= io_enq_4_dec_uops_1_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_is_amo <= io_enq_4_dec_uops_1_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_uses_ldq <= io_enq_4_dec_uops_1_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_uses_stq <= io_enq_4_dec_uops_1_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_is_sys_pc2epc <= io_enq_4_dec_uops_1_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_is_unique <= io_enq_4_dec_uops_1_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_flush_on_commit <= io_enq_4_dec_uops_1_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_ldst_is_rs1 <= io_enq_4_dec_uops_1_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_ldst <= io_enq_4_dec_uops_1_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_lrs1 <= io_enq_4_dec_uops_1_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_lrs2 <= io_enq_4_dec_uops_1_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_lrs3 <= io_enq_4_dec_uops_1_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_ldst_val <= io_enq_4_dec_uops_1_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_dst_rtype <= io_enq_4_dec_uops_1_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_lrs1_rtype <= io_enq_4_dec_uops_1_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_lrs2_rtype <= io_enq_4_dec_uops_1_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_frs3_en <= io_enq_4_dec_uops_1_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_fp_val <= io_enq_4_dec_uops_1_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_fp_single <= io_enq_4_dec_uops_1_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_xcpt_pf_if <= io_enq_4_dec_uops_1_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_xcpt_ae_if <= io_enq_4_dec_uops_1_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_xcpt_ma_if <= io_enq_4_dec_uops_1_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_bp_debug_if <= io_enq_4_dec_uops_1_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_bp_xcpt_if <= io_enq_4_dec_uops_1_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_debug_fsrc <= io_enq_4_dec_uops_1_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_1_debug_tsrc <= io_enq_4_dec_uops_1_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_switch <= io_enq_4_dec_uops_2_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_switch_off <= io_enq_4_dec_uops_2_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_is_unicore <= io_enq_4_dec_uops_2_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_shift <= io_enq_4_dec_uops_2_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_lrs3_rtype <= io_enq_4_dec_uops_2_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_rflag <= io_enq_4_dec_uops_2_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_wflag <= io_enq_4_dec_uops_2_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_prflag <= io_enq_4_dec_uops_2_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_pwflag <= io_enq_4_dec_uops_2_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_pflag_busy <= io_enq_4_dec_uops_2_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_stale_pflag <= io_enq_4_dec_uops_2_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_op1_sel <= io_enq_4_dec_uops_2_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_op2_sel <= io_enq_4_dec_uops_2_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_split_num <= io_enq_4_dec_uops_2_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_self_index <= io_enq_4_dec_uops_2_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_rob_inst_idx <= io_enq_4_dec_uops_2_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_address_num <= io_enq_4_dec_uops_2_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_uopc <= io_enq_4_dec_uops_2_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_inst <= io_enq_4_dec_uops_2_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_debug_inst <= io_enq_4_dec_uops_2_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_is_rvc <= io_enq_4_dec_uops_2_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_debug_pc <= io_enq_4_dec_uops_2_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_iq_type <= io_enq_4_dec_uops_2_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_fu_code <= io_enq_4_dec_uops_2_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_ctrl_br_type <= io_enq_4_dec_uops_2_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_ctrl_op1_sel <= io_enq_4_dec_uops_2_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_ctrl_op2_sel <= io_enq_4_dec_uops_2_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_ctrl_imm_sel <= io_enq_4_dec_uops_2_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_ctrl_op_fcn <= io_enq_4_dec_uops_2_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_ctrl_fcn_dw <= io_enq_4_dec_uops_2_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_ctrl_csr_cmd <= io_enq_4_dec_uops_2_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_ctrl_is_load <= io_enq_4_dec_uops_2_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_ctrl_is_sta <= io_enq_4_dec_uops_2_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_ctrl_is_std <= io_enq_4_dec_uops_2_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_ctrl_op3_sel <= io_enq_4_dec_uops_2_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_iw_state <= io_enq_4_dec_uops_2_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_iw_p1_poisoned <= io_enq_4_dec_uops_2_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_iw_p2_poisoned <= io_enq_4_dec_uops_2_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_is_br <= io_enq_4_dec_uops_2_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_is_jalr <= io_enq_4_dec_uops_2_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_is_jal <= io_enq_4_dec_uops_2_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_is_sfb <= io_enq_4_dec_uops_2_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_br_mask <= io_enq_4_dec_uops_2_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_br_tag <= io_enq_4_dec_uops_2_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_ftq_idx <= io_enq_4_dec_uops_2_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_edge_inst <= io_enq_4_dec_uops_2_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_pc_lob <= io_enq_4_dec_uops_2_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_taken <= io_enq_4_dec_uops_2_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_imm_packed <= io_enq_4_dec_uops_2_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_csr_addr <= io_enq_4_dec_uops_2_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_rob_idx <= io_enq_4_dec_uops_2_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_ldq_idx <= io_enq_4_dec_uops_2_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_stq_idx <= io_enq_4_dec_uops_2_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_rxq_idx <= io_enq_4_dec_uops_2_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_pdst <= io_enq_4_dec_uops_2_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_prs1 <= io_enq_4_dec_uops_2_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_prs2 <= io_enq_4_dec_uops_2_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_prs3 <= io_enq_4_dec_uops_2_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_ppred <= io_enq_4_dec_uops_2_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_prs1_busy <= io_enq_4_dec_uops_2_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_prs2_busy <= io_enq_4_dec_uops_2_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_prs3_busy <= io_enq_4_dec_uops_2_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_ppred_busy <= io_enq_4_dec_uops_2_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_stale_pdst <= io_enq_4_dec_uops_2_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_exception <= io_enq_4_dec_uops_2_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_exc_cause <= io_enq_4_dec_uops_2_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_bypassable <= io_enq_4_dec_uops_2_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_mem_cmd <= io_enq_4_dec_uops_2_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_mem_size <= io_enq_4_dec_uops_2_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_mem_signed <= io_enq_4_dec_uops_2_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_is_fence <= io_enq_4_dec_uops_2_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_is_fencei <= io_enq_4_dec_uops_2_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_is_amo <= io_enq_4_dec_uops_2_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_uses_ldq <= io_enq_4_dec_uops_2_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_uses_stq <= io_enq_4_dec_uops_2_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_is_sys_pc2epc <= io_enq_4_dec_uops_2_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_is_unique <= io_enq_4_dec_uops_2_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_flush_on_commit <= io_enq_4_dec_uops_2_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_ldst_is_rs1 <= io_enq_4_dec_uops_2_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_ldst <= io_enq_4_dec_uops_2_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_lrs1 <= io_enq_4_dec_uops_2_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_lrs2 <= io_enq_4_dec_uops_2_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_lrs3 <= io_enq_4_dec_uops_2_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_ldst_val <= io_enq_4_dec_uops_2_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_dst_rtype <= io_enq_4_dec_uops_2_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_lrs1_rtype <= io_enq_4_dec_uops_2_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_lrs2_rtype <= io_enq_4_dec_uops_2_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_frs3_en <= io_enq_4_dec_uops_2_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_fp_val <= io_enq_4_dec_uops_2_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_fp_single <= io_enq_4_dec_uops_2_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_xcpt_pf_if <= io_enq_4_dec_uops_2_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_xcpt_ae_if <= io_enq_4_dec_uops_2_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_xcpt_ma_if <= io_enq_4_dec_uops_2_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_bp_debug_if <= io_enq_4_dec_uops_2_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_bp_xcpt_if <= io_enq_4_dec_uops_2_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_debug_fsrc <= io_enq_4_dec_uops_2_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_2_debug_tsrc <= io_enq_4_dec_uops_2_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_switch <= io_enq_4_dec_uops_3_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_switch_off <= io_enq_4_dec_uops_3_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_is_unicore <= io_enq_4_dec_uops_3_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_shift <= io_enq_4_dec_uops_3_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_lrs3_rtype <= io_enq_4_dec_uops_3_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_rflag <= io_enq_4_dec_uops_3_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_wflag <= io_enq_4_dec_uops_3_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_prflag <= io_enq_4_dec_uops_3_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_pwflag <= io_enq_4_dec_uops_3_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_pflag_busy <= io_enq_4_dec_uops_3_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_stale_pflag <= io_enq_4_dec_uops_3_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_op1_sel <= io_enq_4_dec_uops_3_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_op2_sel <= io_enq_4_dec_uops_3_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_split_num <= io_enq_4_dec_uops_3_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_self_index <= io_enq_4_dec_uops_3_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_rob_inst_idx <= io_enq_4_dec_uops_3_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_address_num <= io_enq_4_dec_uops_3_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_uopc <= io_enq_4_dec_uops_3_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_inst <= io_enq_4_dec_uops_3_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_debug_inst <= io_enq_4_dec_uops_3_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_is_rvc <= io_enq_4_dec_uops_3_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_debug_pc <= io_enq_4_dec_uops_3_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_iq_type <= io_enq_4_dec_uops_3_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_fu_code <= io_enq_4_dec_uops_3_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_ctrl_br_type <= io_enq_4_dec_uops_3_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_ctrl_op1_sel <= io_enq_4_dec_uops_3_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_ctrl_op2_sel <= io_enq_4_dec_uops_3_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_ctrl_imm_sel <= io_enq_4_dec_uops_3_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_ctrl_op_fcn <= io_enq_4_dec_uops_3_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_ctrl_fcn_dw <= io_enq_4_dec_uops_3_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_ctrl_csr_cmd <= io_enq_4_dec_uops_3_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_ctrl_is_load <= io_enq_4_dec_uops_3_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_ctrl_is_sta <= io_enq_4_dec_uops_3_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_ctrl_is_std <= io_enq_4_dec_uops_3_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_ctrl_op3_sel <= io_enq_4_dec_uops_3_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_iw_state <= io_enq_4_dec_uops_3_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_iw_p1_poisoned <= io_enq_4_dec_uops_3_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_iw_p2_poisoned <= io_enq_4_dec_uops_3_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_is_br <= io_enq_4_dec_uops_3_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_is_jalr <= io_enq_4_dec_uops_3_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_is_jal <= io_enq_4_dec_uops_3_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_is_sfb <= io_enq_4_dec_uops_3_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_br_mask <= io_enq_4_dec_uops_3_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_br_tag <= io_enq_4_dec_uops_3_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_ftq_idx <= io_enq_4_dec_uops_3_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_edge_inst <= io_enq_4_dec_uops_3_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_pc_lob <= io_enq_4_dec_uops_3_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_taken <= io_enq_4_dec_uops_3_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_imm_packed <= io_enq_4_dec_uops_3_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_csr_addr <= io_enq_4_dec_uops_3_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_rob_idx <= io_enq_4_dec_uops_3_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_ldq_idx <= io_enq_4_dec_uops_3_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_stq_idx <= io_enq_4_dec_uops_3_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_rxq_idx <= io_enq_4_dec_uops_3_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_pdst <= io_enq_4_dec_uops_3_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_prs1 <= io_enq_4_dec_uops_3_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_prs2 <= io_enq_4_dec_uops_3_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_prs3 <= io_enq_4_dec_uops_3_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_ppred <= io_enq_4_dec_uops_3_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_prs1_busy <= io_enq_4_dec_uops_3_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_prs2_busy <= io_enq_4_dec_uops_3_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_prs3_busy <= io_enq_4_dec_uops_3_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_ppred_busy <= io_enq_4_dec_uops_3_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_stale_pdst <= io_enq_4_dec_uops_3_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_exception <= io_enq_4_dec_uops_3_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_exc_cause <= io_enq_4_dec_uops_3_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_bypassable <= io_enq_4_dec_uops_3_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_mem_cmd <= io_enq_4_dec_uops_3_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_mem_size <= io_enq_4_dec_uops_3_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_mem_signed <= io_enq_4_dec_uops_3_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_is_fence <= io_enq_4_dec_uops_3_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_is_fencei <= io_enq_4_dec_uops_3_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_is_amo <= io_enq_4_dec_uops_3_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_uses_ldq <= io_enq_4_dec_uops_3_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_uses_stq <= io_enq_4_dec_uops_3_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_is_sys_pc2epc <= io_enq_4_dec_uops_3_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_is_unique <= io_enq_4_dec_uops_3_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_flush_on_commit <= io_enq_4_dec_uops_3_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_ldst_is_rs1 <= io_enq_4_dec_uops_3_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_ldst <= io_enq_4_dec_uops_3_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_lrs1 <= io_enq_4_dec_uops_3_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_lrs2 <= io_enq_4_dec_uops_3_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_lrs3 <= io_enq_4_dec_uops_3_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_ldst_val <= io_enq_4_dec_uops_3_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_dst_rtype <= io_enq_4_dec_uops_3_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_lrs1_rtype <= io_enq_4_dec_uops_3_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_lrs2_rtype <= io_enq_4_dec_uops_3_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_frs3_en <= io_enq_4_dec_uops_3_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_fp_val <= io_enq_4_dec_uops_3_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_fp_single <= io_enq_4_dec_uops_3_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_xcpt_pf_if <= io_enq_4_dec_uops_3_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_xcpt_ae_if <= io_enq_4_dec_uops_3_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_xcpt_ma_if <= io_enq_4_dec_uops_3_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_bp_debug_if <= io_enq_4_dec_uops_3_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_bp_xcpt_if <= io_enq_4_dec_uops_3_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_debug_fsrc <= io_enq_4_dec_uops_3_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_dec_uops_3_debug_tsrc <= io_enq_4_dec_uops_3_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_4_val_mask_0 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_val_mask_0 <= io_enq_4_val_mask_0; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_4_val_mask_1 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_val_mask_1 <= io_enq_4_val_mask_1; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_4_val_mask_2 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_val_mask_2 <= io_enq_4_val_mask_2; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_4_val_mask_3 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_4_val_mask_3 <= io_enq_4_val_mask_3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_switch <= io_enq_5_dec_uops_0_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_switch_off <= io_enq_5_dec_uops_0_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_is_unicore <= io_enq_5_dec_uops_0_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_shift <= io_enq_5_dec_uops_0_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_lrs3_rtype <= io_enq_5_dec_uops_0_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_rflag <= io_enq_5_dec_uops_0_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_wflag <= io_enq_5_dec_uops_0_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_prflag <= io_enq_5_dec_uops_0_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_pwflag <= io_enq_5_dec_uops_0_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_pflag_busy <= io_enq_5_dec_uops_0_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_stale_pflag <= io_enq_5_dec_uops_0_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_op1_sel <= io_enq_5_dec_uops_0_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_op2_sel <= io_enq_5_dec_uops_0_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_split_num <= io_enq_5_dec_uops_0_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_self_index <= io_enq_5_dec_uops_0_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_rob_inst_idx <= io_enq_5_dec_uops_0_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_address_num <= io_enq_5_dec_uops_0_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_uopc <= io_enq_5_dec_uops_0_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_inst <= io_enq_5_dec_uops_0_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_debug_inst <= io_enq_5_dec_uops_0_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_is_rvc <= io_enq_5_dec_uops_0_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_debug_pc <= io_enq_5_dec_uops_0_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_iq_type <= io_enq_5_dec_uops_0_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_fu_code <= io_enq_5_dec_uops_0_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_ctrl_br_type <= io_enq_5_dec_uops_0_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_ctrl_op1_sel <= io_enq_5_dec_uops_0_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_ctrl_op2_sel <= io_enq_5_dec_uops_0_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_ctrl_imm_sel <= io_enq_5_dec_uops_0_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_ctrl_op_fcn <= io_enq_5_dec_uops_0_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_ctrl_fcn_dw <= io_enq_5_dec_uops_0_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_ctrl_csr_cmd <= io_enq_5_dec_uops_0_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_ctrl_is_load <= io_enq_5_dec_uops_0_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_ctrl_is_sta <= io_enq_5_dec_uops_0_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_ctrl_is_std <= io_enq_5_dec_uops_0_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_ctrl_op3_sel <= io_enq_5_dec_uops_0_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_iw_state <= io_enq_5_dec_uops_0_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_iw_p1_poisoned <= io_enq_5_dec_uops_0_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_iw_p2_poisoned <= io_enq_5_dec_uops_0_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_is_br <= io_enq_5_dec_uops_0_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_is_jalr <= io_enq_5_dec_uops_0_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_is_jal <= io_enq_5_dec_uops_0_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_is_sfb <= io_enq_5_dec_uops_0_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_br_mask <= io_enq_5_dec_uops_0_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_br_tag <= io_enq_5_dec_uops_0_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_ftq_idx <= io_enq_5_dec_uops_0_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_edge_inst <= io_enq_5_dec_uops_0_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_pc_lob <= io_enq_5_dec_uops_0_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_taken <= io_enq_5_dec_uops_0_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_imm_packed <= io_enq_5_dec_uops_0_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_csr_addr <= io_enq_5_dec_uops_0_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_rob_idx <= io_enq_5_dec_uops_0_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_ldq_idx <= io_enq_5_dec_uops_0_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_stq_idx <= io_enq_5_dec_uops_0_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_rxq_idx <= io_enq_5_dec_uops_0_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_pdst <= io_enq_5_dec_uops_0_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_prs1 <= io_enq_5_dec_uops_0_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_prs2 <= io_enq_5_dec_uops_0_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_prs3 <= io_enq_5_dec_uops_0_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_ppred <= io_enq_5_dec_uops_0_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_prs1_busy <= io_enq_5_dec_uops_0_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_prs2_busy <= io_enq_5_dec_uops_0_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_prs3_busy <= io_enq_5_dec_uops_0_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_ppred_busy <= io_enq_5_dec_uops_0_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_stale_pdst <= io_enq_5_dec_uops_0_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_exception <= io_enq_5_dec_uops_0_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_exc_cause <= io_enq_5_dec_uops_0_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_bypassable <= io_enq_5_dec_uops_0_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_mem_cmd <= io_enq_5_dec_uops_0_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_mem_size <= io_enq_5_dec_uops_0_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_mem_signed <= io_enq_5_dec_uops_0_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_is_fence <= io_enq_5_dec_uops_0_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_is_fencei <= io_enq_5_dec_uops_0_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_is_amo <= io_enq_5_dec_uops_0_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_uses_ldq <= io_enq_5_dec_uops_0_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_uses_stq <= io_enq_5_dec_uops_0_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_is_sys_pc2epc <= io_enq_5_dec_uops_0_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_is_unique <= io_enq_5_dec_uops_0_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_flush_on_commit <= io_enq_5_dec_uops_0_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_ldst_is_rs1 <= io_enq_5_dec_uops_0_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_ldst <= io_enq_5_dec_uops_0_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_lrs1 <= io_enq_5_dec_uops_0_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_lrs2 <= io_enq_5_dec_uops_0_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_lrs3 <= io_enq_5_dec_uops_0_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_ldst_val <= io_enq_5_dec_uops_0_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_dst_rtype <= io_enq_5_dec_uops_0_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_lrs1_rtype <= io_enq_5_dec_uops_0_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_lrs2_rtype <= io_enq_5_dec_uops_0_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_frs3_en <= io_enq_5_dec_uops_0_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_fp_val <= io_enq_5_dec_uops_0_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_fp_single <= io_enq_5_dec_uops_0_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_xcpt_pf_if <= io_enq_5_dec_uops_0_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_xcpt_ae_if <= io_enq_5_dec_uops_0_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_xcpt_ma_if <= io_enq_5_dec_uops_0_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_bp_debug_if <= io_enq_5_dec_uops_0_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_bp_xcpt_if <= io_enq_5_dec_uops_0_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_debug_fsrc <= io_enq_5_dec_uops_0_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_0_debug_tsrc <= io_enq_5_dec_uops_0_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_switch <= io_enq_5_dec_uops_1_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_switch_off <= io_enq_5_dec_uops_1_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_is_unicore <= io_enq_5_dec_uops_1_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_shift <= io_enq_5_dec_uops_1_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_lrs3_rtype <= io_enq_5_dec_uops_1_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_rflag <= io_enq_5_dec_uops_1_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_wflag <= io_enq_5_dec_uops_1_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_prflag <= io_enq_5_dec_uops_1_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_pwflag <= io_enq_5_dec_uops_1_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_pflag_busy <= io_enq_5_dec_uops_1_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_stale_pflag <= io_enq_5_dec_uops_1_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_op1_sel <= io_enq_5_dec_uops_1_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_op2_sel <= io_enq_5_dec_uops_1_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_split_num <= io_enq_5_dec_uops_1_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_self_index <= io_enq_5_dec_uops_1_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_rob_inst_idx <= io_enq_5_dec_uops_1_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_address_num <= io_enq_5_dec_uops_1_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_uopc <= io_enq_5_dec_uops_1_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_inst <= io_enq_5_dec_uops_1_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_debug_inst <= io_enq_5_dec_uops_1_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_is_rvc <= io_enq_5_dec_uops_1_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_debug_pc <= io_enq_5_dec_uops_1_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_iq_type <= io_enq_5_dec_uops_1_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_fu_code <= io_enq_5_dec_uops_1_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_ctrl_br_type <= io_enq_5_dec_uops_1_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_ctrl_op1_sel <= io_enq_5_dec_uops_1_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_ctrl_op2_sel <= io_enq_5_dec_uops_1_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_ctrl_imm_sel <= io_enq_5_dec_uops_1_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_ctrl_op_fcn <= io_enq_5_dec_uops_1_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_ctrl_fcn_dw <= io_enq_5_dec_uops_1_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_ctrl_csr_cmd <= io_enq_5_dec_uops_1_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_ctrl_is_load <= io_enq_5_dec_uops_1_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_ctrl_is_sta <= io_enq_5_dec_uops_1_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_ctrl_is_std <= io_enq_5_dec_uops_1_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_ctrl_op3_sel <= io_enq_5_dec_uops_1_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_iw_state <= io_enq_5_dec_uops_1_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_iw_p1_poisoned <= io_enq_5_dec_uops_1_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_iw_p2_poisoned <= io_enq_5_dec_uops_1_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_is_br <= io_enq_5_dec_uops_1_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_is_jalr <= io_enq_5_dec_uops_1_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_is_jal <= io_enq_5_dec_uops_1_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_is_sfb <= io_enq_5_dec_uops_1_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_br_mask <= io_enq_5_dec_uops_1_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_br_tag <= io_enq_5_dec_uops_1_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_ftq_idx <= io_enq_5_dec_uops_1_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_edge_inst <= io_enq_5_dec_uops_1_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_pc_lob <= io_enq_5_dec_uops_1_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_taken <= io_enq_5_dec_uops_1_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_imm_packed <= io_enq_5_dec_uops_1_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_csr_addr <= io_enq_5_dec_uops_1_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_rob_idx <= io_enq_5_dec_uops_1_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_ldq_idx <= io_enq_5_dec_uops_1_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_stq_idx <= io_enq_5_dec_uops_1_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_rxq_idx <= io_enq_5_dec_uops_1_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_pdst <= io_enq_5_dec_uops_1_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_prs1 <= io_enq_5_dec_uops_1_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_prs2 <= io_enq_5_dec_uops_1_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_prs3 <= io_enq_5_dec_uops_1_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_ppred <= io_enq_5_dec_uops_1_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_prs1_busy <= io_enq_5_dec_uops_1_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_prs2_busy <= io_enq_5_dec_uops_1_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_prs3_busy <= io_enq_5_dec_uops_1_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_ppred_busy <= io_enq_5_dec_uops_1_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_stale_pdst <= io_enq_5_dec_uops_1_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_exception <= io_enq_5_dec_uops_1_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_exc_cause <= io_enq_5_dec_uops_1_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_bypassable <= io_enq_5_dec_uops_1_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_mem_cmd <= io_enq_5_dec_uops_1_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_mem_size <= io_enq_5_dec_uops_1_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_mem_signed <= io_enq_5_dec_uops_1_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_is_fence <= io_enq_5_dec_uops_1_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_is_fencei <= io_enq_5_dec_uops_1_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_is_amo <= io_enq_5_dec_uops_1_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_uses_ldq <= io_enq_5_dec_uops_1_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_uses_stq <= io_enq_5_dec_uops_1_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_is_sys_pc2epc <= io_enq_5_dec_uops_1_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_is_unique <= io_enq_5_dec_uops_1_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_flush_on_commit <= io_enq_5_dec_uops_1_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_ldst_is_rs1 <= io_enq_5_dec_uops_1_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_ldst <= io_enq_5_dec_uops_1_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_lrs1 <= io_enq_5_dec_uops_1_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_lrs2 <= io_enq_5_dec_uops_1_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_lrs3 <= io_enq_5_dec_uops_1_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_ldst_val <= io_enq_5_dec_uops_1_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_dst_rtype <= io_enq_5_dec_uops_1_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_lrs1_rtype <= io_enq_5_dec_uops_1_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_lrs2_rtype <= io_enq_5_dec_uops_1_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_frs3_en <= io_enq_5_dec_uops_1_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_fp_val <= io_enq_5_dec_uops_1_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_fp_single <= io_enq_5_dec_uops_1_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_xcpt_pf_if <= io_enq_5_dec_uops_1_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_xcpt_ae_if <= io_enq_5_dec_uops_1_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_xcpt_ma_if <= io_enq_5_dec_uops_1_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_bp_debug_if <= io_enq_5_dec_uops_1_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_bp_xcpt_if <= io_enq_5_dec_uops_1_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_debug_fsrc <= io_enq_5_dec_uops_1_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_1_debug_tsrc <= io_enq_5_dec_uops_1_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_switch <= io_enq_5_dec_uops_2_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_switch_off <= io_enq_5_dec_uops_2_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_is_unicore <= io_enq_5_dec_uops_2_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_shift <= io_enq_5_dec_uops_2_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_lrs3_rtype <= io_enq_5_dec_uops_2_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_rflag <= io_enq_5_dec_uops_2_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_wflag <= io_enq_5_dec_uops_2_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_prflag <= io_enq_5_dec_uops_2_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_pwflag <= io_enq_5_dec_uops_2_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_pflag_busy <= io_enq_5_dec_uops_2_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_stale_pflag <= io_enq_5_dec_uops_2_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_op1_sel <= io_enq_5_dec_uops_2_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_op2_sel <= io_enq_5_dec_uops_2_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_split_num <= io_enq_5_dec_uops_2_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_self_index <= io_enq_5_dec_uops_2_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_rob_inst_idx <= io_enq_5_dec_uops_2_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_address_num <= io_enq_5_dec_uops_2_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_uopc <= io_enq_5_dec_uops_2_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_inst <= io_enq_5_dec_uops_2_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_debug_inst <= io_enq_5_dec_uops_2_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_is_rvc <= io_enq_5_dec_uops_2_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_debug_pc <= io_enq_5_dec_uops_2_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_iq_type <= io_enq_5_dec_uops_2_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_fu_code <= io_enq_5_dec_uops_2_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_ctrl_br_type <= io_enq_5_dec_uops_2_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_ctrl_op1_sel <= io_enq_5_dec_uops_2_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_ctrl_op2_sel <= io_enq_5_dec_uops_2_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_ctrl_imm_sel <= io_enq_5_dec_uops_2_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_ctrl_op_fcn <= io_enq_5_dec_uops_2_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_ctrl_fcn_dw <= io_enq_5_dec_uops_2_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_ctrl_csr_cmd <= io_enq_5_dec_uops_2_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_ctrl_is_load <= io_enq_5_dec_uops_2_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_ctrl_is_sta <= io_enq_5_dec_uops_2_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_ctrl_is_std <= io_enq_5_dec_uops_2_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_ctrl_op3_sel <= io_enq_5_dec_uops_2_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_iw_state <= io_enq_5_dec_uops_2_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_iw_p1_poisoned <= io_enq_5_dec_uops_2_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_iw_p2_poisoned <= io_enq_5_dec_uops_2_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_is_br <= io_enq_5_dec_uops_2_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_is_jalr <= io_enq_5_dec_uops_2_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_is_jal <= io_enq_5_dec_uops_2_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_is_sfb <= io_enq_5_dec_uops_2_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_br_mask <= io_enq_5_dec_uops_2_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_br_tag <= io_enq_5_dec_uops_2_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_ftq_idx <= io_enq_5_dec_uops_2_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_edge_inst <= io_enq_5_dec_uops_2_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_pc_lob <= io_enq_5_dec_uops_2_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_taken <= io_enq_5_dec_uops_2_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_imm_packed <= io_enq_5_dec_uops_2_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_csr_addr <= io_enq_5_dec_uops_2_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_rob_idx <= io_enq_5_dec_uops_2_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_ldq_idx <= io_enq_5_dec_uops_2_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_stq_idx <= io_enq_5_dec_uops_2_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_rxq_idx <= io_enq_5_dec_uops_2_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_pdst <= io_enq_5_dec_uops_2_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_prs1 <= io_enq_5_dec_uops_2_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_prs2 <= io_enq_5_dec_uops_2_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_prs3 <= io_enq_5_dec_uops_2_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_ppred <= io_enq_5_dec_uops_2_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_prs1_busy <= io_enq_5_dec_uops_2_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_prs2_busy <= io_enq_5_dec_uops_2_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_prs3_busy <= io_enq_5_dec_uops_2_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_ppred_busy <= io_enq_5_dec_uops_2_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_stale_pdst <= io_enq_5_dec_uops_2_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_exception <= io_enq_5_dec_uops_2_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_exc_cause <= io_enq_5_dec_uops_2_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_bypassable <= io_enq_5_dec_uops_2_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_mem_cmd <= io_enq_5_dec_uops_2_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_mem_size <= io_enq_5_dec_uops_2_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_mem_signed <= io_enq_5_dec_uops_2_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_is_fence <= io_enq_5_dec_uops_2_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_is_fencei <= io_enq_5_dec_uops_2_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_is_amo <= io_enq_5_dec_uops_2_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_uses_ldq <= io_enq_5_dec_uops_2_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_uses_stq <= io_enq_5_dec_uops_2_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_is_sys_pc2epc <= io_enq_5_dec_uops_2_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_is_unique <= io_enq_5_dec_uops_2_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_flush_on_commit <= io_enq_5_dec_uops_2_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_ldst_is_rs1 <= io_enq_5_dec_uops_2_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_ldst <= io_enq_5_dec_uops_2_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_lrs1 <= io_enq_5_dec_uops_2_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_lrs2 <= io_enq_5_dec_uops_2_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_lrs3 <= io_enq_5_dec_uops_2_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_ldst_val <= io_enq_5_dec_uops_2_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_dst_rtype <= io_enq_5_dec_uops_2_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_lrs1_rtype <= io_enq_5_dec_uops_2_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_lrs2_rtype <= io_enq_5_dec_uops_2_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_frs3_en <= io_enq_5_dec_uops_2_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_fp_val <= io_enq_5_dec_uops_2_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_fp_single <= io_enq_5_dec_uops_2_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_xcpt_pf_if <= io_enq_5_dec_uops_2_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_xcpt_ae_if <= io_enq_5_dec_uops_2_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_xcpt_ma_if <= io_enq_5_dec_uops_2_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_bp_debug_if <= io_enq_5_dec_uops_2_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_bp_xcpt_if <= io_enq_5_dec_uops_2_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_debug_fsrc <= io_enq_5_dec_uops_2_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_2_debug_tsrc <= io_enq_5_dec_uops_2_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_switch <= io_enq_5_dec_uops_3_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_switch_off <= io_enq_5_dec_uops_3_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_is_unicore <= io_enq_5_dec_uops_3_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_shift <= io_enq_5_dec_uops_3_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_lrs3_rtype <= io_enq_5_dec_uops_3_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_rflag <= io_enq_5_dec_uops_3_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_wflag <= io_enq_5_dec_uops_3_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_prflag <= io_enq_5_dec_uops_3_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_pwflag <= io_enq_5_dec_uops_3_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_pflag_busy <= io_enq_5_dec_uops_3_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_stale_pflag <= io_enq_5_dec_uops_3_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_op1_sel <= io_enq_5_dec_uops_3_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_op2_sel <= io_enq_5_dec_uops_3_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_split_num <= io_enq_5_dec_uops_3_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_self_index <= io_enq_5_dec_uops_3_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_rob_inst_idx <= io_enq_5_dec_uops_3_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_address_num <= io_enq_5_dec_uops_3_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_uopc <= io_enq_5_dec_uops_3_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_inst <= io_enq_5_dec_uops_3_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_debug_inst <= io_enq_5_dec_uops_3_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_is_rvc <= io_enq_5_dec_uops_3_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_debug_pc <= io_enq_5_dec_uops_3_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_iq_type <= io_enq_5_dec_uops_3_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_fu_code <= io_enq_5_dec_uops_3_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_ctrl_br_type <= io_enq_5_dec_uops_3_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_ctrl_op1_sel <= io_enq_5_dec_uops_3_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_ctrl_op2_sel <= io_enq_5_dec_uops_3_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_ctrl_imm_sel <= io_enq_5_dec_uops_3_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_ctrl_op_fcn <= io_enq_5_dec_uops_3_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_ctrl_fcn_dw <= io_enq_5_dec_uops_3_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_ctrl_csr_cmd <= io_enq_5_dec_uops_3_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_ctrl_is_load <= io_enq_5_dec_uops_3_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_ctrl_is_sta <= io_enq_5_dec_uops_3_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_ctrl_is_std <= io_enq_5_dec_uops_3_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_ctrl_op3_sel <= io_enq_5_dec_uops_3_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_iw_state <= io_enq_5_dec_uops_3_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_iw_p1_poisoned <= io_enq_5_dec_uops_3_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_iw_p2_poisoned <= io_enq_5_dec_uops_3_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_is_br <= io_enq_5_dec_uops_3_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_is_jalr <= io_enq_5_dec_uops_3_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_is_jal <= io_enq_5_dec_uops_3_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_is_sfb <= io_enq_5_dec_uops_3_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_br_mask <= io_enq_5_dec_uops_3_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_br_tag <= io_enq_5_dec_uops_3_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_ftq_idx <= io_enq_5_dec_uops_3_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_edge_inst <= io_enq_5_dec_uops_3_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_pc_lob <= io_enq_5_dec_uops_3_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_taken <= io_enq_5_dec_uops_3_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_imm_packed <= io_enq_5_dec_uops_3_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_csr_addr <= io_enq_5_dec_uops_3_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_rob_idx <= io_enq_5_dec_uops_3_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_ldq_idx <= io_enq_5_dec_uops_3_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_stq_idx <= io_enq_5_dec_uops_3_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_rxq_idx <= io_enq_5_dec_uops_3_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_pdst <= io_enq_5_dec_uops_3_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_prs1 <= io_enq_5_dec_uops_3_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_prs2 <= io_enq_5_dec_uops_3_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_prs3 <= io_enq_5_dec_uops_3_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_ppred <= io_enq_5_dec_uops_3_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_prs1_busy <= io_enq_5_dec_uops_3_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_prs2_busy <= io_enq_5_dec_uops_3_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_prs3_busy <= io_enq_5_dec_uops_3_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_ppred_busy <= io_enq_5_dec_uops_3_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_stale_pdst <= io_enq_5_dec_uops_3_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_exception <= io_enq_5_dec_uops_3_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_exc_cause <= io_enq_5_dec_uops_3_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_bypassable <= io_enq_5_dec_uops_3_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_mem_cmd <= io_enq_5_dec_uops_3_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_mem_size <= io_enq_5_dec_uops_3_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_mem_signed <= io_enq_5_dec_uops_3_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_is_fence <= io_enq_5_dec_uops_3_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_is_fencei <= io_enq_5_dec_uops_3_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_is_amo <= io_enq_5_dec_uops_3_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_uses_ldq <= io_enq_5_dec_uops_3_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_uses_stq <= io_enq_5_dec_uops_3_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_is_sys_pc2epc <= io_enq_5_dec_uops_3_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_is_unique <= io_enq_5_dec_uops_3_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_flush_on_commit <= io_enq_5_dec_uops_3_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_ldst_is_rs1 <= io_enq_5_dec_uops_3_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_ldst <= io_enq_5_dec_uops_3_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_lrs1 <= io_enq_5_dec_uops_3_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_lrs2 <= io_enq_5_dec_uops_3_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_lrs3 <= io_enq_5_dec_uops_3_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_ldst_val <= io_enq_5_dec_uops_3_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_dst_rtype <= io_enq_5_dec_uops_3_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_lrs1_rtype <= io_enq_5_dec_uops_3_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_lrs2_rtype <= io_enq_5_dec_uops_3_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_frs3_en <= io_enq_5_dec_uops_3_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_fp_val <= io_enq_5_dec_uops_3_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_fp_single <= io_enq_5_dec_uops_3_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_xcpt_pf_if <= io_enq_5_dec_uops_3_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_xcpt_ae_if <= io_enq_5_dec_uops_3_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_xcpt_ma_if <= io_enq_5_dec_uops_3_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_bp_debug_if <= io_enq_5_dec_uops_3_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_bp_xcpt_if <= io_enq_5_dec_uops_3_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_debug_fsrc <= io_enq_5_dec_uops_3_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_dec_uops_3_debug_tsrc <= io_enq_5_dec_uops_3_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_5_val_mask_0 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_val_mask_0 <= io_enq_5_val_mask_0; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_5_val_mask_1 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_val_mask_1 <= io_enq_5_val_mask_1; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_5_val_mask_2 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_val_mask_2 <= io_enq_5_val_mask_2; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_5_val_mask_3 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_5_val_mask_3 <= io_enq_5_val_mask_3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_switch <= io_enq_6_dec_uops_0_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_switch_off <= io_enq_6_dec_uops_0_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_is_unicore <= io_enq_6_dec_uops_0_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_shift <= io_enq_6_dec_uops_0_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_lrs3_rtype <= io_enq_6_dec_uops_0_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_rflag <= io_enq_6_dec_uops_0_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_wflag <= io_enq_6_dec_uops_0_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_prflag <= io_enq_6_dec_uops_0_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_pwflag <= io_enq_6_dec_uops_0_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_pflag_busy <= io_enq_6_dec_uops_0_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_stale_pflag <= io_enq_6_dec_uops_0_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_op1_sel <= io_enq_6_dec_uops_0_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_op2_sel <= io_enq_6_dec_uops_0_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_split_num <= io_enq_6_dec_uops_0_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_self_index <= io_enq_6_dec_uops_0_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_rob_inst_idx <= io_enq_6_dec_uops_0_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_address_num <= io_enq_6_dec_uops_0_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_uopc <= io_enq_6_dec_uops_0_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_inst <= io_enq_6_dec_uops_0_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_debug_inst <= io_enq_6_dec_uops_0_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_is_rvc <= io_enq_6_dec_uops_0_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_debug_pc <= io_enq_6_dec_uops_0_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_iq_type <= io_enq_6_dec_uops_0_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_fu_code <= io_enq_6_dec_uops_0_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_ctrl_br_type <= io_enq_6_dec_uops_0_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_ctrl_op1_sel <= io_enq_6_dec_uops_0_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_ctrl_op2_sel <= io_enq_6_dec_uops_0_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_ctrl_imm_sel <= io_enq_6_dec_uops_0_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_ctrl_op_fcn <= io_enq_6_dec_uops_0_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_ctrl_fcn_dw <= io_enq_6_dec_uops_0_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_ctrl_csr_cmd <= io_enq_6_dec_uops_0_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_ctrl_is_load <= io_enq_6_dec_uops_0_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_ctrl_is_sta <= io_enq_6_dec_uops_0_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_ctrl_is_std <= io_enq_6_dec_uops_0_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_ctrl_op3_sel <= io_enq_6_dec_uops_0_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_iw_state <= io_enq_6_dec_uops_0_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_iw_p1_poisoned <= io_enq_6_dec_uops_0_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_iw_p2_poisoned <= io_enq_6_dec_uops_0_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_is_br <= io_enq_6_dec_uops_0_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_is_jalr <= io_enq_6_dec_uops_0_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_is_jal <= io_enq_6_dec_uops_0_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_is_sfb <= io_enq_6_dec_uops_0_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_br_mask <= io_enq_6_dec_uops_0_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_br_tag <= io_enq_6_dec_uops_0_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_ftq_idx <= io_enq_6_dec_uops_0_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_edge_inst <= io_enq_6_dec_uops_0_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_pc_lob <= io_enq_6_dec_uops_0_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_taken <= io_enq_6_dec_uops_0_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_imm_packed <= io_enq_6_dec_uops_0_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_csr_addr <= io_enq_6_dec_uops_0_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_rob_idx <= io_enq_6_dec_uops_0_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_ldq_idx <= io_enq_6_dec_uops_0_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_stq_idx <= io_enq_6_dec_uops_0_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_rxq_idx <= io_enq_6_dec_uops_0_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_pdst <= io_enq_6_dec_uops_0_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_prs1 <= io_enq_6_dec_uops_0_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_prs2 <= io_enq_6_dec_uops_0_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_prs3 <= io_enq_6_dec_uops_0_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_ppred <= io_enq_6_dec_uops_0_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_prs1_busy <= io_enq_6_dec_uops_0_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_prs2_busy <= io_enq_6_dec_uops_0_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_prs3_busy <= io_enq_6_dec_uops_0_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_ppred_busy <= io_enq_6_dec_uops_0_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_stale_pdst <= io_enq_6_dec_uops_0_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_exception <= io_enq_6_dec_uops_0_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_exc_cause <= io_enq_6_dec_uops_0_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_bypassable <= io_enq_6_dec_uops_0_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_mem_cmd <= io_enq_6_dec_uops_0_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_mem_size <= io_enq_6_dec_uops_0_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_mem_signed <= io_enq_6_dec_uops_0_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_is_fence <= io_enq_6_dec_uops_0_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_is_fencei <= io_enq_6_dec_uops_0_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_is_amo <= io_enq_6_dec_uops_0_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_uses_ldq <= io_enq_6_dec_uops_0_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_uses_stq <= io_enq_6_dec_uops_0_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_is_sys_pc2epc <= io_enq_6_dec_uops_0_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_is_unique <= io_enq_6_dec_uops_0_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_flush_on_commit <= io_enq_6_dec_uops_0_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_ldst_is_rs1 <= io_enq_6_dec_uops_0_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_ldst <= io_enq_6_dec_uops_0_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_lrs1 <= io_enq_6_dec_uops_0_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_lrs2 <= io_enq_6_dec_uops_0_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_lrs3 <= io_enq_6_dec_uops_0_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_ldst_val <= io_enq_6_dec_uops_0_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_dst_rtype <= io_enq_6_dec_uops_0_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_lrs1_rtype <= io_enq_6_dec_uops_0_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_lrs2_rtype <= io_enq_6_dec_uops_0_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_frs3_en <= io_enq_6_dec_uops_0_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_fp_val <= io_enq_6_dec_uops_0_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_fp_single <= io_enq_6_dec_uops_0_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_xcpt_pf_if <= io_enq_6_dec_uops_0_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_xcpt_ae_if <= io_enq_6_dec_uops_0_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_xcpt_ma_if <= io_enq_6_dec_uops_0_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_bp_debug_if <= io_enq_6_dec_uops_0_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_bp_xcpt_if <= io_enq_6_dec_uops_0_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_debug_fsrc <= io_enq_6_dec_uops_0_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_0_debug_tsrc <= io_enq_6_dec_uops_0_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_switch <= io_enq_6_dec_uops_1_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_switch_off <= io_enq_6_dec_uops_1_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_is_unicore <= io_enq_6_dec_uops_1_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_shift <= io_enq_6_dec_uops_1_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_lrs3_rtype <= io_enq_6_dec_uops_1_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_rflag <= io_enq_6_dec_uops_1_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_wflag <= io_enq_6_dec_uops_1_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_prflag <= io_enq_6_dec_uops_1_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_pwflag <= io_enq_6_dec_uops_1_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_pflag_busy <= io_enq_6_dec_uops_1_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_stale_pflag <= io_enq_6_dec_uops_1_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_op1_sel <= io_enq_6_dec_uops_1_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_op2_sel <= io_enq_6_dec_uops_1_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_split_num <= io_enq_6_dec_uops_1_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_self_index <= io_enq_6_dec_uops_1_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_rob_inst_idx <= io_enq_6_dec_uops_1_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_address_num <= io_enq_6_dec_uops_1_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_uopc <= io_enq_6_dec_uops_1_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_inst <= io_enq_6_dec_uops_1_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_debug_inst <= io_enq_6_dec_uops_1_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_is_rvc <= io_enq_6_dec_uops_1_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_debug_pc <= io_enq_6_dec_uops_1_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_iq_type <= io_enq_6_dec_uops_1_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_fu_code <= io_enq_6_dec_uops_1_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_ctrl_br_type <= io_enq_6_dec_uops_1_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_ctrl_op1_sel <= io_enq_6_dec_uops_1_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_ctrl_op2_sel <= io_enq_6_dec_uops_1_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_ctrl_imm_sel <= io_enq_6_dec_uops_1_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_ctrl_op_fcn <= io_enq_6_dec_uops_1_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_ctrl_fcn_dw <= io_enq_6_dec_uops_1_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_ctrl_csr_cmd <= io_enq_6_dec_uops_1_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_ctrl_is_load <= io_enq_6_dec_uops_1_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_ctrl_is_sta <= io_enq_6_dec_uops_1_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_ctrl_is_std <= io_enq_6_dec_uops_1_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_ctrl_op3_sel <= io_enq_6_dec_uops_1_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_iw_state <= io_enq_6_dec_uops_1_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_iw_p1_poisoned <= io_enq_6_dec_uops_1_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_iw_p2_poisoned <= io_enq_6_dec_uops_1_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_is_br <= io_enq_6_dec_uops_1_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_is_jalr <= io_enq_6_dec_uops_1_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_is_jal <= io_enq_6_dec_uops_1_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_is_sfb <= io_enq_6_dec_uops_1_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_br_mask <= io_enq_6_dec_uops_1_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_br_tag <= io_enq_6_dec_uops_1_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_ftq_idx <= io_enq_6_dec_uops_1_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_edge_inst <= io_enq_6_dec_uops_1_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_pc_lob <= io_enq_6_dec_uops_1_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_taken <= io_enq_6_dec_uops_1_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_imm_packed <= io_enq_6_dec_uops_1_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_csr_addr <= io_enq_6_dec_uops_1_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_rob_idx <= io_enq_6_dec_uops_1_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_ldq_idx <= io_enq_6_dec_uops_1_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_stq_idx <= io_enq_6_dec_uops_1_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_rxq_idx <= io_enq_6_dec_uops_1_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_pdst <= io_enq_6_dec_uops_1_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_prs1 <= io_enq_6_dec_uops_1_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_prs2 <= io_enq_6_dec_uops_1_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_prs3 <= io_enq_6_dec_uops_1_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_ppred <= io_enq_6_dec_uops_1_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_prs1_busy <= io_enq_6_dec_uops_1_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_prs2_busy <= io_enq_6_dec_uops_1_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_prs3_busy <= io_enq_6_dec_uops_1_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_ppred_busy <= io_enq_6_dec_uops_1_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_stale_pdst <= io_enq_6_dec_uops_1_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_exception <= io_enq_6_dec_uops_1_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_exc_cause <= io_enq_6_dec_uops_1_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_bypassable <= io_enq_6_dec_uops_1_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_mem_cmd <= io_enq_6_dec_uops_1_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_mem_size <= io_enq_6_dec_uops_1_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_mem_signed <= io_enq_6_dec_uops_1_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_is_fence <= io_enq_6_dec_uops_1_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_is_fencei <= io_enq_6_dec_uops_1_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_is_amo <= io_enq_6_dec_uops_1_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_uses_ldq <= io_enq_6_dec_uops_1_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_uses_stq <= io_enq_6_dec_uops_1_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_is_sys_pc2epc <= io_enq_6_dec_uops_1_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_is_unique <= io_enq_6_dec_uops_1_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_flush_on_commit <= io_enq_6_dec_uops_1_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_ldst_is_rs1 <= io_enq_6_dec_uops_1_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_ldst <= io_enq_6_dec_uops_1_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_lrs1 <= io_enq_6_dec_uops_1_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_lrs2 <= io_enq_6_dec_uops_1_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_lrs3 <= io_enq_6_dec_uops_1_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_ldst_val <= io_enq_6_dec_uops_1_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_dst_rtype <= io_enq_6_dec_uops_1_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_lrs1_rtype <= io_enq_6_dec_uops_1_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_lrs2_rtype <= io_enq_6_dec_uops_1_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_frs3_en <= io_enq_6_dec_uops_1_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_fp_val <= io_enq_6_dec_uops_1_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_fp_single <= io_enq_6_dec_uops_1_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_xcpt_pf_if <= io_enq_6_dec_uops_1_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_xcpt_ae_if <= io_enq_6_dec_uops_1_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_xcpt_ma_if <= io_enq_6_dec_uops_1_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_bp_debug_if <= io_enq_6_dec_uops_1_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_bp_xcpt_if <= io_enq_6_dec_uops_1_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_debug_fsrc <= io_enq_6_dec_uops_1_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_1_debug_tsrc <= io_enq_6_dec_uops_1_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_switch <= io_enq_6_dec_uops_2_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_switch_off <= io_enq_6_dec_uops_2_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_is_unicore <= io_enq_6_dec_uops_2_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_shift <= io_enq_6_dec_uops_2_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_lrs3_rtype <= io_enq_6_dec_uops_2_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_rflag <= io_enq_6_dec_uops_2_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_wflag <= io_enq_6_dec_uops_2_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_prflag <= io_enq_6_dec_uops_2_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_pwflag <= io_enq_6_dec_uops_2_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_pflag_busy <= io_enq_6_dec_uops_2_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_stale_pflag <= io_enq_6_dec_uops_2_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_op1_sel <= io_enq_6_dec_uops_2_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_op2_sel <= io_enq_6_dec_uops_2_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_split_num <= io_enq_6_dec_uops_2_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_self_index <= io_enq_6_dec_uops_2_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_rob_inst_idx <= io_enq_6_dec_uops_2_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_address_num <= io_enq_6_dec_uops_2_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_uopc <= io_enq_6_dec_uops_2_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_inst <= io_enq_6_dec_uops_2_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_debug_inst <= io_enq_6_dec_uops_2_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_is_rvc <= io_enq_6_dec_uops_2_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_debug_pc <= io_enq_6_dec_uops_2_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_iq_type <= io_enq_6_dec_uops_2_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_fu_code <= io_enq_6_dec_uops_2_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_ctrl_br_type <= io_enq_6_dec_uops_2_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_ctrl_op1_sel <= io_enq_6_dec_uops_2_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_ctrl_op2_sel <= io_enq_6_dec_uops_2_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_ctrl_imm_sel <= io_enq_6_dec_uops_2_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_ctrl_op_fcn <= io_enq_6_dec_uops_2_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_ctrl_fcn_dw <= io_enq_6_dec_uops_2_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_ctrl_csr_cmd <= io_enq_6_dec_uops_2_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_ctrl_is_load <= io_enq_6_dec_uops_2_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_ctrl_is_sta <= io_enq_6_dec_uops_2_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_ctrl_is_std <= io_enq_6_dec_uops_2_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_ctrl_op3_sel <= io_enq_6_dec_uops_2_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_iw_state <= io_enq_6_dec_uops_2_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_iw_p1_poisoned <= io_enq_6_dec_uops_2_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_iw_p2_poisoned <= io_enq_6_dec_uops_2_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_is_br <= io_enq_6_dec_uops_2_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_is_jalr <= io_enq_6_dec_uops_2_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_is_jal <= io_enq_6_dec_uops_2_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_is_sfb <= io_enq_6_dec_uops_2_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_br_mask <= io_enq_6_dec_uops_2_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_br_tag <= io_enq_6_dec_uops_2_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_ftq_idx <= io_enq_6_dec_uops_2_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_edge_inst <= io_enq_6_dec_uops_2_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_pc_lob <= io_enq_6_dec_uops_2_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_taken <= io_enq_6_dec_uops_2_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_imm_packed <= io_enq_6_dec_uops_2_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_csr_addr <= io_enq_6_dec_uops_2_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_rob_idx <= io_enq_6_dec_uops_2_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_ldq_idx <= io_enq_6_dec_uops_2_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_stq_idx <= io_enq_6_dec_uops_2_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_rxq_idx <= io_enq_6_dec_uops_2_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_pdst <= io_enq_6_dec_uops_2_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_prs1 <= io_enq_6_dec_uops_2_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_prs2 <= io_enq_6_dec_uops_2_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_prs3 <= io_enq_6_dec_uops_2_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_ppred <= io_enq_6_dec_uops_2_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_prs1_busy <= io_enq_6_dec_uops_2_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_prs2_busy <= io_enq_6_dec_uops_2_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_prs3_busy <= io_enq_6_dec_uops_2_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_ppred_busy <= io_enq_6_dec_uops_2_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_stale_pdst <= io_enq_6_dec_uops_2_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_exception <= io_enq_6_dec_uops_2_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_exc_cause <= io_enq_6_dec_uops_2_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_bypassable <= io_enq_6_dec_uops_2_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_mem_cmd <= io_enq_6_dec_uops_2_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_mem_size <= io_enq_6_dec_uops_2_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_mem_signed <= io_enq_6_dec_uops_2_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_is_fence <= io_enq_6_dec_uops_2_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_is_fencei <= io_enq_6_dec_uops_2_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_is_amo <= io_enq_6_dec_uops_2_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_uses_ldq <= io_enq_6_dec_uops_2_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_uses_stq <= io_enq_6_dec_uops_2_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_is_sys_pc2epc <= io_enq_6_dec_uops_2_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_is_unique <= io_enq_6_dec_uops_2_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_flush_on_commit <= io_enq_6_dec_uops_2_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_ldst_is_rs1 <= io_enq_6_dec_uops_2_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_ldst <= io_enq_6_dec_uops_2_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_lrs1 <= io_enq_6_dec_uops_2_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_lrs2 <= io_enq_6_dec_uops_2_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_lrs3 <= io_enq_6_dec_uops_2_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_ldst_val <= io_enq_6_dec_uops_2_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_dst_rtype <= io_enq_6_dec_uops_2_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_lrs1_rtype <= io_enq_6_dec_uops_2_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_lrs2_rtype <= io_enq_6_dec_uops_2_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_frs3_en <= io_enq_6_dec_uops_2_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_fp_val <= io_enq_6_dec_uops_2_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_fp_single <= io_enq_6_dec_uops_2_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_xcpt_pf_if <= io_enq_6_dec_uops_2_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_xcpt_ae_if <= io_enq_6_dec_uops_2_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_xcpt_ma_if <= io_enq_6_dec_uops_2_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_bp_debug_if <= io_enq_6_dec_uops_2_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_bp_xcpt_if <= io_enq_6_dec_uops_2_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_debug_fsrc <= io_enq_6_dec_uops_2_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_2_debug_tsrc <= io_enq_6_dec_uops_2_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_switch <= io_enq_6_dec_uops_3_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_switch_off <= io_enq_6_dec_uops_3_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_is_unicore <= io_enq_6_dec_uops_3_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_shift <= io_enq_6_dec_uops_3_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_lrs3_rtype <= io_enq_6_dec_uops_3_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_rflag <= io_enq_6_dec_uops_3_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_wflag <= io_enq_6_dec_uops_3_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_prflag <= io_enq_6_dec_uops_3_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_pwflag <= io_enq_6_dec_uops_3_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_pflag_busy <= io_enq_6_dec_uops_3_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_stale_pflag <= io_enq_6_dec_uops_3_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_op1_sel <= io_enq_6_dec_uops_3_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_op2_sel <= io_enq_6_dec_uops_3_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_split_num <= io_enq_6_dec_uops_3_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_self_index <= io_enq_6_dec_uops_3_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_rob_inst_idx <= io_enq_6_dec_uops_3_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_address_num <= io_enq_6_dec_uops_3_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_uopc <= io_enq_6_dec_uops_3_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_inst <= io_enq_6_dec_uops_3_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_debug_inst <= io_enq_6_dec_uops_3_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_is_rvc <= io_enq_6_dec_uops_3_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_debug_pc <= io_enq_6_dec_uops_3_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_iq_type <= io_enq_6_dec_uops_3_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_fu_code <= io_enq_6_dec_uops_3_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_ctrl_br_type <= io_enq_6_dec_uops_3_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_ctrl_op1_sel <= io_enq_6_dec_uops_3_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_ctrl_op2_sel <= io_enq_6_dec_uops_3_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_ctrl_imm_sel <= io_enq_6_dec_uops_3_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_ctrl_op_fcn <= io_enq_6_dec_uops_3_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_ctrl_fcn_dw <= io_enq_6_dec_uops_3_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_ctrl_csr_cmd <= io_enq_6_dec_uops_3_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_ctrl_is_load <= io_enq_6_dec_uops_3_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_ctrl_is_sta <= io_enq_6_dec_uops_3_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_ctrl_is_std <= io_enq_6_dec_uops_3_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_ctrl_op3_sel <= io_enq_6_dec_uops_3_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_iw_state <= io_enq_6_dec_uops_3_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_iw_p1_poisoned <= io_enq_6_dec_uops_3_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_iw_p2_poisoned <= io_enq_6_dec_uops_3_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_is_br <= io_enq_6_dec_uops_3_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_is_jalr <= io_enq_6_dec_uops_3_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_is_jal <= io_enq_6_dec_uops_3_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_is_sfb <= io_enq_6_dec_uops_3_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_br_mask <= io_enq_6_dec_uops_3_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_br_tag <= io_enq_6_dec_uops_3_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_ftq_idx <= io_enq_6_dec_uops_3_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_edge_inst <= io_enq_6_dec_uops_3_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_pc_lob <= io_enq_6_dec_uops_3_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_taken <= io_enq_6_dec_uops_3_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_imm_packed <= io_enq_6_dec_uops_3_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_csr_addr <= io_enq_6_dec_uops_3_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_rob_idx <= io_enq_6_dec_uops_3_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_ldq_idx <= io_enq_6_dec_uops_3_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_stq_idx <= io_enq_6_dec_uops_3_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_rxq_idx <= io_enq_6_dec_uops_3_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_pdst <= io_enq_6_dec_uops_3_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_prs1 <= io_enq_6_dec_uops_3_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_prs2 <= io_enq_6_dec_uops_3_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_prs3 <= io_enq_6_dec_uops_3_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_ppred <= io_enq_6_dec_uops_3_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_prs1_busy <= io_enq_6_dec_uops_3_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_prs2_busy <= io_enq_6_dec_uops_3_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_prs3_busy <= io_enq_6_dec_uops_3_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_ppred_busy <= io_enq_6_dec_uops_3_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_stale_pdst <= io_enq_6_dec_uops_3_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_exception <= io_enq_6_dec_uops_3_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_exc_cause <= io_enq_6_dec_uops_3_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_bypassable <= io_enq_6_dec_uops_3_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_mem_cmd <= io_enq_6_dec_uops_3_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_mem_size <= io_enq_6_dec_uops_3_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_mem_signed <= io_enq_6_dec_uops_3_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_is_fence <= io_enq_6_dec_uops_3_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_is_fencei <= io_enq_6_dec_uops_3_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_is_amo <= io_enq_6_dec_uops_3_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_uses_ldq <= io_enq_6_dec_uops_3_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_uses_stq <= io_enq_6_dec_uops_3_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_is_sys_pc2epc <= io_enq_6_dec_uops_3_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_is_unique <= io_enq_6_dec_uops_3_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_flush_on_commit <= io_enq_6_dec_uops_3_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_ldst_is_rs1 <= io_enq_6_dec_uops_3_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_ldst <= io_enq_6_dec_uops_3_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_lrs1 <= io_enq_6_dec_uops_3_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_lrs2 <= io_enq_6_dec_uops_3_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_lrs3 <= io_enq_6_dec_uops_3_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_ldst_val <= io_enq_6_dec_uops_3_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_dst_rtype <= io_enq_6_dec_uops_3_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_lrs1_rtype <= io_enq_6_dec_uops_3_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_lrs2_rtype <= io_enq_6_dec_uops_3_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_frs3_en <= io_enq_6_dec_uops_3_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_fp_val <= io_enq_6_dec_uops_3_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_fp_single <= io_enq_6_dec_uops_3_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_xcpt_pf_if <= io_enq_6_dec_uops_3_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_xcpt_ae_if <= io_enq_6_dec_uops_3_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_xcpt_ma_if <= io_enq_6_dec_uops_3_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_bp_debug_if <= io_enq_6_dec_uops_3_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_bp_xcpt_if <= io_enq_6_dec_uops_3_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_debug_fsrc <= io_enq_6_dec_uops_3_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_dec_uops_3_debug_tsrc <= io_enq_6_dec_uops_3_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_6_val_mask_0 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_val_mask_0 <= io_enq_6_val_mask_0; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_6_val_mask_1 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_val_mask_1 <= io_enq_6_val_mask_1; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_6_val_mask_2 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_val_mask_2 <= io_enq_6_val_mask_2; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_6_val_mask_3 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_6_val_mask_3 <= io_enq_6_val_mask_3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_switch <= io_enq_7_dec_uops_0_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_switch_off <= io_enq_7_dec_uops_0_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_is_unicore <= io_enq_7_dec_uops_0_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_shift <= io_enq_7_dec_uops_0_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_lrs3_rtype <= io_enq_7_dec_uops_0_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_rflag <= io_enq_7_dec_uops_0_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_wflag <= io_enq_7_dec_uops_0_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_prflag <= io_enq_7_dec_uops_0_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_pwflag <= io_enq_7_dec_uops_0_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_pflag_busy <= io_enq_7_dec_uops_0_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_stale_pflag <= io_enq_7_dec_uops_0_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_op1_sel <= io_enq_7_dec_uops_0_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_op2_sel <= io_enq_7_dec_uops_0_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_split_num <= io_enq_7_dec_uops_0_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_self_index <= io_enq_7_dec_uops_0_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_rob_inst_idx <= io_enq_7_dec_uops_0_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_address_num <= io_enq_7_dec_uops_0_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_uopc <= io_enq_7_dec_uops_0_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_inst <= io_enq_7_dec_uops_0_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_debug_inst <= io_enq_7_dec_uops_0_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_is_rvc <= io_enq_7_dec_uops_0_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_debug_pc <= io_enq_7_dec_uops_0_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_iq_type <= io_enq_7_dec_uops_0_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_fu_code <= io_enq_7_dec_uops_0_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_ctrl_br_type <= io_enq_7_dec_uops_0_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_ctrl_op1_sel <= io_enq_7_dec_uops_0_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_ctrl_op2_sel <= io_enq_7_dec_uops_0_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_ctrl_imm_sel <= io_enq_7_dec_uops_0_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_ctrl_op_fcn <= io_enq_7_dec_uops_0_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_ctrl_fcn_dw <= io_enq_7_dec_uops_0_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_ctrl_csr_cmd <= io_enq_7_dec_uops_0_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_ctrl_is_load <= io_enq_7_dec_uops_0_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_ctrl_is_sta <= io_enq_7_dec_uops_0_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_ctrl_is_std <= io_enq_7_dec_uops_0_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_ctrl_op3_sel <= io_enq_7_dec_uops_0_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_iw_state <= io_enq_7_dec_uops_0_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_iw_p1_poisoned <= io_enq_7_dec_uops_0_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_iw_p2_poisoned <= io_enq_7_dec_uops_0_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_is_br <= io_enq_7_dec_uops_0_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_is_jalr <= io_enq_7_dec_uops_0_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_is_jal <= io_enq_7_dec_uops_0_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_is_sfb <= io_enq_7_dec_uops_0_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_br_mask <= io_enq_7_dec_uops_0_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_br_tag <= io_enq_7_dec_uops_0_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_ftq_idx <= io_enq_7_dec_uops_0_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_edge_inst <= io_enq_7_dec_uops_0_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_pc_lob <= io_enq_7_dec_uops_0_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_taken <= io_enq_7_dec_uops_0_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_imm_packed <= io_enq_7_dec_uops_0_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_csr_addr <= io_enq_7_dec_uops_0_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_rob_idx <= io_enq_7_dec_uops_0_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_ldq_idx <= io_enq_7_dec_uops_0_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_stq_idx <= io_enq_7_dec_uops_0_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_rxq_idx <= io_enq_7_dec_uops_0_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_pdst <= io_enq_7_dec_uops_0_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_prs1 <= io_enq_7_dec_uops_0_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_prs2 <= io_enq_7_dec_uops_0_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_prs3 <= io_enq_7_dec_uops_0_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_ppred <= io_enq_7_dec_uops_0_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_prs1_busy <= io_enq_7_dec_uops_0_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_prs2_busy <= io_enq_7_dec_uops_0_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_prs3_busy <= io_enq_7_dec_uops_0_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_ppred_busy <= io_enq_7_dec_uops_0_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_stale_pdst <= io_enq_7_dec_uops_0_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_exception <= io_enq_7_dec_uops_0_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_exc_cause <= io_enq_7_dec_uops_0_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_bypassable <= io_enq_7_dec_uops_0_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_mem_cmd <= io_enq_7_dec_uops_0_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_mem_size <= io_enq_7_dec_uops_0_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_mem_signed <= io_enq_7_dec_uops_0_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_is_fence <= io_enq_7_dec_uops_0_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_is_fencei <= io_enq_7_dec_uops_0_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_is_amo <= io_enq_7_dec_uops_0_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_uses_ldq <= io_enq_7_dec_uops_0_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_uses_stq <= io_enq_7_dec_uops_0_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_is_sys_pc2epc <= io_enq_7_dec_uops_0_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_is_unique <= io_enq_7_dec_uops_0_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_flush_on_commit <= io_enq_7_dec_uops_0_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_ldst_is_rs1 <= io_enq_7_dec_uops_0_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_ldst <= io_enq_7_dec_uops_0_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_lrs1 <= io_enq_7_dec_uops_0_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_lrs2 <= io_enq_7_dec_uops_0_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_lrs3 <= io_enq_7_dec_uops_0_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_ldst_val <= io_enq_7_dec_uops_0_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_dst_rtype <= io_enq_7_dec_uops_0_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_lrs1_rtype <= io_enq_7_dec_uops_0_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_lrs2_rtype <= io_enq_7_dec_uops_0_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_frs3_en <= io_enq_7_dec_uops_0_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_fp_val <= io_enq_7_dec_uops_0_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_fp_single <= io_enq_7_dec_uops_0_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_xcpt_pf_if <= io_enq_7_dec_uops_0_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_xcpt_ae_if <= io_enq_7_dec_uops_0_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_xcpt_ma_if <= io_enq_7_dec_uops_0_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_bp_debug_if <= io_enq_7_dec_uops_0_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_bp_xcpt_if <= io_enq_7_dec_uops_0_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_debug_fsrc <= io_enq_7_dec_uops_0_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_0_debug_tsrc <= io_enq_7_dec_uops_0_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_switch <= io_enq_7_dec_uops_1_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_switch_off <= io_enq_7_dec_uops_1_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_is_unicore <= io_enq_7_dec_uops_1_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_shift <= io_enq_7_dec_uops_1_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_lrs3_rtype <= io_enq_7_dec_uops_1_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_rflag <= io_enq_7_dec_uops_1_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_wflag <= io_enq_7_dec_uops_1_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_prflag <= io_enq_7_dec_uops_1_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_pwflag <= io_enq_7_dec_uops_1_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_pflag_busy <= io_enq_7_dec_uops_1_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_stale_pflag <= io_enq_7_dec_uops_1_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_op1_sel <= io_enq_7_dec_uops_1_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_op2_sel <= io_enq_7_dec_uops_1_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_split_num <= io_enq_7_dec_uops_1_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_self_index <= io_enq_7_dec_uops_1_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_rob_inst_idx <= io_enq_7_dec_uops_1_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_address_num <= io_enq_7_dec_uops_1_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_uopc <= io_enq_7_dec_uops_1_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_inst <= io_enq_7_dec_uops_1_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_debug_inst <= io_enq_7_dec_uops_1_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_is_rvc <= io_enq_7_dec_uops_1_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_debug_pc <= io_enq_7_dec_uops_1_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_iq_type <= io_enq_7_dec_uops_1_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_fu_code <= io_enq_7_dec_uops_1_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_ctrl_br_type <= io_enq_7_dec_uops_1_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_ctrl_op1_sel <= io_enq_7_dec_uops_1_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_ctrl_op2_sel <= io_enq_7_dec_uops_1_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_ctrl_imm_sel <= io_enq_7_dec_uops_1_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_ctrl_op_fcn <= io_enq_7_dec_uops_1_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_ctrl_fcn_dw <= io_enq_7_dec_uops_1_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_ctrl_csr_cmd <= io_enq_7_dec_uops_1_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_ctrl_is_load <= io_enq_7_dec_uops_1_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_ctrl_is_sta <= io_enq_7_dec_uops_1_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_ctrl_is_std <= io_enq_7_dec_uops_1_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_ctrl_op3_sel <= io_enq_7_dec_uops_1_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_iw_state <= io_enq_7_dec_uops_1_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_iw_p1_poisoned <= io_enq_7_dec_uops_1_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_iw_p2_poisoned <= io_enq_7_dec_uops_1_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_is_br <= io_enq_7_dec_uops_1_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_is_jalr <= io_enq_7_dec_uops_1_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_is_jal <= io_enq_7_dec_uops_1_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_is_sfb <= io_enq_7_dec_uops_1_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_br_mask <= io_enq_7_dec_uops_1_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_br_tag <= io_enq_7_dec_uops_1_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_ftq_idx <= io_enq_7_dec_uops_1_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_edge_inst <= io_enq_7_dec_uops_1_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_pc_lob <= io_enq_7_dec_uops_1_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_taken <= io_enq_7_dec_uops_1_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_imm_packed <= io_enq_7_dec_uops_1_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_csr_addr <= io_enq_7_dec_uops_1_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_rob_idx <= io_enq_7_dec_uops_1_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_ldq_idx <= io_enq_7_dec_uops_1_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_stq_idx <= io_enq_7_dec_uops_1_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_rxq_idx <= io_enq_7_dec_uops_1_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_pdst <= io_enq_7_dec_uops_1_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_prs1 <= io_enq_7_dec_uops_1_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_prs2 <= io_enq_7_dec_uops_1_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_prs3 <= io_enq_7_dec_uops_1_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_ppred <= io_enq_7_dec_uops_1_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_prs1_busy <= io_enq_7_dec_uops_1_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_prs2_busy <= io_enq_7_dec_uops_1_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_prs3_busy <= io_enq_7_dec_uops_1_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_ppred_busy <= io_enq_7_dec_uops_1_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_stale_pdst <= io_enq_7_dec_uops_1_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_exception <= io_enq_7_dec_uops_1_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_exc_cause <= io_enq_7_dec_uops_1_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_bypassable <= io_enq_7_dec_uops_1_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_mem_cmd <= io_enq_7_dec_uops_1_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_mem_size <= io_enq_7_dec_uops_1_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_mem_signed <= io_enq_7_dec_uops_1_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_is_fence <= io_enq_7_dec_uops_1_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_is_fencei <= io_enq_7_dec_uops_1_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_is_amo <= io_enq_7_dec_uops_1_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_uses_ldq <= io_enq_7_dec_uops_1_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_uses_stq <= io_enq_7_dec_uops_1_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_is_sys_pc2epc <= io_enq_7_dec_uops_1_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_is_unique <= io_enq_7_dec_uops_1_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_flush_on_commit <= io_enq_7_dec_uops_1_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_ldst_is_rs1 <= io_enq_7_dec_uops_1_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_ldst <= io_enq_7_dec_uops_1_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_lrs1 <= io_enq_7_dec_uops_1_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_lrs2 <= io_enq_7_dec_uops_1_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_lrs3 <= io_enq_7_dec_uops_1_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_ldst_val <= io_enq_7_dec_uops_1_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_dst_rtype <= io_enq_7_dec_uops_1_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_lrs1_rtype <= io_enq_7_dec_uops_1_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_lrs2_rtype <= io_enq_7_dec_uops_1_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_frs3_en <= io_enq_7_dec_uops_1_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_fp_val <= io_enq_7_dec_uops_1_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_fp_single <= io_enq_7_dec_uops_1_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_xcpt_pf_if <= io_enq_7_dec_uops_1_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_xcpt_ae_if <= io_enq_7_dec_uops_1_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_xcpt_ma_if <= io_enq_7_dec_uops_1_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_bp_debug_if <= io_enq_7_dec_uops_1_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_bp_xcpt_if <= io_enq_7_dec_uops_1_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_debug_fsrc <= io_enq_7_dec_uops_1_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_1_debug_tsrc <= io_enq_7_dec_uops_1_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_switch <= io_enq_7_dec_uops_2_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_switch_off <= io_enq_7_dec_uops_2_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_is_unicore <= io_enq_7_dec_uops_2_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_shift <= io_enq_7_dec_uops_2_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_lrs3_rtype <= io_enq_7_dec_uops_2_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_rflag <= io_enq_7_dec_uops_2_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_wflag <= io_enq_7_dec_uops_2_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_prflag <= io_enq_7_dec_uops_2_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_pwflag <= io_enq_7_dec_uops_2_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_pflag_busy <= io_enq_7_dec_uops_2_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_stale_pflag <= io_enq_7_dec_uops_2_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_op1_sel <= io_enq_7_dec_uops_2_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_op2_sel <= io_enq_7_dec_uops_2_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_split_num <= io_enq_7_dec_uops_2_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_self_index <= io_enq_7_dec_uops_2_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_rob_inst_idx <= io_enq_7_dec_uops_2_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_address_num <= io_enq_7_dec_uops_2_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_uopc <= io_enq_7_dec_uops_2_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_inst <= io_enq_7_dec_uops_2_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_debug_inst <= io_enq_7_dec_uops_2_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_is_rvc <= io_enq_7_dec_uops_2_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_debug_pc <= io_enq_7_dec_uops_2_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_iq_type <= io_enq_7_dec_uops_2_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_fu_code <= io_enq_7_dec_uops_2_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_ctrl_br_type <= io_enq_7_dec_uops_2_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_ctrl_op1_sel <= io_enq_7_dec_uops_2_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_ctrl_op2_sel <= io_enq_7_dec_uops_2_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_ctrl_imm_sel <= io_enq_7_dec_uops_2_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_ctrl_op_fcn <= io_enq_7_dec_uops_2_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_ctrl_fcn_dw <= io_enq_7_dec_uops_2_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_ctrl_csr_cmd <= io_enq_7_dec_uops_2_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_ctrl_is_load <= io_enq_7_dec_uops_2_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_ctrl_is_sta <= io_enq_7_dec_uops_2_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_ctrl_is_std <= io_enq_7_dec_uops_2_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_ctrl_op3_sel <= io_enq_7_dec_uops_2_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_iw_state <= io_enq_7_dec_uops_2_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_iw_p1_poisoned <= io_enq_7_dec_uops_2_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_iw_p2_poisoned <= io_enq_7_dec_uops_2_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_is_br <= io_enq_7_dec_uops_2_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_is_jalr <= io_enq_7_dec_uops_2_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_is_jal <= io_enq_7_dec_uops_2_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_is_sfb <= io_enq_7_dec_uops_2_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_br_mask <= io_enq_7_dec_uops_2_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_br_tag <= io_enq_7_dec_uops_2_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_ftq_idx <= io_enq_7_dec_uops_2_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_edge_inst <= io_enq_7_dec_uops_2_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_pc_lob <= io_enq_7_dec_uops_2_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_taken <= io_enq_7_dec_uops_2_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_imm_packed <= io_enq_7_dec_uops_2_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_csr_addr <= io_enq_7_dec_uops_2_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_rob_idx <= io_enq_7_dec_uops_2_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_ldq_idx <= io_enq_7_dec_uops_2_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_stq_idx <= io_enq_7_dec_uops_2_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_rxq_idx <= io_enq_7_dec_uops_2_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_pdst <= io_enq_7_dec_uops_2_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_prs1 <= io_enq_7_dec_uops_2_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_prs2 <= io_enq_7_dec_uops_2_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_prs3 <= io_enq_7_dec_uops_2_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_ppred <= io_enq_7_dec_uops_2_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_prs1_busy <= io_enq_7_dec_uops_2_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_prs2_busy <= io_enq_7_dec_uops_2_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_prs3_busy <= io_enq_7_dec_uops_2_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_ppred_busy <= io_enq_7_dec_uops_2_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_stale_pdst <= io_enq_7_dec_uops_2_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_exception <= io_enq_7_dec_uops_2_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_exc_cause <= io_enq_7_dec_uops_2_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_bypassable <= io_enq_7_dec_uops_2_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_mem_cmd <= io_enq_7_dec_uops_2_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_mem_size <= io_enq_7_dec_uops_2_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_mem_signed <= io_enq_7_dec_uops_2_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_is_fence <= io_enq_7_dec_uops_2_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_is_fencei <= io_enq_7_dec_uops_2_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_is_amo <= io_enq_7_dec_uops_2_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_uses_ldq <= io_enq_7_dec_uops_2_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_uses_stq <= io_enq_7_dec_uops_2_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_is_sys_pc2epc <= io_enq_7_dec_uops_2_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_is_unique <= io_enq_7_dec_uops_2_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_flush_on_commit <= io_enq_7_dec_uops_2_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_ldst_is_rs1 <= io_enq_7_dec_uops_2_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_ldst <= io_enq_7_dec_uops_2_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_lrs1 <= io_enq_7_dec_uops_2_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_lrs2 <= io_enq_7_dec_uops_2_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_lrs3 <= io_enq_7_dec_uops_2_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_ldst_val <= io_enq_7_dec_uops_2_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_dst_rtype <= io_enq_7_dec_uops_2_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_lrs1_rtype <= io_enq_7_dec_uops_2_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_lrs2_rtype <= io_enq_7_dec_uops_2_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_frs3_en <= io_enq_7_dec_uops_2_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_fp_val <= io_enq_7_dec_uops_2_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_fp_single <= io_enq_7_dec_uops_2_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_xcpt_pf_if <= io_enq_7_dec_uops_2_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_xcpt_ae_if <= io_enq_7_dec_uops_2_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_xcpt_ma_if <= io_enq_7_dec_uops_2_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_bp_debug_if <= io_enq_7_dec_uops_2_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_bp_xcpt_if <= io_enq_7_dec_uops_2_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_debug_fsrc <= io_enq_7_dec_uops_2_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_2_debug_tsrc <= io_enq_7_dec_uops_2_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_switch <= io_enq_7_dec_uops_3_switch; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_switch_off <= io_enq_7_dec_uops_3_switch_off; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_is_unicore <= io_enq_7_dec_uops_3_is_unicore; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_shift <= io_enq_7_dec_uops_3_shift; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_lrs3_rtype <= io_enq_7_dec_uops_3_lrs3_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_rflag <= io_enq_7_dec_uops_3_rflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_wflag <= io_enq_7_dec_uops_3_wflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_prflag <= io_enq_7_dec_uops_3_prflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_pwflag <= io_enq_7_dec_uops_3_pwflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_pflag_busy <= io_enq_7_dec_uops_3_pflag_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_stale_pflag <= io_enq_7_dec_uops_3_stale_pflag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_op1_sel <= io_enq_7_dec_uops_3_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_op2_sel <= io_enq_7_dec_uops_3_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_split_num <= io_enq_7_dec_uops_3_split_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_self_index <= io_enq_7_dec_uops_3_self_index; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_rob_inst_idx <= io_enq_7_dec_uops_3_rob_inst_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_address_num <= io_enq_7_dec_uops_3_address_num; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_uopc <= io_enq_7_dec_uops_3_uopc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_inst <= io_enq_7_dec_uops_3_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_debug_inst <= io_enq_7_dec_uops_3_debug_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_is_rvc <= io_enq_7_dec_uops_3_is_rvc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_debug_pc <= io_enq_7_dec_uops_3_debug_pc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_iq_type <= io_enq_7_dec_uops_3_iq_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_fu_code <= io_enq_7_dec_uops_3_fu_code; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_ctrl_br_type <= io_enq_7_dec_uops_3_ctrl_br_type; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_ctrl_op1_sel <= io_enq_7_dec_uops_3_ctrl_op1_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_ctrl_op2_sel <= io_enq_7_dec_uops_3_ctrl_op2_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_ctrl_imm_sel <= io_enq_7_dec_uops_3_ctrl_imm_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_ctrl_op_fcn <= io_enq_7_dec_uops_3_ctrl_op_fcn; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_ctrl_fcn_dw <= io_enq_7_dec_uops_3_ctrl_fcn_dw; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_ctrl_csr_cmd <= io_enq_7_dec_uops_3_ctrl_csr_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_ctrl_is_load <= io_enq_7_dec_uops_3_ctrl_is_load; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_ctrl_is_sta <= io_enq_7_dec_uops_3_ctrl_is_sta; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_ctrl_is_std <= io_enq_7_dec_uops_3_ctrl_is_std; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_ctrl_op3_sel <= io_enq_7_dec_uops_3_ctrl_op3_sel; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_iw_state <= io_enq_7_dec_uops_3_iw_state; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_iw_p1_poisoned <= io_enq_7_dec_uops_3_iw_p1_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_iw_p2_poisoned <= io_enq_7_dec_uops_3_iw_p2_poisoned; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_is_br <= io_enq_7_dec_uops_3_is_br; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_is_jalr <= io_enq_7_dec_uops_3_is_jalr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_is_jal <= io_enq_7_dec_uops_3_is_jal; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_is_sfb <= io_enq_7_dec_uops_3_is_sfb; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_br_mask <= io_enq_7_dec_uops_3_br_mask; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_br_tag <= io_enq_7_dec_uops_3_br_tag; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_ftq_idx <= io_enq_7_dec_uops_3_ftq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_edge_inst <= io_enq_7_dec_uops_3_edge_inst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_pc_lob <= io_enq_7_dec_uops_3_pc_lob; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_taken <= io_enq_7_dec_uops_3_taken; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_imm_packed <= io_enq_7_dec_uops_3_imm_packed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_csr_addr <= io_enq_7_dec_uops_3_csr_addr; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_rob_idx <= io_enq_7_dec_uops_3_rob_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_ldq_idx <= io_enq_7_dec_uops_3_ldq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_stq_idx <= io_enq_7_dec_uops_3_stq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_rxq_idx <= io_enq_7_dec_uops_3_rxq_idx; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_pdst <= io_enq_7_dec_uops_3_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_prs1 <= io_enq_7_dec_uops_3_prs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_prs2 <= io_enq_7_dec_uops_3_prs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_prs3 <= io_enq_7_dec_uops_3_prs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_ppred <= io_enq_7_dec_uops_3_ppred; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_prs1_busy <= io_enq_7_dec_uops_3_prs1_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_prs2_busy <= io_enq_7_dec_uops_3_prs2_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_prs3_busy <= io_enq_7_dec_uops_3_prs3_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_ppred_busy <= io_enq_7_dec_uops_3_ppred_busy; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_stale_pdst <= io_enq_7_dec_uops_3_stale_pdst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_exception <= io_enq_7_dec_uops_3_exception; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_exc_cause <= io_enq_7_dec_uops_3_exc_cause; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_bypassable <= io_enq_7_dec_uops_3_bypassable; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_mem_cmd <= io_enq_7_dec_uops_3_mem_cmd; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_mem_size <= io_enq_7_dec_uops_3_mem_size; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_mem_signed <= io_enq_7_dec_uops_3_mem_signed; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_is_fence <= io_enq_7_dec_uops_3_is_fence; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_is_fencei <= io_enq_7_dec_uops_3_is_fencei; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_is_amo <= io_enq_7_dec_uops_3_is_amo; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_uses_ldq <= io_enq_7_dec_uops_3_uses_ldq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_uses_stq <= io_enq_7_dec_uops_3_uses_stq; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_is_sys_pc2epc <= io_enq_7_dec_uops_3_is_sys_pc2epc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_is_unique <= io_enq_7_dec_uops_3_is_unique; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_flush_on_commit <= io_enq_7_dec_uops_3_flush_on_commit; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_ldst_is_rs1 <= io_enq_7_dec_uops_3_ldst_is_rs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_ldst <= io_enq_7_dec_uops_3_ldst; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_lrs1 <= io_enq_7_dec_uops_3_lrs1; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_lrs2 <= io_enq_7_dec_uops_3_lrs2; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_lrs3 <= io_enq_7_dec_uops_3_lrs3; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_ldst_val <= io_enq_7_dec_uops_3_ldst_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_dst_rtype <= io_enq_7_dec_uops_3_dst_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_lrs1_rtype <= io_enq_7_dec_uops_3_lrs1_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_lrs2_rtype <= io_enq_7_dec_uops_3_lrs2_rtype; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_frs3_en <= io_enq_7_dec_uops_3_frs3_en; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_fp_val <= io_enq_7_dec_uops_3_fp_val; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_fp_single <= io_enq_7_dec_uops_3_fp_single; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_xcpt_pf_if <= io_enq_7_dec_uops_3_xcpt_pf_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_xcpt_ae_if <= io_enq_7_dec_uops_3_xcpt_ae_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_xcpt_ma_if <= io_enq_7_dec_uops_3_xcpt_ma_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_bp_debug_if <= io_enq_7_dec_uops_3_bp_debug_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_bp_xcpt_if <= io_enq_7_dec_uops_3_bp_xcpt_if; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_debug_fsrc <= io_enq_7_dec_uops_3_debug_fsrc; // @[enq_transBuff.scala 119:20]
    end
    if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_dec_uops_3_debug_tsrc <= io_enq_7_dec_uops_3_debug_tsrc; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_7_val_mask_0 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_val_mask_0 <= io_enq_7_val_mask_0; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_7_val_mask_1 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_val_mask_1 <= io_enq_7_val_mask_1; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_7_val_mask_2 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_val_mask_2 <= io_enq_7_val_mask_2; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_buffer_7_val_mask_3 <= 1'h0; // @[enq_transBuff.scala 141:43]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_buffer_7_val_mask_3 <= io_enq_7_val_mask_3; // @[enq_transBuff.scala 119:20]
    end
    if (io_clear) begin // @[enq_transBuff.scala 135:19]
      enq_valid <= 1'h0; // @[enq_transBuff.scala 138:19]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      enq_valid <= io_enq_valid; // @[enq_transBuff.scala 120:19]
    end else if (last_cycle_over) begin // @[enq_transBuff.scala 84:28]
      enq_valid <= 1'h0; // @[enq_transBuff.scala 85:18]
    end
    if (reset) begin // @[enq_transBuff.scala 53:26]
      set_idx <= 5'h0; // @[enq_transBuff.scala 53:26]
    end else if (io_clear) begin // @[enq_transBuff.scala 135:19]
      set_idx <= 5'h0; // @[enq_transBuff.scala 136:17]
    end else if (~io_enq_valid & ~enq_valid) begin // @[enq_transBuff.scala 102:38]
      set_idx <= 5'h0; // @[enq_transBuff.scala 104:17]
    end else if (trans_buffer_io_enq_ready) begin // @[enq_transBuff.scala 106:41]
      set_idx <= _GEN_1;
    end
    if (reset) begin // @[enq_transBuff.scala 54:26]
      set_num <= 5'h0; // @[enq_transBuff.scala 54:26]
    end else if (io_clear) begin // @[enq_transBuff.scala 135:19]
      set_num <= 5'h0; // @[enq_transBuff.scala 137:17]
    end else if (_T_2) begin // @[enq_transBuff.scala 118:71]
      set_num <= io_set_num; // @[enq_transBuff.scala 121:17]
    end else if (~io_enq_valid & ~enq_valid) begin // @[enq_transBuff.scala 102:38]
      set_num <= 5'h0; // @[enq_transBuff.scala 103:17]
    end
    if (_T_2) begin // @[enq_transBuff.scala 78:27]
      REG <= _T_3;
    end else if (enq_valid) begin // @[enq_transBuff.scala 79:28]
      REG <= _T_6 & trans_buffer_io_enq_ready;
    end else begin
      REG <= 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_switch = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_switch_off = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_is_unicore = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_shift = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_lrs3_rtype = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_rflag = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_wflag = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_prflag = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_pwflag = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_pflag_busy = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_stale_pflag = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_op1_sel = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_op2_sel = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_split_num = _RAND_13[5:0];
  _RAND_14 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_self_index = _RAND_14[5:0];
  _RAND_15 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_rob_inst_idx = _RAND_15[5:0];
  _RAND_16 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_address_num = _RAND_16[5:0];
  _RAND_17 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_uopc = _RAND_17[6:0];
  _RAND_18 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_inst = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_debug_inst = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_is_rvc = _RAND_20[0:0];
  _RAND_21 = {2{`RANDOM}};
  enq_buffer_0_dec_uops_0_debug_pc = _RAND_21[39:0];
  _RAND_22 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_iq_type = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_fu_code = _RAND_23[9:0];
  _RAND_24 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_ctrl_br_type = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_ctrl_op1_sel = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_ctrl_op2_sel = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_ctrl_imm_sel = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_ctrl_op_fcn = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_ctrl_fcn_dw = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_ctrl_csr_cmd = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_ctrl_is_load = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_ctrl_is_sta = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_ctrl_is_std = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_ctrl_op3_sel = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_iw_state = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_iw_p1_poisoned = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_iw_p2_poisoned = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_is_br = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_is_jalr = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_is_jal = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_is_sfb = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_br_mask = _RAND_42[11:0];
  _RAND_43 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_br_tag = _RAND_43[3:0];
  _RAND_44 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_ftq_idx = _RAND_44[4:0];
  _RAND_45 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_edge_inst = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_pc_lob = _RAND_46[5:0];
  _RAND_47 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_taken = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_imm_packed = _RAND_48[19:0];
  _RAND_49 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_csr_addr = _RAND_49[11:0];
  _RAND_50 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_rob_idx = _RAND_50[5:0];
  _RAND_51 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_ldq_idx = _RAND_51[4:0];
  _RAND_52 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_stq_idx = _RAND_52[4:0];
  _RAND_53 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_rxq_idx = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_pdst = _RAND_54[6:0];
  _RAND_55 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_prs1 = _RAND_55[6:0];
  _RAND_56 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_prs2 = _RAND_56[6:0];
  _RAND_57 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_prs3 = _RAND_57[6:0];
  _RAND_58 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_ppred = _RAND_58[4:0];
  _RAND_59 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_prs1_busy = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_prs2_busy = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_prs3_busy = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_ppred_busy = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_stale_pdst = _RAND_63[6:0];
  _RAND_64 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_exception = _RAND_64[0:0];
  _RAND_65 = {2{`RANDOM}};
  enq_buffer_0_dec_uops_0_exc_cause = _RAND_65[63:0];
  _RAND_66 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_bypassable = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_mem_cmd = _RAND_67[4:0];
  _RAND_68 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_mem_size = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_mem_signed = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_is_fence = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_is_fencei = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_is_amo = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_uses_ldq = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_uses_stq = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_is_sys_pc2epc = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_is_unique = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_flush_on_commit = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_ldst_is_rs1 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_ldst = _RAND_79[5:0];
  _RAND_80 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_lrs1 = _RAND_80[5:0];
  _RAND_81 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_lrs2 = _RAND_81[5:0];
  _RAND_82 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_lrs3 = _RAND_82[5:0];
  _RAND_83 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_ldst_val = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_dst_rtype = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_lrs1_rtype = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_lrs2_rtype = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_frs3_en = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_fp_val = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_fp_single = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_xcpt_pf_if = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_xcpt_ae_if = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_xcpt_ma_if = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_bp_debug_if = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_bp_xcpt_if = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_debug_fsrc = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_0_debug_tsrc = _RAND_96[1:0];
  _RAND_97 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_switch = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_switch_off = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_is_unicore = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_shift = _RAND_100[2:0];
  _RAND_101 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_lrs3_rtype = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_rflag = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_wflag = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_prflag = _RAND_104[3:0];
  _RAND_105 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_pwflag = _RAND_105[3:0];
  _RAND_106 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_pflag_busy = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_stale_pflag = _RAND_107[3:0];
  _RAND_108 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_op1_sel = _RAND_108[3:0];
  _RAND_109 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_op2_sel = _RAND_109[3:0];
  _RAND_110 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_split_num = _RAND_110[5:0];
  _RAND_111 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_self_index = _RAND_111[5:0];
  _RAND_112 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_rob_inst_idx = _RAND_112[5:0];
  _RAND_113 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_address_num = _RAND_113[5:0];
  _RAND_114 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_uopc = _RAND_114[6:0];
  _RAND_115 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_inst = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_debug_inst = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_is_rvc = _RAND_117[0:0];
  _RAND_118 = {2{`RANDOM}};
  enq_buffer_0_dec_uops_1_debug_pc = _RAND_118[39:0];
  _RAND_119 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_iq_type = _RAND_119[2:0];
  _RAND_120 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_fu_code = _RAND_120[9:0];
  _RAND_121 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_ctrl_br_type = _RAND_121[3:0];
  _RAND_122 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_ctrl_op1_sel = _RAND_122[1:0];
  _RAND_123 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_ctrl_op2_sel = _RAND_123[2:0];
  _RAND_124 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_ctrl_imm_sel = _RAND_124[2:0];
  _RAND_125 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_ctrl_op_fcn = _RAND_125[3:0];
  _RAND_126 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_ctrl_fcn_dw = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_ctrl_csr_cmd = _RAND_127[2:0];
  _RAND_128 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_ctrl_is_load = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_ctrl_is_sta = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_ctrl_is_std = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_ctrl_op3_sel = _RAND_131[1:0];
  _RAND_132 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_iw_state = _RAND_132[1:0];
  _RAND_133 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_iw_p1_poisoned = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_iw_p2_poisoned = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_is_br = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_is_jalr = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_is_jal = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_is_sfb = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_br_mask = _RAND_139[11:0];
  _RAND_140 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_br_tag = _RAND_140[3:0];
  _RAND_141 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_ftq_idx = _RAND_141[4:0];
  _RAND_142 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_edge_inst = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_pc_lob = _RAND_143[5:0];
  _RAND_144 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_taken = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_imm_packed = _RAND_145[19:0];
  _RAND_146 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_csr_addr = _RAND_146[11:0];
  _RAND_147 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_rob_idx = _RAND_147[5:0];
  _RAND_148 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_ldq_idx = _RAND_148[4:0];
  _RAND_149 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_stq_idx = _RAND_149[4:0];
  _RAND_150 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_rxq_idx = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_pdst = _RAND_151[6:0];
  _RAND_152 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_prs1 = _RAND_152[6:0];
  _RAND_153 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_prs2 = _RAND_153[6:0];
  _RAND_154 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_prs3 = _RAND_154[6:0];
  _RAND_155 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_ppred = _RAND_155[4:0];
  _RAND_156 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_prs1_busy = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_prs2_busy = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_prs3_busy = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_ppred_busy = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_stale_pdst = _RAND_160[6:0];
  _RAND_161 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_exception = _RAND_161[0:0];
  _RAND_162 = {2{`RANDOM}};
  enq_buffer_0_dec_uops_1_exc_cause = _RAND_162[63:0];
  _RAND_163 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_bypassable = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_mem_cmd = _RAND_164[4:0];
  _RAND_165 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_mem_size = _RAND_165[1:0];
  _RAND_166 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_mem_signed = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_is_fence = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_is_fencei = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_is_amo = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_uses_ldq = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_uses_stq = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_is_sys_pc2epc = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_is_unique = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_flush_on_commit = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_ldst_is_rs1 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_ldst = _RAND_176[5:0];
  _RAND_177 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_lrs1 = _RAND_177[5:0];
  _RAND_178 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_lrs2 = _RAND_178[5:0];
  _RAND_179 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_lrs3 = _RAND_179[5:0];
  _RAND_180 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_ldst_val = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_dst_rtype = _RAND_181[1:0];
  _RAND_182 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_lrs1_rtype = _RAND_182[1:0];
  _RAND_183 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_lrs2_rtype = _RAND_183[1:0];
  _RAND_184 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_frs3_en = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_fp_val = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_fp_single = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_xcpt_pf_if = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_xcpt_ae_if = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_xcpt_ma_if = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_bp_debug_if = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_bp_xcpt_if = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_debug_fsrc = _RAND_192[1:0];
  _RAND_193 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_1_debug_tsrc = _RAND_193[1:0];
  _RAND_194 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_switch = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_switch_off = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_is_unicore = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_shift = _RAND_197[2:0];
  _RAND_198 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_lrs3_rtype = _RAND_198[1:0];
  _RAND_199 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_rflag = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_wflag = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_prflag = _RAND_201[3:0];
  _RAND_202 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_pwflag = _RAND_202[3:0];
  _RAND_203 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_pflag_busy = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_stale_pflag = _RAND_204[3:0];
  _RAND_205 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_op1_sel = _RAND_205[3:0];
  _RAND_206 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_op2_sel = _RAND_206[3:0];
  _RAND_207 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_split_num = _RAND_207[5:0];
  _RAND_208 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_self_index = _RAND_208[5:0];
  _RAND_209 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_rob_inst_idx = _RAND_209[5:0];
  _RAND_210 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_address_num = _RAND_210[5:0];
  _RAND_211 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_uopc = _RAND_211[6:0];
  _RAND_212 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_inst = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_debug_inst = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_is_rvc = _RAND_214[0:0];
  _RAND_215 = {2{`RANDOM}};
  enq_buffer_0_dec_uops_2_debug_pc = _RAND_215[39:0];
  _RAND_216 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_iq_type = _RAND_216[2:0];
  _RAND_217 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_fu_code = _RAND_217[9:0];
  _RAND_218 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_ctrl_br_type = _RAND_218[3:0];
  _RAND_219 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_ctrl_op1_sel = _RAND_219[1:0];
  _RAND_220 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_ctrl_op2_sel = _RAND_220[2:0];
  _RAND_221 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_ctrl_imm_sel = _RAND_221[2:0];
  _RAND_222 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_ctrl_op_fcn = _RAND_222[3:0];
  _RAND_223 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_ctrl_fcn_dw = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_ctrl_csr_cmd = _RAND_224[2:0];
  _RAND_225 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_ctrl_is_load = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_ctrl_is_sta = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_ctrl_is_std = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_ctrl_op3_sel = _RAND_228[1:0];
  _RAND_229 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_iw_state = _RAND_229[1:0];
  _RAND_230 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_iw_p1_poisoned = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_iw_p2_poisoned = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_is_br = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_is_jalr = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_is_jal = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_is_sfb = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_br_mask = _RAND_236[11:0];
  _RAND_237 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_br_tag = _RAND_237[3:0];
  _RAND_238 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_ftq_idx = _RAND_238[4:0];
  _RAND_239 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_edge_inst = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_pc_lob = _RAND_240[5:0];
  _RAND_241 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_taken = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_imm_packed = _RAND_242[19:0];
  _RAND_243 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_csr_addr = _RAND_243[11:0];
  _RAND_244 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_rob_idx = _RAND_244[5:0];
  _RAND_245 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_ldq_idx = _RAND_245[4:0];
  _RAND_246 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_stq_idx = _RAND_246[4:0];
  _RAND_247 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_rxq_idx = _RAND_247[1:0];
  _RAND_248 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_pdst = _RAND_248[6:0];
  _RAND_249 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_prs1 = _RAND_249[6:0];
  _RAND_250 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_prs2 = _RAND_250[6:0];
  _RAND_251 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_prs3 = _RAND_251[6:0];
  _RAND_252 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_ppred = _RAND_252[4:0];
  _RAND_253 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_prs1_busy = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_prs2_busy = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_prs3_busy = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_ppred_busy = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_stale_pdst = _RAND_257[6:0];
  _RAND_258 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_exception = _RAND_258[0:0];
  _RAND_259 = {2{`RANDOM}};
  enq_buffer_0_dec_uops_2_exc_cause = _RAND_259[63:0];
  _RAND_260 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_bypassable = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_mem_cmd = _RAND_261[4:0];
  _RAND_262 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_mem_size = _RAND_262[1:0];
  _RAND_263 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_mem_signed = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_is_fence = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_is_fencei = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_is_amo = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_uses_ldq = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_uses_stq = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_is_sys_pc2epc = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_is_unique = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_flush_on_commit = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_ldst_is_rs1 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_ldst = _RAND_273[5:0];
  _RAND_274 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_lrs1 = _RAND_274[5:0];
  _RAND_275 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_lrs2 = _RAND_275[5:0];
  _RAND_276 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_lrs3 = _RAND_276[5:0];
  _RAND_277 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_ldst_val = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_dst_rtype = _RAND_278[1:0];
  _RAND_279 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_lrs1_rtype = _RAND_279[1:0];
  _RAND_280 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_lrs2_rtype = _RAND_280[1:0];
  _RAND_281 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_frs3_en = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_fp_val = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_fp_single = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_xcpt_pf_if = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_xcpt_ae_if = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_xcpt_ma_if = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_bp_debug_if = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_bp_xcpt_if = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_debug_fsrc = _RAND_289[1:0];
  _RAND_290 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_2_debug_tsrc = _RAND_290[1:0];
  _RAND_291 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_switch = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_switch_off = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_is_unicore = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_shift = _RAND_294[2:0];
  _RAND_295 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_lrs3_rtype = _RAND_295[1:0];
  _RAND_296 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_rflag = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_wflag = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_prflag = _RAND_298[3:0];
  _RAND_299 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_pwflag = _RAND_299[3:0];
  _RAND_300 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_pflag_busy = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_stale_pflag = _RAND_301[3:0];
  _RAND_302 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_op1_sel = _RAND_302[3:0];
  _RAND_303 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_op2_sel = _RAND_303[3:0];
  _RAND_304 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_split_num = _RAND_304[5:0];
  _RAND_305 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_self_index = _RAND_305[5:0];
  _RAND_306 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_rob_inst_idx = _RAND_306[5:0];
  _RAND_307 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_address_num = _RAND_307[5:0];
  _RAND_308 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_uopc = _RAND_308[6:0];
  _RAND_309 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_inst = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_debug_inst = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_is_rvc = _RAND_311[0:0];
  _RAND_312 = {2{`RANDOM}};
  enq_buffer_0_dec_uops_3_debug_pc = _RAND_312[39:0];
  _RAND_313 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_iq_type = _RAND_313[2:0];
  _RAND_314 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_fu_code = _RAND_314[9:0];
  _RAND_315 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_ctrl_br_type = _RAND_315[3:0];
  _RAND_316 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_ctrl_op1_sel = _RAND_316[1:0];
  _RAND_317 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_ctrl_op2_sel = _RAND_317[2:0];
  _RAND_318 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_ctrl_imm_sel = _RAND_318[2:0];
  _RAND_319 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_ctrl_op_fcn = _RAND_319[3:0];
  _RAND_320 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_ctrl_fcn_dw = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_ctrl_csr_cmd = _RAND_321[2:0];
  _RAND_322 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_ctrl_is_load = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_ctrl_is_sta = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_ctrl_is_std = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_ctrl_op3_sel = _RAND_325[1:0];
  _RAND_326 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_iw_state = _RAND_326[1:0];
  _RAND_327 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_iw_p1_poisoned = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_iw_p2_poisoned = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_is_br = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_is_jalr = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_is_jal = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_is_sfb = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_br_mask = _RAND_333[11:0];
  _RAND_334 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_br_tag = _RAND_334[3:0];
  _RAND_335 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_ftq_idx = _RAND_335[4:0];
  _RAND_336 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_edge_inst = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_pc_lob = _RAND_337[5:0];
  _RAND_338 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_taken = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_imm_packed = _RAND_339[19:0];
  _RAND_340 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_csr_addr = _RAND_340[11:0];
  _RAND_341 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_rob_idx = _RAND_341[5:0];
  _RAND_342 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_ldq_idx = _RAND_342[4:0];
  _RAND_343 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_stq_idx = _RAND_343[4:0];
  _RAND_344 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_rxq_idx = _RAND_344[1:0];
  _RAND_345 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_pdst = _RAND_345[6:0];
  _RAND_346 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_prs1 = _RAND_346[6:0];
  _RAND_347 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_prs2 = _RAND_347[6:0];
  _RAND_348 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_prs3 = _RAND_348[6:0];
  _RAND_349 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_ppred = _RAND_349[4:0];
  _RAND_350 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_prs1_busy = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_prs2_busy = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_prs3_busy = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_ppred_busy = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_stale_pdst = _RAND_354[6:0];
  _RAND_355 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_exception = _RAND_355[0:0];
  _RAND_356 = {2{`RANDOM}};
  enq_buffer_0_dec_uops_3_exc_cause = _RAND_356[63:0];
  _RAND_357 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_bypassable = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_mem_cmd = _RAND_358[4:0];
  _RAND_359 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_mem_size = _RAND_359[1:0];
  _RAND_360 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_mem_signed = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_is_fence = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_is_fencei = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_is_amo = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_uses_ldq = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_uses_stq = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_is_sys_pc2epc = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_is_unique = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_flush_on_commit = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_ldst_is_rs1 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_ldst = _RAND_370[5:0];
  _RAND_371 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_lrs1 = _RAND_371[5:0];
  _RAND_372 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_lrs2 = _RAND_372[5:0];
  _RAND_373 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_lrs3 = _RAND_373[5:0];
  _RAND_374 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_ldst_val = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_dst_rtype = _RAND_375[1:0];
  _RAND_376 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_lrs1_rtype = _RAND_376[1:0];
  _RAND_377 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_lrs2_rtype = _RAND_377[1:0];
  _RAND_378 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_frs3_en = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_fp_val = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_fp_single = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_xcpt_pf_if = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_xcpt_ae_if = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_xcpt_ma_if = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_bp_debug_if = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_bp_xcpt_if = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_debug_fsrc = _RAND_386[1:0];
  _RAND_387 = {1{`RANDOM}};
  enq_buffer_0_dec_uops_3_debug_tsrc = _RAND_387[1:0];
  _RAND_388 = {1{`RANDOM}};
  enq_buffer_0_val_mask_0 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  enq_buffer_0_val_mask_1 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  enq_buffer_0_val_mask_2 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  enq_buffer_0_val_mask_3 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_switch = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_switch_off = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_is_unicore = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_shift = _RAND_395[2:0];
  _RAND_396 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_lrs3_rtype = _RAND_396[1:0];
  _RAND_397 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_rflag = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_wflag = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_prflag = _RAND_399[3:0];
  _RAND_400 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_pwflag = _RAND_400[3:0];
  _RAND_401 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_pflag_busy = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_stale_pflag = _RAND_402[3:0];
  _RAND_403 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_op1_sel = _RAND_403[3:0];
  _RAND_404 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_op2_sel = _RAND_404[3:0];
  _RAND_405 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_split_num = _RAND_405[5:0];
  _RAND_406 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_self_index = _RAND_406[5:0];
  _RAND_407 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_rob_inst_idx = _RAND_407[5:0];
  _RAND_408 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_address_num = _RAND_408[5:0];
  _RAND_409 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_uopc = _RAND_409[6:0];
  _RAND_410 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_inst = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_debug_inst = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_is_rvc = _RAND_412[0:0];
  _RAND_413 = {2{`RANDOM}};
  enq_buffer_1_dec_uops_0_debug_pc = _RAND_413[39:0];
  _RAND_414 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_iq_type = _RAND_414[2:0];
  _RAND_415 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_fu_code = _RAND_415[9:0];
  _RAND_416 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_ctrl_br_type = _RAND_416[3:0];
  _RAND_417 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_ctrl_op1_sel = _RAND_417[1:0];
  _RAND_418 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_ctrl_op2_sel = _RAND_418[2:0];
  _RAND_419 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_ctrl_imm_sel = _RAND_419[2:0];
  _RAND_420 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_ctrl_op_fcn = _RAND_420[3:0];
  _RAND_421 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_ctrl_fcn_dw = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_ctrl_csr_cmd = _RAND_422[2:0];
  _RAND_423 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_ctrl_is_load = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_ctrl_is_sta = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_ctrl_is_std = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_ctrl_op3_sel = _RAND_426[1:0];
  _RAND_427 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_iw_state = _RAND_427[1:0];
  _RAND_428 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_iw_p1_poisoned = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_iw_p2_poisoned = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_is_br = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_is_jalr = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_is_jal = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_is_sfb = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_br_mask = _RAND_434[11:0];
  _RAND_435 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_br_tag = _RAND_435[3:0];
  _RAND_436 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_ftq_idx = _RAND_436[4:0];
  _RAND_437 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_edge_inst = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_pc_lob = _RAND_438[5:0];
  _RAND_439 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_taken = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_imm_packed = _RAND_440[19:0];
  _RAND_441 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_csr_addr = _RAND_441[11:0];
  _RAND_442 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_rob_idx = _RAND_442[5:0];
  _RAND_443 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_ldq_idx = _RAND_443[4:0];
  _RAND_444 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_stq_idx = _RAND_444[4:0];
  _RAND_445 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_rxq_idx = _RAND_445[1:0];
  _RAND_446 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_pdst = _RAND_446[6:0];
  _RAND_447 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_prs1 = _RAND_447[6:0];
  _RAND_448 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_prs2 = _RAND_448[6:0];
  _RAND_449 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_prs3 = _RAND_449[6:0];
  _RAND_450 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_ppred = _RAND_450[4:0];
  _RAND_451 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_prs1_busy = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_prs2_busy = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_prs3_busy = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_ppred_busy = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_stale_pdst = _RAND_455[6:0];
  _RAND_456 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_exception = _RAND_456[0:0];
  _RAND_457 = {2{`RANDOM}};
  enq_buffer_1_dec_uops_0_exc_cause = _RAND_457[63:0];
  _RAND_458 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_bypassable = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_mem_cmd = _RAND_459[4:0];
  _RAND_460 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_mem_size = _RAND_460[1:0];
  _RAND_461 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_mem_signed = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_is_fence = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_is_fencei = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_is_amo = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_uses_ldq = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_uses_stq = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_is_sys_pc2epc = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_is_unique = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_flush_on_commit = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_ldst_is_rs1 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_ldst = _RAND_471[5:0];
  _RAND_472 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_lrs1 = _RAND_472[5:0];
  _RAND_473 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_lrs2 = _RAND_473[5:0];
  _RAND_474 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_lrs3 = _RAND_474[5:0];
  _RAND_475 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_ldst_val = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_dst_rtype = _RAND_476[1:0];
  _RAND_477 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_lrs1_rtype = _RAND_477[1:0];
  _RAND_478 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_lrs2_rtype = _RAND_478[1:0];
  _RAND_479 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_frs3_en = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_fp_val = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_fp_single = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_xcpt_pf_if = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_xcpt_ae_if = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_xcpt_ma_if = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_bp_debug_if = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_bp_xcpt_if = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_debug_fsrc = _RAND_487[1:0];
  _RAND_488 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_0_debug_tsrc = _RAND_488[1:0];
  _RAND_489 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_switch = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_switch_off = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_is_unicore = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_shift = _RAND_492[2:0];
  _RAND_493 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_lrs3_rtype = _RAND_493[1:0];
  _RAND_494 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_rflag = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_wflag = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_prflag = _RAND_496[3:0];
  _RAND_497 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_pwflag = _RAND_497[3:0];
  _RAND_498 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_pflag_busy = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_stale_pflag = _RAND_499[3:0];
  _RAND_500 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_op1_sel = _RAND_500[3:0];
  _RAND_501 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_op2_sel = _RAND_501[3:0];
  _RAND_502 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_split_num = _RAND_502[5:0];
  _RAND_503 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_self_index = _RAND_503[5:0];
  _RAND_504 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_rob_inst_idx = _RAND_504[5:0];
  _RAND_505 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_address_num = _RAND_505[5:0];
  _RAND_506 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_uopc = _RAND_506[6:0];
  _RAND_507 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_inst = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_debug_inst = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_is_rvc = _RAND_509[0:0];
  _RAND_510 = {2{`RANDOM}};
  enq_buffer_1_dec_uops_1_debug_pc = _RAND_510[39:0];
  _RAND_511 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_iq_type = _RAND_511[2:0];
  _RAND_512 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_fu_code = _RAND_512[9:0];
  _RAND_513 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_ctrl_br_type = _RAND_513[3:0];
  _RAND_514 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_ctrl_op1_sel = _RAND_514[1:0];
  _RAND_515 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_ctrl_op2_sel = _RAND_515[2:0];
  _RAND_516 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_ctrl_imm_sel = _RAND_516[2:0];
  _RAND_517 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_ctrl_op_fcn = _RAND_517[3:0];
  _RAND_518 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_ctrl_fcn_dw = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_ctrl_csr_cmd = _RAND_519[2:0];
  _RAND_520 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_ctrl_is_load = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_ctrl_is_sta = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_ctrl_is_std = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_ctrl_op3_sel = _RAND_523[1:0];
  _RAND_524 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_iw_state = _RAND_524[1:0];
  _RAND_525 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_iw_p1_poisoned = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_iw_p2_poisoned = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_is_br = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_is_jalr = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_is_jal = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_is_sfb = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_br_mask = _RAND_531[11:0];
  _RAND_532 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_br_tag = _RAND_532[3:0];
  _RAND_533 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_ftq_idx = _RAND_533[4:0];
  _RAND_534 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_edge_inst = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_pc_lob = _RAND_535[5:0];
  _RAND_536 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_taken = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_imm_packed = _RAND_537[19:0];
  _RAND_538 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_csr_addr = _RAND_538[11:0];
  _RAND_539 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_rob_idx = _RAND_539[5:0];
  _RAND_540 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_ldq_idx = _RAND_540[4:0];
  _RAND_541 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_stq_idx = _RAND_541[4:0];
  _RAND_542 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_rxq_idx = _RAND_542[1:0];
  _RAND_543 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_pdst = _RAND_543[6:0];
  _RAND_544 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_prs1 = _RAND_544[6:0];
  _RAND_545 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_prs2 = _RAND_545[6:0];
  _RAND_546 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_prs3 = _RAND_546[6:0];
  _RAND_547 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_ppred = _RAND_547[4:0];
  _RAND_548 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_prs1_busy = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_prs2_busy = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_prs3_busy = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_ppred_busy = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_stale_pdst = _RAND_552[6:0];
  _RAND_553 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_exception = _RAND_553[0:0];
  _RAND_554 = {2{`RANDOM}};
  enq_buffer_1_dec_uops_1_exc_cause = _RAND_554[63:0];
  _RAND_555 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_bypassable = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_mem_cmd = _RAND_556[4:0];
  _RAND_557 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_mem_size = _RAND_557[1:0];
  _RAND_558 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_mem_signed = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_is_fence = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_is_fencei = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_is_amo = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_uses_ldq = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_uses_stq = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_is_sys_pc2epc = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_is_unique = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_flush_on_commit = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_ldst_is_rs1 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_ldst = _RAND_568[5:0];
  _RAND_569 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_lrs1 = _RAND_569[5:0];
  _RAND_570 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_lrs2 = _RAND_570[5:0];
  _RAND_571 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_lrs3 = _RAND_571[5:0];
  _RAND_572 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_ldst_val = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_dst_rtype = _RAND_573[1:0];
  _RAND_574 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_lrs1_rtype = _RAND_574[1:0];
  _RAND_575 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_lrs2_rtype = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_frs3_en = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_fp_val = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_fp_single = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_xcpt_pf_if = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_xcpt_ae_if = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_xcpt_ma_if = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_bp_debug_if = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_bp_xcpt_if = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_debug_fsrc = _RAND_584[1:0];
  _RAND_585 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_1_debug_tsrc = _RAND_585[1:0];
  _RAND_586 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_switch = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_switch_off = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_is_unicore = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_shift = _RAND_589[2:0];
  _RAND_590 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_lrs3_rtype = _RAND_590[1:0];
  _RAND_591 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_rflag = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_wflag = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_prflag = _RAND_593[3:0];
  _RAND_594 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_pwflag = _RAND_594[3:0];
  _RAND_595 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_pflag_busy = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_stale_pflag = _RAND_596[3:0];
  _RAND_597 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_op1_sel = _RAND_597[3:0];
  _RAND_598 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_op2_sel = _RAND_598[3:0];
  _RAND_599 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_split_num = _RAND_599[5:0];
  _RAND_600 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_self_index = _RAND_600[5:0];
  _RAND_601 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_rob_inst_idx = _RAND_601[5:0];
  _RAND_602 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_address_num = _RAND_602[5:0];
  _RAND_603 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_uopc = _RAND_603[6:0];
  _RAND_604 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_inst = _RAND_604[31:0];
  _RAND_605 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_debug_inst = _RAND_605[31:0];
  _RAND_606 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_is_rvc = _RAND_606[0:0];
  _RAND_607 = {2{`RANDOM}};
  enq_buffer_1_dec_uops_2_debug_pc = _RAND_607[39:0];
  _RAND_608 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_iq_type = _RAND_608[2:0];
  _RAND_609 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_fu_code = _RAND_609[9:0];
  _RAND_610 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_ctrl_br_type = _RAND_610[3:0];
  _RAND_611 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_ctrl_op1_sel = _RAND_611[1:0];
  _RAND_612 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_ctrl_op2_sel = _RAND_612[2:0];
  _RAND_613 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_ctrl_imm_sel = _RAND_613[2:0];
  _RAND_614 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_ctrl_op_fcn = _RAND_614[3:0];
  _RAND_615 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_ctrl_fcn_dw = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_ctrl_csr_cmd = _RAND_616[2:0];
  _RAND_617 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_ctrl_is_load = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_ctrl_is_sta = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_ctrl_is_std = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_ctrl_op3_sel = _RAND_620[1:0];
  _RAND_621 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_iw_state = _RAND_621[1:0];
  _RAND_622 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_iw_p1_poisoned = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_iw_p2_poisoned = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_is_br = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_is_jalr = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_is_jal = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_is_sfb = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_br_mask = _RAND_628[11:0];
  _RAND_629 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_br_tag = _RAND_629[3:0];
  _RAND_630 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_ftq_idx = _RAND_630[4:0];
  _RAND_631 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_edge_inst = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_pc_lob = _RAND_632[5:0];
  _RAND_633 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_taken = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_imm_packed = _RAND_634[19:0];
  _RAND_635 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_csr_addr = _RAND_635[11:0];
  _RAND_636 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_rob_idx = _RAND_636[5:0];
  _RAND_637 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_ldq_idx = _RAND_637[4:0];
  _RAND_638 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_stq_idx = _RAND_638[4:0];
  _RAND_639 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_rxq_idx = _RAND_639[1:0];
  _RAND_640 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_pdst = _RAND_640[6:0];
  _RAND_641 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_prs1 = _RAND_641[6:0];
  _RAND_642 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_prs2 = _RAND_642[6:0];
  _RAND_643 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_prs3 = _RAND_643[6:0];
  _RAND_644 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_ppred = _RAND_644[4:0];
  _RAND_645 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_prs1_busy = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_prs2_busy = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_prs3_busy = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_ppred_busy = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_stale_pdst = _RAND_649[6:0];
  _RAND_650 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_exception = _RAND_650[0:0];
  _RAND_651 = {2{`RANDOM}};
  enq_buffer_1_dec_uops_2_exc_cause = _RAND_651[63:0];
  _RAND_652 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_bypassable = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_mem_cmd = _RAND_653[4:0];
  _RAND_654 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_mem_size = _RAND_654[1:0];
  _RAND_655 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_mem_signed = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_is_fence = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_is_fencei = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_is_amo = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_uses_ldq = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_uses_stq = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_is_sys_pc2epc = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_is_unique = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_flush_on_commit = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_ldst_is_rs1 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_ldst = _RAND_665[5:0];
  _RAND_666 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_lrs1 = _RAND_666[5:0];
  _RAND_667 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_lrs2 = _RAND_667[5:0];
  _RAND_668 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_lrs3 = _RAND_668[5:0];
  _RAND_669 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_ldst_val = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_dst_rtype = _RAND_670[1:0];
  _RAND_671 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_lrs1_rtype = _RAND_671[1:0];
  _RAND_672 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_lrs2_rtype = _RAND_672[1:0];
  _RAND_673 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_frs3_en = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_fp_val = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_fp_single = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_xcpt_pf_if = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_xcpt_ae_if = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_xcpt_ma_if = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_bp_debug_if = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_bp_xcpt_if = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_debug_fsrc = _RAND_681[1:0];
  _RAND_682 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_2_debug_tsrc = _RAND_682[1:0];
  _RAND_683 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_switch = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_switch_off = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_is_unicore = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_shift = _RAND_686[2:0];
  _RAND_687 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_lrs3_rtype = _RAND_687[1:0];
  _RAND_688 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_rflag = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_wflag = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_prflag = _RAND_690[3:0];
  _RAND_691 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_pwflag = _RAND_691[3:0];
  _RAND_692 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_pflag_busy = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_stale_pflag = _RAND_693[3:0];
  _RAND_694 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_op1_sel = _RAND_694[3:0];
  _RAND_695 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_op2_sel = _RAND_695[3:0];
  _RAND_696 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_split_num = _RAND_696[5:0];
  _RAND_697 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_self_index = _RAND_697[5:0];
  _RAND_698 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_rob_inst_idx = _RAND_698[5:0];
  _RAND_699 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_address_num = _RAND_699[5:0];
  _RAND_700 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_uopc = _RAND_700[6:0];
  _RAND_701 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_inst = _RAND_701[31:0];
  _RAND_702 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_debug_inst = _RAND_702[31:0];
  _RAND_703 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_is_rvc = _RAND_703[0:0];
  _RAND_704 = {2{`RANDOM}};
  enq_buffer_1_dec_uops_3_debug_pc = _RAND_704[39:0];
  _RAND_705 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_iq_type = _RAND_705[2:0];
  _RAND_706 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_fu_code = _RAND_706[9:0];
  _RAND_707 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_ctrl_br_type = _RAND_707[3:0];
  _RAND_708 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_ctrl_op1_sel = _RAND_708[1:0];
  _RAND_709 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_ctrl_op2_sel = _RAND_709[2:0];
  _RAND_710 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_ctrl_imm_sel = _RAND_710[2:0];
  _RAND_711 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_ctrl_op_fcn = _RAND_711[3:0];
  _RAND_712 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_ctrl_fcn_dw = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_ctrl_csr_cmd = _RAND_713[2:0];
  _RAND_714 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_ctrl_is_load = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_ctrl_is_sta = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_ctrl_is_std = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_ctrl_op3_sel = _RAND_717[1:0];
  _RAND_718 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_iw_state = _RAND_718[1:0];
  _RAND_719 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_iw_p1_poisoned = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_iw_p2_poisoned = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_is_br = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_is_jalr = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_is_jal = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_is_sfb = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_br_mask = _RAND_725[11:0];
  _RAND_726 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_br_tag = _RAND_726[3:0];
  _RAND_727 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_ftq_idx = _RAND_727[4:0];
  _RAND_728 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_edge_inst = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_pc_lob = _RAND_729[5:0];
  _RAND_730 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_taken = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_imm_packed = _RAND_731[19:0];
  _RAND_732 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_csr_addr = _RAND_732[11:0];
  _RAND_733 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_rob_idx = _RAND_733[5:0];
  _RAND_734 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_ldq_idx = _RAND_734[4:0];
  _RAND_735 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_stq_idx = _RAND_735[4:0];
  _RAND_736 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_rxq_idx = _RAND_736[1:0];
  _RAND_737 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_pdst = _RAND_737[6:0];
  _RAND_738 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_prs1 = _RAND_738[6:0];
  _RAND_739 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_prs2 = _RAND_739[6:0];
  _RAND_740 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_prs3 = _RAND_740[6:0];
  _RAND_741 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_ppred = _RAND_741[4:0];
  _RAND_742 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_prs1_busy = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_prs2_busy = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_prs3_busy = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_ppred_busy = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_stale_pdst = _RAND_746[6:0];
  _RAND_747 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_exception = _RAND_747[0:0];
  _RAND_748 = {2{`RANDOM}};
  enq_buffer_1_dec_uops_3_exc_cause = _RAND_748[63:0];
  _RAND_749 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_bypassable = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_mem_cmd = _RAND_750[4:0];
  _RAND_751 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_mem_size = _RAND_751[1:0];
  _RAND_752 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_mem_signed = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_is_fence = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_is_fencei = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_is_amo = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_uses_ldq = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_uses_stq = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_is_sys_pc2epc = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_is_unique = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_flush_on_commit = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_ldst_is_rs1 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_ldst = _RAND_762[5:0];
  _RAND_763 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_lrs1 = _RAND_763[5:0];
  _RAND_764 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_lrs2 = _RAND_764[5:0];
  _RAND_765 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_lrs3 = _RAND_765[5:0];
  _RAND_766 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_ldst_val = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_dst_rtype = _RAND_767[1:0];
  _RAND_768 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_lrs1_rtype = _RAND_768[1:0];
  _RAND_769 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_lrs2_rtype = _RAND_769[1:0];
  _RAND_770 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_frs3_en = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_fp_val = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_fp_single = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_xcpt_pf_if = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_xcpt_ae_if = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_xcpt_ma_if = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_bp_debug_if = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_bp_xcpt_if = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_debug_fsrc = _RAND_778[1:0];
  _RAND_779 = {1{`RANDOM}};
  enq_buffer_1_dec_uops_3_debug_tsrc = _RAND_779[1:0];
  _RAND_780 = {1{`RANDOM}};
  enq_buffer_1_val_mask_0 = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  enq_buffer_1_val_mask_1 = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  enq_buffer_1_val_mask_2 = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  enq_buffer_1_val_mask_3 = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_switch = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_switch_off = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_is_unicore = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_shift = _RAND_787[2:0];
  _RAND_788 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_lrs3_rtype = _RAND_788[1:0];
  _RAND_789 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_rflag = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_wflag = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_prflag = _RAND_791[3:0];
  _RAND_792 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_pwflag = _RAND_792[3:0];
  _RAND_793 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_pflag_busy = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_stale_pflag = _RAND_794[3:0];
  _RAND_795 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_op1_sel = _RAND_795[3:0];
  _RAND_796 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_op2_sel = _RAND_796[3:0];
  _RAND_797 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_split_num = _RAND_797[5:0];
  _RAND_798 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_self_index = _RAND_798[5:0];
  _RAND_799 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_rob_inst_idx = _RAND_799[5:0];
  _RAND_800 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_address_num = _RAND_800[5:0];
  _RAND_801 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_uopc = _RAND_801[6:0];
  _RAND_802 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_inst = _RAND_802[31:0];
  _RAND_803 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_debug_inst = _RAND_803[31:0];
  _RAND_804 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_is_rvc = _RAND_804[0:0];
  _RAND_805 = {2{`RANDOM}};
  enq_buffer_2_dec_uops_0_debug_pc = _RAND_805[39:0];
  _RAND_806 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_iq_type = _RAND_806[2:0];
  _RAND_807 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_fu_code = _RAND_807[9:0];
  _RAND_808 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_ctrl_br_type = _RAND_808[3:0];
  _RAND_809 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_ctrl_op1_sel = _RAND_809[1:0];
  _RAND_810 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_ctrl_op2_sel = _RAND_810[2:0];
  _RAND_811 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_ctrl_imm_sel = _RAND_811[2:0];
  _RAND_812 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_ctrl_op_fcn = _RAND_812[3:0];
  _RAND_813 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_ctrl_fcn_dw = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_ctrl_csr_cmd = _RAND_814[2:0];
  _RAND_815 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_ctrl_is_load = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_ctrl_is_sta = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_ctrl_is_std = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_ctrl_op3_sel = _RAND_818[1:0];
  _RAND_819 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_iw_state = _RAND_819[1:0];
  _RAND_820 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_iw_p1_poisoned = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_iw_p2_poisoned = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_is_br = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_is_jalr = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_is_jal = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_is_sfb = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_br_mask = _RAND_826[11:0];
  _RAND_827 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_br_tag = _RAND_827[3:0];
  _RAND_828 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_ftq_idx = _RAND_828[4:0];
  _RAND_829 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_edge_inst = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_pc_lob = _RAND_830[5:0];
  _RAND_831 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_taken = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_imm_packed = _RAND_832[19:0];
  _RAND_833 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_csr_addr = _RAND_833[11:0];
  _RAND_834 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_rob_idx = _RAND_834[5:0];
  _RAND_835 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_ldq_idx = _RAND_835[4:0];
  _RAND_836 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_stq_idx = _RAND_836[4:0];
  _RAND_837 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_rxq_idx = _RAND_837[1:0];
  _RAND_838 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_pdst = _RAND_838[6:0];
  _RAND_839 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_prs1 = _RAND_839[6:0];
  _RAND_840 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_prs2 = _RAND_840[6:0];
  _RAND_841 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_prs3 = _RAND_841[6:0];
  _RAND_842 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_ppred = _RAND_842[4:0];
  _RAND_843 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_prs1_busy = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_prs2_busy = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_prs3_busy = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_ppred_busy = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_stale_pdst = _RAND_847[6:0];
  _RAND_848 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_exception = _RAND_848[0:0];
  _RAND_849 = {2{`RANDOM}};
  enq_buffer_2_dec_uops_0_exc_cause = _RAND_849[63:0];
  _RAND_850 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_bypassable = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_mem_cmd = _RAND_851[4:0];
  _RAND_852 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_mem_size = _RAND_852[1:0];
  _RAND_853 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_mem_signed = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_is_fence = _RAND_854[0:0];
  _RAND_855 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_is_fencei = _RAND_855[0:0];
  _RAND_856 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_is_amo = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_uses_ldq = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_uses_stq = _RAND_858[0:0];
  _RAND_859 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_is_sys_pc2epc = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_is_unique = _RAND_860[0:0];
  _RAND_861 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_flush_on_commit = _RAND_861[0:0];
  _RAND_862 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_ldst_is_rs1 = _RAND_862[0:0];
  _RAND_863 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_ldst = _RAND_863[5:0];
  _RAND_864 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_lrs1 = _RAND_864[5:0];
  _RAND_865 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_lrs2 = _RAND_865[5:0];
  _RAND_866 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_lrs3 = _RAND_866[5:0];
  _RAND_867 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_ldst_val = _RAND_867[0:0];
  _RAND_868 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_dst_rtype = _RAND_868[1:0];
  _RAND_869 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_lrs1_rtype = _RAND_869[1:0];
  _RAND_870 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_lrs2_rtype = _RAND_870[1:0];
  _RAND_871 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_frs3_en = _RAND_871[0:0];
  _RAND_872 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_fp_val = _RAND_872[0:0];
  _RAND_873 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_fp_single = _RAND_873[0:0];
  _RAND_874 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_xcpt_pf_if = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_xcpt_ae_if = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_xcpt_ma_if = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_bp_debug_if = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_bp_xcpt_if = _RAND_878[0:0];
  _RAND_879 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_debug_fsrc = _RAND_879[1:0];
  _RAND_880 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_0_debug_tsrc = _RAND_880[1:0];
  _RAND_881 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_switch = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_switch_off = _RAND_882[0:0];
  _RAND_883 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_is_unicore = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_shift = _RAND_884[2:0];
  _RAND_885 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_lrs3_rtype = _RAND_885[1:0];
  _RAND_886 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_rflag = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_wflag = _RAND_887[0:0];
  _RAND_888 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_prflag = _RAND_888[3:0];
  _RAND_889 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_pwflag = _RAND_889[3:0];
  _RAND_890 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_pflag_busy = _RAND_890[0:0];
  _RAND_891 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_stale_pflag = _RAND_891[3:0];
  _RAND_892 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_op1_sel = _RAND_892[3:0];
  _RAND_893 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_op2_sel = _RAND_893[3:0];
  _RAND_894 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_split_num = _RAND_894[5:0];
  _RAND_895 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_self_index = _RAND_895[5:0];
  _RAND_896 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_rob_inst_idx = _RAND_896[5:0];
  _RAND_897 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_address_num = _RAND_897[5:0];
  _RAND_898 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_uopc = _RAND_898[6:0];
  _RAND_899 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_inst = _RAND_899[31:0];
  _RAND_900 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_debug_inst = _RAND_900[31:0];
  _RAND_901 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_is_rvc = _RAND_901[0:0];
  _RAND_902 = {2{`RANDOM}};
  enq_buffer_2_dec_uops_1_debug_pc = _RAND_902[39:0];
  _RAND_903 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_iq_type = _RAND_903[2:0];
  _RAND_904 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_fu_code = _RAND_904[9:0];
  _RAND_905 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_ctrl_br_type = _RAND_905[3:0];
  _RAND_906 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_ctrl_op1_sel = _RAND_906[1:0];
  _RAND_907 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_ctrl_op2_sel = _RAND_907[2:0];
  _RAND_908 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_ctrl_imm_sel = _RAND_908[2:0];
  _RAND_909 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_ctrl_op_fcn = _RAND_909[3:0];
  _RAND_910 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_ctrl_fcn_dw = _RAND_910[0:0];
  _RAND_911 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_ctrl_csr_cmd = _RAND_911[2:0];
  _RAND_912 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_ctrl_is_load = _RAND_912[0:0];
  _RAND_913 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_ctrl_is_sta = _RAND_913[0:0];
  _RAND_914 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_ctrl_is_std = _RAND_914[0:0];
  _RAND_915 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_ctrl_op3_sel = _RAND_915[1:0];
  _RAND_916 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_iw_state = _RAND_916[1:0];
  _RAND_917 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_iw_p1_poisoned = _RAND_917[0:0];
  _RAND_918 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_iw_p2_poisoned = _RAND_918[0:0];
  _RAND_919 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_is_br = _RAND_919[0:0];
  _RAND_920 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_is_jalr = _RAND_920[0:0];
  _RAND_921 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_is_jal = _RAND_921[0:0];
  _RAND_922 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_is_sfb = _RAND_922[0:0];
  _RAND_923 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_br_mask = _RAND_923[11:0];
  _RAND_924 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_br_tag = _RAND_924[3:0];
  _RAND_925 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_ftq_idx = _RAND_925[4:0];
  _RAND_926 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_edge_inst = _RAND_926[0:0];
  _RAND_927 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_pc_lob = _RAND_927[5:0];
  _RAND_928 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_taken = _RAND_928[0:0];
  _RAND_929 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_imm_packed = _RAND_929[19:0];
  _RAND_930 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_csr_addr = _RAND_930[11:0];
  _RAND_931 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_rob_idx = _RAND_931[5:0];
  _RAND_932 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_ldq_idx = _RAND_932[4:0];
  _RAND_933 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_stq_idx = _RAND_933[4:0];
  _RAND_934 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_rxq_idx = _RAND_934[1:0];
  _RAND_935 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_pdst = _RAND_935[6:0];
  _RAND_936 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_prs1 = _RAND_936[6:0];
  _RAND_937 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_prs2 = _RAND_937[6:0];
  _RAND_938 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_prs3 = _RAND_938[6:0];
  _RAND_939 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_ppred = _RAND_939[4:0];
  _RAND_940 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_prs1_busy = _RAND_940[0:0];
  _RAND_941 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_prs2_busy = _RAND_941[0:0];
  _RAND_942 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_prs3_busy = _RAND_942[0:0];
  _RAND_943 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_ppred_busy = _RAND_943[0:0];
  _RAND_944 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_stale_pdst = _RAND_944[6:0];
  _RAND_945 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_exception = _RAND_945[0:0];
  _RAND_946 = {2{`RANDOM}};
  enq_buffer_2_dec_uops_1_exc_cause = _RAND_946[63:0];
  _RAND_947 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_bypassable = _RAND_947[0:0];
  _RAND_948 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_mem_cmd = _RAND_948[4:0];
  _RAND_949 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_mem_size = _RAND_949[1:0];
  _RAND_950 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_mem_signed = _RAND_950[0:0];
  _RAND_951 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_is_fence = _RAND_951[0:0];
  _RAND_952 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_is_fencei = _RAND_952[0:0];
  _RAND_953 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_is_amo = _RAND_953[0:0];
  _RAND_954 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_uses_ldq = _RAND_954[0:0];
  _RAND_955 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_uses_stq = _RAND_955[0:0];
  _RAND_956 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_is_sys_pc2epc = _RAND_956[0:0];
  _RAND_957 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_is_unique = _RAND_957[0:0];
  _RAND_958 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_flush_on_commit = _RAND_958[0:0];
  _RAND_959 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_ldst_is_rs1 = _RAND_959[0:0];
  _RAND_960 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_ldst = _RAND_960[5:0];
  _RAND_961 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_lrs1 = _RAND_961[5:0];
  _RAND_962 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_lrs2 = _RAND_962[5:0];
  _RAND_963 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_lrs3 = _RAND_963[5:0];
  _RAND_964 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_ldst_val = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_dst_rtype = _RAND_965[1:0];
  _RAND_966 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_lrs1_rtype = _RAND_966[1:0];
  _RAND_967 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_lrs2_rtype = _RAND_967[1:0];
  _RAND_968 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_frs3_en = _RAND_968[0:0];
  _RAND_969 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_fp_val = _RAND_969[0:0];
  _RAND_970 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_fp_single = _RAND_970[0:0];
  _RAND_971 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_xcpt_pf_if = _RAND_971[0:0];
  _RAND_972 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_xcpt_ae_if = _RAND_972[0:0];
  _RAND_973 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_xcpt_ma_if = _RAND_973[0:0];
  _RAND_974 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_bp_debug_if = _RAND_974[0:0];
  _RAND_975 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_bp_xcpt_if = _RAND_975[0:0];
  _RAND_976 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_debug_fsrc = _RAND_976[1:0];
  _RAND_977 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_1_debug_tsrc = _RAND_977[1:0];
  _RAND_978 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_switch = _RAND_978[0:0];
  _RAND_979 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_switch_off = _RAND_979[0:0];
  _RAND_980 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_is_unicore = _RAND_980[0:0];
  _RAND_981 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_shift = _RAND_981[2:0];
  _RAND_982 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_lrs3_rtype = _RAND_982[1:0];
  _RAND_983 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_rflag = _RAND_983[0:0];
  _RAND_984 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_wflag = _RAND_984[0:0];
  _RAND_985 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_prflag = _RAND_985[3:0];
  _RAND_986 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_pwflag = _RAND_986[3:0];
  _RAND_987 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_pflag_busy = _RAND_987[0:0];
  _RAND_988 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_stale_pflag = _RAND_988[3:0];
  _RAND_989 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_op1_sel = _RAND_989[3:0];
  _RAND_990 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_op2_sel = _RAND_990[3:0];
  _RAND_991 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_split_num = _RAND_991[5:0];
  _RAND_992 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_self_index = _RAND_992[5:0];
  _RAND_993 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_rob_inst_idx = _RAND_993[5:0];
  _RAND_994 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_address_num = _RAND_994[5:0];
  _RAND_995 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_uopc = _RAND_995[6:0];
  _RAND_996 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_inst = _RAND_996[31:0];
  _RAND_997 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_debug_inst = _RAND_997[31:0];
  _RAND_998 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_is_rvc = _RAND_998[0:0];
  _RAND_999 = {2{`RANDOM}};
  enq_buffer_2_dec_uops_2_debug_pc = _RAND_999[39:0];
  _RAND_1000 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_iq_type = _RAND_1000[2:0];
  _RAND_1001 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_fu_code = _RAND_1001[9:0];
  _RAND_1002 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_ctrl_br_type = _RAND_1002[3:0];
  _RAND_1003 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_ctrl_op1_sel = _RAND_1003[1:0];
  _RAND_1004 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_ctrl_op2_sel = _RAND_1004[2:0];
  _RAND_1005 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_ctrl_imm_sel = _RAND_1005[2:0];
  _RAND_1006 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_ctrl_op_fcn = _RAND_1006[3:0];
  _RAND_1007 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_ctrl_fcn_dw = _RAND_1007[0:0];
  _RAND_1008 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_ctrl_csr_cmd = _RAND_1008[2:0];
  _RAND_1009 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_ctrl_is_load = _RAND_1009[0:0];
  _RAND_1010 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_ctrl_is_sta = _RAND_1010[0:0];
  _RAND_1011 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_ctrl_is_std = _RAND_1011[0:0];
  _RAND_1012 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_ctrl_op3_sel = _RAND_1012[1:0];
  _RAND_1013 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_iw_state = _RAND_1013[1:0];
  _RAND_1014 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_iw_p1_poisoned = _RAND_1014[0:0];
  _RAND_1015 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_iw_p2_poisoned = _RAND_1015[0:0];
  _RAND_1016 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_is_br = _RAND_1016[0:0];
  _RAND_1017 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_is_jalr = _RAND_1017[0:0];
  _RAND_1018 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_is_jal = _RAND_1018[0:0];
  _RAND_1019 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_is_sfb = _RAND_1019[0:0];
  _RAND_1020 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_br_mask = _RAND_1020[11:0];
  _RAND_1021 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_br_tag = _RAND_1021[3:0];
  _RAND_1022 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_ftq_idx = _RAND_1022[4:0];
  _RAND_1023 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_edge_inst = _RAND_1023[0:0];
  _RAND_1024 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_pc_lob = _RAND_1024[5:0];
  _RAND_1025 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_taken = _RAND_1025[0:0];
  _RAND_1026 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_imm_packed = _RAND_1026[19:0];
  _RAND_1027 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_csr_addr = _RAND_1027[11:0];
  _RAND_1028 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_rob_idx = _RAND_1028[5:0];
  _RAND_1029 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_ldq_idx = _RAND_1029[4:0];
  _RAND_1030 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_stq_idx = _RAND_1030[4:0];
  _RAND_1031 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_rxq_idx = _RAND_1031[1:0];
  _RAND_1032 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_pdst = _RAND_1032[6:0];
  _RAND_1033 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_prs1 = _RAND_1033[6:0];
  _RAND_1034 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_prs2 = _RAND_1034[6:0];
  _RAND_1035 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_prs3 = _RAND_1035[6:0];
  _RAND_1036 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_ppred = _RAND_1036[4:0];
  _RAND_1037 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_prs1_busy = _RAND_1037[0:0];
  _RAND_1038 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_prs2_busy = _RAND_1038[0:0];
  _RAND_1039 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_prs3_busy = _RAND_1039[0:0];
  _RAND_1040 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_ppred_busy = _RAND_1040[0:0];
  _RAND_1041 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_stale_pdst = _RAND_1041[6:0];
  _RAND_1042 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_exception = _RAND_1042[0:0];
  _RAND_1043 = {2{`RANDOM}};
  enq_buffer_2_dec_uops_2_exc_cause = _RAND_1043[63:0];
  _RAND_1044 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_bypassable = _RAND_1044[0:0];
  _RAND_1045 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_mem_cmd = _RAND_1045[4:0];
  _RAND_1046 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_mem_size = _RAND_1046[1:0];
  _RAND_1047 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_mem_signed = _RAND_1047[0:0];
  _RAND_1048 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_is_fence = _RAND_1048[0:0];
  _RAND_1049 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_is_fencei = _RAND_1049[0:0];
  _RAND_1050 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_is_amo = _RAND_1050[0:0];
  _RAND_1051 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_uses_ldq = _RAND_1051[0:0];
  _RAND_1052 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_uses_stq = _RAND_1052[0:0];
  _RAND_1053 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_is_sys_pc2epc = _RAND_1053[0:0];
  _RAND_1054 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_is_unique = _RAND_1054[0:0];
  _RAND_1055 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_flush_on_commit = _RAND_1055[0:0];
  _RAND_1056 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_ldst_is_rs1 = _RAND_1056[0:0];
  _RAND_1057 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_ldst = _RAND_1057[5:0];
  _RAND_1058 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_lrs1 = _RAND_1058[5:0];
  _RAND_1059 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_lrs2 = _RAND_1059[5:0];
  _RAND_1060 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_lrs3 = _RAND_1060[5:0];
  _RAND_1061 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_ldst_val = _RAND_1061[0:0];
  _RAND_1062 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_dst_rtype = _RAND_1062[1:0];
  _RAND_1063 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_lrs1_rtype = _RAND_1063[1:0];
  _RAND_1064 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_lrs2_rtype = _RAND_1064[1:0];
  _RAND_1065 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_frs3_en = _RAND_1065[0:0];
  _RAND_1066 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_fp_val = _RAND_1066[0:0];
  _RAND_1067 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_fp_single = _RAND_1067[0:0];
  _RAND_1068 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_xcpt_pf_if = _RAND_1068[0:0];
  _RAND_1069 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_xcpt_ae_if = _RAND_1069[0:0];
  _RAND_1070 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_xcpt_ma_if = _RAND_1070[0:0];
  _RAND_1071 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_bp_debug_if = _RAND_1071[0:0];
  _RAND_1072 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_bp_xcpt_if = _RAND_1072[0:0];
  _RAND_1073 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_debug_fsrc = _RAND_1073[1:0];
  _RAND_1074 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_2_debug_tsrc = _RAND_1074[1:0];
  _RAND_1075 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_switch = _RAND_1075[0:0];
  _RAND_1076 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_switch_off = _RAND_1076[0:0];
  _RAND_1077 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_is_unicore = _RAND_1077[0:0];
  _RAND_1078 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_shift = _RAND_1078[2:0];
  _RAND_1079 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_lrs3_rtype = _RAND_1079[1:0];
  _RAND_1080 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_rflag = _RAND_1080[0:0];
  _RAND_1081 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_wflag = _RAND_1081[0:0];
  _RAND_1082 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_prflag = _RAND_1082[3:0];
  _RAND_1083 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_pwflag = _RAND_1083[3:0];
  _RAND_1084 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_pflag_busy = _RAND_1084[0:0];
  _RAND_1085 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_stale_pflag = _RAND_1085[3:0];
  _RAND_1086 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_op1_sel = _RAND_1086[3:0];
  _RAND_1087 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_op2_sel = _RAND_1087[3:0];
  _RAND_1088 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_split_num = _RAND_1088[5:0];
  _RAND_1089 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_self_index = _RAND_1089[5:0];
  _RAND_1090 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_rob_inst_idx = _RAND_1090[5:0];
  _RAND_1091 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_address_num = _RAND_1091[5:0];
  _RAND_1092 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_uopc = _RAND_1092[6:0];
  _RAND_1093 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_inst = _RAND_1093[31:0];
  _RAND_1094 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_debug_inst = _RAND_1094[31:0];
  _RAND_1095 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_is_rvc = _RAND_1095[0:0];
  _RAND_1096 = {2{`RANDOM}};
  enq_buffer_2_dec_uops_3_debug_pc = _RAND_1096[39:0];
  _RAND_1097 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_iq_type = _RAND_1097[2:0];
  _RAND_1098 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_fu_code = _RAND_1098[9:0];
  _RAND_1099 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_ctrl_br_type = _RAND_1099[3:0];
  _RAND_1100 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_ctrl_op1_sel = _RAND_1100[1:0];
  _RAND_1101 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_ctrl_op2_sel = _RAND_1101[2:0];
  _RAND_1102 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_ctrl_imm_sel = _RAND_1102[2:0];
  _RAND_1103 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_ctrl_op_fcn = _RAND_1103[3:0];
  _RAND_1104 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_ctrl_fcn_dw = _RAND_1104[0:0];
  _RAND_1105 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_ctrl_csr_cmd = _RAND_1105[2:0];
  _RAND_1106 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_ctrl_is_load = _RAND_1106[0:0];
  _RAND_1107 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_ctrl_is_sta = _RAND_1107[0:0];
  _RAND_1108 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_ctrl_is_std = _RAND_1108[0:0];
  _RAND_1109 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_ctrl_op3_sel = _RAND_1109[1:0];
  _RAND_1110 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_iw_state = _RAND_1110[1:0];
  _RAND_1111 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_iw_p1_poisoned = _RAND_1111[0:0];
  _RAND_1112 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_iw_p2_poisoned = _RAND_1112[0:0];
  _RAND_1113 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_is_br = _RAND_1113[0:0];
  _RAND_1114 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_is_jalr = _RAND_1114[0:0];
  _RAND_1115 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_is_jal = _RAND_1115[0:0];
  _RAND_1116 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_is_sfb = _RAND_1116[0:0];
  _RAND_1117 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_br_mask = _RAND_1117[11:0];
  _RAND_1118 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_br_tag = _RAND_1118[3:0];
  _RAND_1119 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_ftq_idx = _RAND_1119[4:0];
  _RAND_1120 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_edge_inst = _RAND_1120[0:0];
  _RAND_1121 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_pc_lob = _RAND_1121[5:0];
  _RAND_1122 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_taken = _RAND_1122[0:0];
  _RAND_1123 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_imm_packed = _RAND_1123[19:0];
  _RAND_1124 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_csr_addr = _RAND_1124[11:0];
  _RAND_1125 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_rob_idx = _RAND_1125[5:0];
  _RAND_1126 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_ldq_idx = _RAND_1126[4:0];
  _RAND_1127 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_stq_idx = _RAND_1127[4:0];
  _RAND_1128 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_rxq_idx = _RAND_1128[1:0];
  _RAND_1129 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_pdst = _RAND_1129[6:0];
  _RAND_1130 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_prs1 = _RAND_1130[6:0];
  _RAND_1131 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_prs2 = _RAND_1131[6:0];
  _RAND_1132 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_prs3 = _RAND_1132[6:0];
  _RAND_1133 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_ppred = _RAND_1133[4:0];
  _RAND_1134 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_prs1_busy = _RAND_1134[0:0];
  _RAND_1135 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_prs2_busy = _RAND_1135[0:0];
  _RAND_1136 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_prs3_busy = _RAND_1136[0:0];
  _RAND_1137 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_ppred_busy = _RAND_1137[0:0];
  _RAND_1138 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_stale_pdst = _RAND_1138[6:0];
  _RAND_1139 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_exception = _RAND_1139[0:0];
  _RAND_1140 = {2{`RANDOM}};
  enq_buffer_2_dec_uops_3_exc_cause = _RAND_1140[63:0];
  _RAND_1141 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_bypassable = _RAND_1141[0:0];
  _RAND_1142 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_mem_cmd = _RAND_1142[4:0];
  _RAND_1143 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_mem_size = _RAND_1143[1:0];
  _RAND_1144 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_mem_signed = _RAND_1144[0:0];
  _RAND_1145 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_is_fence = _RAND_1145[0:0];
  _RAND_1146 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_is_fencei = _RAND_1146[0:0];
  _RAND_1147 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_is_amo = _RAND_1147[0:0];
  _RAND_1148 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_uses_ldq = _RAND_1148[0:0];
  _RAND_1149 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_uses_stq = _RAND_1149[0:0];
  _RAND_1150 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_is_sys_pc2epc = _RAND_1150[0:0];
  _RAND_1151 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_is_unique = _RAND_1151[0:0];
  _RAND_1152 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_flush_on_commit = _RAND_1152[0:0];
  _RAND_1153 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_ldst_is_rs1 = _RAND_1153[0:0];
  _RAND_1154 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_ldst = _RAND_1154[5:0];
  _RAND_1155 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_lrs1 = _RAND_1155[5:0];
  _RAND_1156 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_lrs2 = _RAND_1156[5:0];
  _RAND_1157 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_lrs3 = _RAND_1157[5:0];
  _RAND_1158 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_ldst_val = _RAND_1158[0:0];
  _RAND_1159 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_dst_rtype = _RAND_1159[1:0];
  _RAND_1160 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_lrs1_rtype = _RAND_1160[1:0];
  _RAND_1161 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_lrs2_rtype = _RAND_1161[1:0];
  _RAND_1162 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_frs3_en = _RAND_1162[0:0];
  _RAND_1163 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_fp_val = _RAND_1163[0:0];
  _RAND_1164 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_fp_single = _RAND_1164[0:0];
  _RAND_1165 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_xcpt_pf_if = _RAND_1165[0:0];
  _RAND_1166 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_xcpt_ae_if = _RAND_1166[0:0];
  _RAND_1167 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_xcpt_ma_if = _RAND_1167[0:0];
  _RAND_1168 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_bp_debug_if = _RAND_1168[0:0];
  _RAND_1169 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_bp_xcpt_if = _RAND_1169[0:0];
  _RAND_1170 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_debug_fsrc = _RAND_1170[1:0];
  _RAND_1171 = {1{`RANDOM}};
  enq_buffer_2_dec_uops_3_debug_tsrc = _RAND_1171[1:0];
  _RAND_1172 = {1{`RANDOM}};
  enq_buffer_2_val_mask_0 = _RAND_1172[0:0];
  _RAND_1173 = {1{`RANDOM}};
  enq_buffer_2_val_mask_1 = _RAND_1173[0:0];
  _RAND_1174 = {1{`RANDOM}};
  enq_buffer_2_val_mask_2 = _RAND_1174[0:0];
  _RAND_1175 = {1{`RANDOM}};
  enq_buffer_2_val_mask_3 = _RAND_1175[0:0];
  _RAND_1176 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_switch = _RAND_1176[0:0];
  _RAND_1177 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_switch_off = _RAND_1177[0:0];
  _RAND_1178 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_is_unicore = _RAND_1178[0:0];
  _RAND_1179 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_shift = _RAND_1179[2:0];
  _RAND_1180 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_lrs3_rtype = _RAND_1180[1:0];
  _RAND_1181 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_rflag = _RAND_1181[0:0];
  _RAND_1182 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_wflag = _RAND_1182[0:0];
  _RAND_1183 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_prflag = _RAND_1183[3:0];
  _RAND_1184 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_pwflag = _RAND_1184[3:0];
  _RAND_1185 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_pflag_busy = _RAND_1185[0:0];
  _RAND_1186 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_stale_pflag = _RAND_1186[3:0];
  _RAND_1187 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_op1_sel = _RAND_1187[3:0];
  _RAND_1188 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_op2_sel = _RAND_1188[3:0];
  _RAND_1189 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_split_num = _RAND_1189[5:0];
  _RAND_1190 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_self_index = _RAND_1190[5:0];
  _RAND_1191 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_rob_inst_idx = _RAND_1191[5:0];
  _RAND_1192 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_address_num = _RAND_1192[5:0];
  _RAND_1193 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_uopc = _RAND_1193[6:0];
  _RAND_1194 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_inst = _RAND_1194[31:0];
  _RAND_1195 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_debug_inst = _RAND_1195[31:0];
  _RAND_1196 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_is_rvc = _RAND_1196[0:0];
  _RAND_1197 = {2{`RANDOM}};
  enq_buffer_3_dec_uops_0_debug_pc = _RAND_1197[39:0];
  _RAND_1198 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_iq_type = _RAND_1198[2:0];
  _RAND_1199 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_fu_code = _RAND_1199[9:0];
  _RAND_1200 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_ctrl_br_type = _RAND_1200[3:0];
  _RAND_1201 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_ctrl_op1_sel = _RAND_1201[1:0];
  _RAND_1202 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_ctrl_op2_sel = _RAND_1202[2:0];
  _RAND_1203 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_ctrl_imm_sel = _RAND_1203[2:0];
  _RAND_1204 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_ctrl_op_fcn = _RAND_1204[3:0];
  _RAND_1205 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_ctrl_fcn_dw = _RAND_1205[0:0];
  _RAND_1206 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_ctrl_csr_cmd = _RAND_1206[2:0];
  _RAND_1207 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_ctrl_is_load = _RAND_1207[0:0];
  _RAND_1208 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_ctrl_is_sta = _RAND_1208[0:0];
  _RAND_1209 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_ctrl_is_std = _RAND_1209[0:0];
  _RAND_1210 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_ctrl_op3_sel = _RAND_1210[1:0];
  _RAND_1211 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_iw_state = _RAND_1211[1:0];
  _RAND_1212 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_iw_p1_poisoned = _RAND_1212[0:0];
  _RAND_1213 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_iw_p2_poisoned = _RAND_1213[0:0];
  _RAND_1214 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_is_br = _RAND_1214[0:0];
  _RAND_1215 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_is_jalr = _RAND_1215[0:0];
  _RAND_1216 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_is_jal = _RAND_1216[0:0];
  _RAND_1217 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_is_sfb = _RAND_1217[0:0];
  _RAND_1218 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_br_mask = _RAND_1218[11:0];
  _RAND_1219 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_br_tag = _RAND_1219[3:0];
  _RAND_1220 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_ftq_idx = _RAND_1220[4:0];
  _RAND_1221 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_edge_inst = _RAND_1221[0:0];
  _RAND_1222 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_pc_lob = _RAND_1222[5:0];
  _RAND_1223 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_taken = _RAND_1223[0:0];
  _RAND_1224 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_imm_packed = _RAND_1224[19:0];
  _RAND_1225 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_csr_addr = _RAND_1225[11:0];
  _RAND_1226 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_rob_idx = _RAND_1226[5:0];
  _RAND_1227 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_ldq_idx = _RAND_1227[4:0];
  _RAND_1228 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_stq_idx = _RAND_1228[4:0];
  _RAND_1229 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_rxq_idx = _RAND_1229[1:0];
  _RAND_1230 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_pdst = _RAND_1230[6:0];
  _RAND_1231 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_prs1 = _RAND_1231[6:0];
  _RAND_1232 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_prs2 = _RAND_1232[6:0];
  _RAND_1233 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_prs3 = _RAND_1233[6:0];
  _RAND_1234 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_ppred = _RAND_1234[4:0];
  _RAND_1235 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_prs1_busy = _RAND_1235[0:0];
  _RAND_1236 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_prs2_busy = _RAND_1236[0:0];
  _RAND_1237 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_prs3_busy = _RAND_1237[0:0];
  _RAND_1238 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_ppred_busy = _RAND_1238[0:0];
  _RAND_1239 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_stale_pdst = _RAND_1239[6:0];
  _RAND_1240 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_exception = _RAND_1240[0:0];
  _RAND_1241 = {2{`RANDOM}};
  enq_buffer_3_dec_uops_0_exc_cause = _RAND_1241[63:0];
  _RAND_1242 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_bypassable = _RAND_1242[0:0];
  _RAND_1243 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_mem_cmd = _RAND_1243[4:0];
  _RAND_1244 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_mem_size = _RAND_1244[1:0];
  _RAND_1245 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_mem_signed = _RAND_1245[0:0];
  _RAND_1246 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_is_fence = _RAND_1246[0:0];
  _RAND_1247 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_is_fencei = _RAND_1247[0:0];
  _RAND_1248 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_is_amo = _RAND_1248[0:0];
  _RAND_1249 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_uses_ldq = _RAND_1249[0:0];
  _RAND_1250 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_uses_stq = _RAND_1250[0:0];
  _RAND_1251 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_is_sys_pc2epc = _RAND_1251[0:0];
  _RAND_1252 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_is_unique = _RAND_1252[0:0];
  _RAND_1253 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_flush_on_commit = _RAND_1253[0:0];
  _RAND_1254 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_ldst_is_rs1 = _RAND_1254[0:0];
  _RAND_1255 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_ldst = _RAND_1255[5:0];
  _RAND_1256 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_lrs1 = _RAND_1256[5:0];
  _RAND_1257 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_lrs2 = _RAND_1257[5:0];
  _RAND_1258 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_lrs3 = _RAND_1258[5:0];
  _RAND_1259 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_ldst_val = _RAND_1259[0:0];
  _RAND_1260 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_dst_rtype = _RAND_1260[1:0];
  _RAND_1261 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_lrs1_rtype = _RAND_1261[1:0];
  _RAND_1262 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_lrs2_rtype = _RAND_1262[1:0];
  _RAND_1263 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_frs3_en = _RAND_1263[0:0];
  _RAND_1264 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_fp_val = _RAND_1264[0:0];
  _RAND_1265 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_fp_single = _RAND_1265[0:0];
  _RAND_1266 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_xcpt_pf_if = _RAND_1266[0:0];
  _RAND_1267 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_xcpt_ae_if = _RAND_1267[0:0];
  _RAND_1268 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_xcpt_ma_if = _RAND_1268[0:0];
  _RAND_1269 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_bp_debug_if = _RAND_1269[0:0];
  _RAND_1270 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_bp_xcpt_if = _RAND_1270[0:0];
  _RAND_1271 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_debug_fsrc = _RAND_1271[1:0];
  _RAND_1272 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_0_debug_tsrc = _RAND_1272[1:0];
  _RAND_1273 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_switch = _RAND_1273[0:0];
  _RAND_1274 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_switch_off = _RAND_1274[0:0];
  _RAND_1275 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_is_unicore = _RAND_1275[0:0];
  _RAND_1276 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_shift = _RAND_1276[2:0];
  _RAND_1277 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_lrs3_rtype = _RAND_1277[1:0];
  _RAND_1278 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_rflag = _RAND_1278[0:0];
  _RAND_1279 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_wflag = _RAND_1279[0:0];
  _RAND_1280 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_prflag = _RAND_1280[3:0];
  _RAND_1281 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_pwflag = _RAND_1281[3:0];
  _RAND_1282 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_pflag_busy = _RAND_1282[0:0];
  _RAND_1283 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_stale_pflag = _RAND_1283[3:0];
  _RAND_1284 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_op1_sel = _RAND_1284[3:0];
  _RAND_1285 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_op2_sel = _RAND_1285[3:0];
  _RAND_1286 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_split_num = _RAND_1286[5:0];
  _RAND_1287 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_self_index = _RAND_1287[5:0];
  _RAND_1288 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_rob_inst_idx = _RAND_1288[5:0];
  _RAND_1289 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_address_num = _RAND_1289[5:0];
  _RAND_1290 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_uopc = _RAND_1290[6:0];
  _RAND_1291 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_inst = _RAND_1291[31:0];
  _RAND_1292 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_debug_inst = _RAND_1292[31:0];
  _RAND_1293 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_is_rvc = _RAND_1293[0:0];
  _RAND_1294 = {2{`RANDOM}};
  enq_buffer_3_dec_uops_1_debug_pc = _RAND_1294[39:0];
  _RAND_1295 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_iq_type = _RAND_1295[2:0];
  _RAND_1296 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_fu_code = _RAND_1296[9:0];
  _RAND_1297 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_ctrl_br_type = _RAND_1297[3:0];
  _RAND_1298 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_ctrl_op1_sel = _RAND_1298[1:0];
  _RAND_1299 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_ctrl_op2_sel = _RAND_1299[2:0];
  _RAND_1300 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_ctrl_imm_sel = _RAND_1300[2:0];
  _RAND_1301 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_ctrl_op_fcn = _RAND_1301[3:0];
  _RAND_1302 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_ctrl_fcn_dw = _RAND_1302[0:0];
  _RAND_1303 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_ctrl_csr_cmd = _RAND_1303[2:0];
  _RAND_1304 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_ctrl_is_load = _RAND_1304[0:0];
  _RAND_1305 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_ctrl_is_sta = _RAND_1305[0:0];
  _RAND_1306 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_ctrl_is_std = _RAND_1306[0:0];
  _RAND_1307 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_ctrl_op3_sel = _RAND_1307[1:0];
  _RAND_1308 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_iw_state = _RAND_1308[1:0];
  _RAND_1309 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_iw_p1_poisoned = _RAND_1309[0:0];
  _RAND_1310 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_iw_p2_poisoned = _RAND_1310[0:0];
  _RAND_1311 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_is_br = _RAND_1311[0:0];
  _RAND_1312 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_is_jalr = _RAND_1312[0:0];
  _RAND_1313 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_is_jal = _RAND_1313[0:0];
  _RAND_1314 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_is_sfb = _RAND_1314[0:0];
  _RAND_1315 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_br_mask = _RAND_1315[11:0];
  _RAND_1316 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_br_tag = _RAND_1316[3:0];
  _RAND_1317 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_ftq_idx = _RAND_1317[4:0];
  _RAND_1318 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_edge_inst = _RAND_1318[0:0];
  _RAND_1319 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_pc_lob = _RAND_1319[5:0];
  _RAND_1320 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_taken = _RAND_1320[0:0];
  _RAND_1321 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_imm_packed = _RAND_1321[19:0];
  _RAND_1322 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_csr_addr = _RAND_1322[11:0];
  _RAND_1323 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_rob_idx = _RAND_1323[5:0];
  _RAND_1324 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_ldq_idx = _RAND_1324[4:0];
  _RAND_1325 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_stq_idx = _RAND_1325[4:0];
  _RAND_1326 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_rxq_idx = _RAND_1326[1:0];
  _RAND_1327 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_pdst = _RAND_1327[6:0];
  _RAND_1328 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_prs1 = _RAND_1328[6:0];
  _RAND_1329 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_prs2 = _RAND_1329[6:0];
  _RAND_1330 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_prs3 = _RAND_1330[6:0];
  _RAND_1331 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_ppred = _RAND_1331[4:0];
  _RAND_1332 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_prs1_busy = _RAND_1332[0:0];
  _RAND_1333 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_prs2_busy = _RAND_1333[0:0];
  _RAND_1334 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_prs3_busy = _RAND_1334[0:0];
  _RAND_1335 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_ppred_busy = _RAND_1335[0:0];
  _RAND_1336 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_stale_pdst = _RAND_1336[6:0];
  _RAND_1337 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_exception = _RAND_1337[0:0];
  _RAND_1338 = {2{`RANDOM}};
  enq_buffer_3_dec_uops_1_exc_cause = _RAND_1338[63:0];
  _RAND_1339 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_bypassable = _RAND_1339[0:0];
  _RAND_1340 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_mem_cmd = _RAND_1340[4:0];
  _RAND_1341 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_mem_size = _RAND_1341[1:0];
  _RAND_1342 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_mem_signed = _RAND_1342[0:0];
  _RAND_1343 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_is_fence = _RAND_1343[0:0];
  _RAND_1344 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_is_fencei = _RAND_1344[0:0];
  _RAND_1345 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_is_amo = _RAND_1345[0:0];
  _RAND_1346 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_uses_ldq = _RAND_1346[0:0];
  _RAND_1347 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_uses_stq = _RAND_1347[0:0];
  _RAND_1348 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_is_sys_pc2epc = _RAND_1348[0:0];
  _RAND_1349 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_is_unique = _RAND_1349[0:0];
  _RAND_1350 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_flush_on_commit = _RAND_1350[0:0];
  _RAND_1351 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_ldst_is_rs1 = _RAND_1351[0:0];
  _RAND_1352 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_ldst = _RAND_1352[5:0];
  _RAND_1353 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_lrs1 = _RAND_1353[5:0];
  _RAND_1354 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_lrs2 = _RAND_1354[5:0];
  _RAND_1355 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_lrs3 = _RAND_1355[5:0];
  _RAND_1356 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_ldst_val = _RAND_1356[0:0];
  _RAND_1357 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_dst_rtype = _RAND_1357[1:0];
  _RAND_1358 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_lrs1_rtype = _RAND_1358[1:0];
  _RAND_1359 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_lrs2_rtype = _RAND_1359[1:0];
  _RAND_1360 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_frs3_en = _RAND_1360[0:0];
  _RAND_1361 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_fp_val = _RAND_1361[0:0];
  _RAND_1362 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_fp_single = _RAND_1362[0:0];
  _RAND_1363 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_xcpt_pf_if = _RAND_1363[0:0];
  _RAND_1364 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_xcpt_ae_if = _RAND_1364[0:0];
  _RAND_1365 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_xcpt_ma_if = _RAND_1365[0:0];
  _RAND_1366 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_bp_debug_if = _RAND_1366[0:0];
  _RAND_1367 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_bp_xcpt_if = _RAND_1367[0:0];
  _RAND_1368 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_debug_fsrc = _RAND_1368[1:0];
  _RAND_1369 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_1_debug_tsrc = _RAND_1369[1:0];
  _RAND_1370 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_switch = _RAND_1370[0:0];
  _RAND_1371 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_switch_off = _RAND_1371[0:0];
  _RAND_1372 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_is_unicore = _RAND_1372[0:0];
  _RAND_1373 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_shift = _RAND_1373[2:0];
  _RAND_1374 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_lrs3_rtype = _RAND_1374[1:0];
  _RAND_1375 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_rflag = _RAND_1375[0:0];
  _RAND_1376 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_wflag = _RAND_1376[0:0];
  _RAND_1377 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_prflag = _RAND_1377[3:0];
  _RAND_1378 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_pwflag = _RAND_1378[3:0];
  _RAND_1379 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_pflag_busy = _RAND_1379[0:0];
  _RAND_1380 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_stale_pflag = _RAND_1380[3:0];
  _RAND_1381 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_op1_sel = _RAND_1381[3:0];
  _RAND_1382 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_op2_sel = _RAND_1382[3:0];
  _RAND_1383 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_split_num = _RAND_1383[5:0];
  _RAND_1384 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_self_index = _RAND_1384[5:0];
  _RAND_1385 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_rob_inst_idx = _RAND_1385[5:0];
  _RAND_1386 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_address_num = _RAND_1386[5:0];
  _RAND_1387 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_uopc = _RAND_1387[6:0];
  _RAND_1388 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_inst = _RAND_1388[31:0];
  _RAND_1389 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_debug_inst = _RAND_1389[31:0];
  _RAND_1390 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_is_rvc = _RAND_1390[0:0];
  _RAND_1391 = {2{`RANDOM}};
  enq_buffer_3_dec_uops_2_debug_pc = _RAND_1391[39:0];
  _RAND_1392 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_iq_type = _RAND_1392[2:0];
  _RAND_1393 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_fu_code = _RAND_1393[9:0];
  _RAND_1394 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_ctrl_br_type = _RAND_1394[3:0];
  _RAND_1395 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_ctrl_op1_sel = _RAND_1395[1:0];
  _RAND_1396 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_ctrl_op2_sel = _RAND_1396[2:0];
  _RAND_1397 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_ctrl_imm_sel = _RAND_1397[2:0];
  _RAND_1398 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_ctrl_op_fcn = _RAND_1398[3:0];
  _RAND_1399 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_ctrl_fcn_dw = _RAND_1399[0:0];
  _RAND_1400 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_ctrl_csr_cmd = _RAND_1400[2:0];
  _RAND_1401 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_ctrl_is_load = _RAND_1401[0:0];
  _RAND_1402 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_ctrl_is_sta = _RAND_1402[0:0];
  _RAND_1403 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_ctrl_is_std = _RAND_1403[0:0];
  _RAND_1404 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_ctrl_op3_sel = _RAND_1404[1:0];
  _RAND_1405 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_iw_state = _RAND_1405[1:0];
  _RAND_1406 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_iw_p1_poisoned = _RAND_1406[0:0];
  _RAND_1407 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_iw_p2_poisoned = _RAND_1407[0:0];
  _RAND_1408 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_is_br = _RAND_1408[0:0];
  _RAND_1409 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_is_jalr = _RAND_1409[0:0];
  _RAND_1410 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_is_jal = _RAND_1410[0:0];
  _RAND_1411 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_is_sfb = _RAND_1411[0:0];
  _RAND_1412 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_br_mask = _RAND_1412[11:0];
  _RAND_1413 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_br_tag = _RAND_1413[3:0];
  _RAND_1414 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_ftq_idx = _RAND_1414[4:0];
  _RAND_1415 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_edge_inst = _RAND_1415[0:0];
  _RAND_1416 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_pc_lob = _RAND_1416[5:0];
  _RAND_1417 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_taken = _RAND_1417[0:0];
  _RAND_1418 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_imm_packed = _RAND_1418[19:0];
  _RAND_1419 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_csr_addr = _RAND_1419[11:0];
  _RAND_1420 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_rob_idx = _RAND_1420[5:0];
  _RAND_1421 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_ldq_idx = _RAND_1421[4:0];
  _RAND_1422 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_stq_idx = _RAND_1422[4:0];
  _RAND_1423 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_rxq_idx = _RAND_1423[1:0];
  _RAND_1424 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_pdst = _RAND_1424[6:0];
  _RAND_1425 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_prs1 = _RAND_1425[6:0];
  _RAND_1426 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_prs2 = _RAND_1426[6:0];
  _RAND_1427 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_prs3 = _RAND_1427[6:0];
  _RAND_1428 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_ppred = _RAND_1428[4:0];
  _RAND_1429 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_prs1_busy = _RAND_1429[0:0];
  _RAND_1430 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_prs2_busy = _RAND_1430[0:0];
  _RAND_1431 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_prs3_busy = _RAND_1431[0:0];
  _RAND_1432 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_ppred_busy = _RAND_1432[0:0];
  _RAND_1433 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_stale_pdst = _RAND_1433[6:0];
  _RAND_1434 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_exception = _RAND_1434[0:0];
  _RAND_1435 = {2{`RANDOM}};
  enq_buffer_3_dec_uops_2_exc_cause = _RAND_1435[63:0];
  _RAND_1436 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_bypassable = _RAND_1436[0:0];
  _RAND_1437 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_mem_cmd = _RAND_1437[4:0];
  _RAND_1438 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_mem_size = _RAND_1438[1:0];
  _RAND_1439 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_mem_signed = _RAND_1439[0:0];
  _RAND_1440 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_is_fence = _RAND_1440[0:0];
  _RAND_1441 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_is_fencei = _RAND_1441[0:0];
  _RAND_1442 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_is_amo = _RAND_1442[0:0];
  _RAND_1443 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_uses_ldq = _RAND_1443[0:0];
  _RAND_1444 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_uses_stq = _RAND_1444[0:0];
  _RAND_1445 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_is_sys_pc2epc = _RAND_1445[0:0];
  _RAND_1446 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_is_unique = _RAND_1446[0:0];
  _RAND_1447 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_flush_on_commit = _RAND_1447[0:0];
  _RAND_1448 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_ldst_is_rs1 = _RAND_1448[0:0];
  _RAND_1449 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_ldst = _RAND_1449[5:0];
  _RAND_1450 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_lrs1 = _RAND_1450[5:0];
  _RAND_1451 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_lrs2 = _RAND_1451[5:0];
  _RAND_1452 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_lrs3 = _RAND_1452[5:0];
  _RAND_1453 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_ldst_val = _RAND_1453[0:0];
  _RAND_1454 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_dst_rtype = _RAND_1454[1:0];
  _RAND_1455 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_lrs1_rtype = _RAND_1455[1:0];
  _RAND_1456 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_lrs2_rtype = _RAND_1456[1:0];
  _RAND_1457 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_frs3_en = _RAND_1457[0:0];
  _RAND_1458 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_fp_val = _RAND_1458[0:0];
  _RAND_1459 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_fp_single = _RAND_1459[0:0];
  _RAND_1460 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_xcpt_pf_if = _RAND_1460[0:0];
  _RAND_1461 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_xcpt_ae_if = _RAND_1461[0:0];
  _RAND_1462 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_xcpt_ma_if = _RAND_1462[0:0];
  _RAND_1463 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_bp_debug_if = _RAND_1463[0:0];
  _RAND_1464 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_bp_xcpt_if = _RAND_1464[0:0];
  _RAND_1465 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_debug_fsrc = _RAND_1465[1:0];
  _RAND_1466 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_2_debug_tsrc = _RAND_1466[1:0];
  _RAND_1467 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_switch = _RAND_1467[0:0];
  _RAND_1468 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_switch_off = _RAND_1468[0:0];
  _RAND_1469 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_is_unicore = _RAND_1469[0:0];
  _RAND_1470 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_shift = _RAND_1470[2:0];
  _RAND_1471 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_lrs3_rtype = _RAND_1471[1:0];
  _RAND_1472 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_rflag = _RAND_1472[0:0];
  _RAND_1473 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_wflag = _RAND_1473[0:0];
  _RAND_1474 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_prflag = _RAND_1474[3:0];
  _RAND_1475 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_pwflag = _RAND_1475[3:0];
  _RAND_1476 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_pflag_busy = _RAND_1476[0:0];
  _RAND_1477 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_stale_pflag = _RAND_1477[3:0];
  _RAND_1478 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_op1_sel = _RAND_1478[3:0];
  _RAND_1479 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_op2_sel = _RAND_1479[3:0];
  _RAND_1480 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_split_num = _RAND_1480[5:0];
  _RAND_1481 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_self_index = _RAND_1481[5:0];
  _RAND_1482 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_rob_inst_idx = _RAND_1482[5:0];
  _RAND_1483 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_address_num = _RAND_1483[5:0];
  _RAND_1484 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_uopc = _RAND_1484[6:0];
  _RAND_1485 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_inst = _RAND_1485[31:0];
  _RAND_1486 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_debug_inst = _RAND_1486[31:0];
  _RAND_1487 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_is_rvc = _RAND_1487[0:0];
  _RAND_1488 = {2{`RANDOM}};
  enq_buffer_3_dec_uops_3_debug_pc = _RAND_1488[39:0];
  _RAND_1489 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_iq_type = _RAND_1489[2:0];
  _RAND_1490 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_fu_code = _RAND_1490[9:0];
  _RAND_1491 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_ctrl_br_type = _RAND_1491[3:0];
  _RAND_1492 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_ctrl_op1_sel = _RAND_1492[1:0];
  _RAND_1493 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_ctrl_op2_sel = _RAND_1493[2:0];
  _RAND_1494 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_ctrl_imm_sel = _RAND_1494[2:0];
  _RAND_1495 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_ctrl_op_fcn = _RAND_1495[3:0];
  _RAND_1496 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_ctrl_fcn_dw = _RAND_1496[0:0];
  _RAND_1497 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_ctrl_csr_cmd = _RAND_1497[2:0];
  _RAND_1498 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_ctrl_is_load = _RAND_1498[0:0];
  _RAND_1499 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_ctrl_is_sta = _RAND_1499[0:0];
  _RAND_1500 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_ctrl_is_std = _RAND_1500[0:0];
  _RAND_1501 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_ctrl_op3_sel = _RAND_1501[1:0];
  _RAND_1502 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_iw_state = _RAND_1502[1:0];
  _RAND_1503 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_iw_p1_poisoned = _RAND_1503[0:0];
  _RAND_1504 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_iw_p2_poisoned = _RAND_1504[0:0];
  _RAND_1505 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_is_br = _RAND_1505[0:0];
  _RAND_1506 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_is_jalr = _RAND_1506[0:0];
  _RAND_1507 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_is_jal = _RAND_1507[0:0];
  _RAND_1508 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_is_sfb = _RAND_1508[0:0];
  _RAND_1509 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_br_mask = _RAND_1509[11:0];
  _RAND_1510 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_br_tag = _RAND_1510[3:0];
  _RAND_1511 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_ftq_idx = _RAND_1511[4:0];
  _RAND_1512 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_edge_inst = _RAND_1512[0:0];
  _RAND_1513 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_pc_lob = _RAND_1513[5:0];
  _RAND_1514 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_taken = _RAND_1514[0:0];
  _RAND_1515 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_imm_packed = _RAND_1515[19:0];
  _RAND_1516 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_csr_addr = _RAND_1516[11:0];
  _RAND_1517 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_rob_idx = _RAND_1517[5:0];
  _RAND_1518 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_ldq_idx = _RAND_1518[4:0];
  _RAND_1519 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_stq_idx = _RAND_1519[4:0];
  _RAND_1520 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_rxq_idx = _RAND_1520[1:0];
  _RAND_1521 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_pdst = _RAND_1521[6:0];
  _RAND_1522 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_prs1 = _RAND_1522[6:0];
  _RAND_1523 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_prs2 = _RAND_1523[6:0];
  _RAND_1524 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_prs3 = _RAND_1524[6:0];
  _RAND_1525 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_ppred = _RAND_1525[4:0];
  _RAND_1526 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_prs1_busy = _RAND_1526[0:0];
  _RAND_1527 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_prs2_busy = _RAND_1527[0:0];
  _RAND_1528 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_prs3_busy = _RAND_1528[0:0];
  _RAND_1529 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_ppred_busy = _RAND_1529[0:0];
  _RAND_1530 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_stale_pdst = _RAND_1530[6:0];
  _RAND_1531 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_exception = _RAND_1531[0:0];
  _RAND_1532 = {2{`RANDOM}};
  enq_buffer_3_dec_uops_3_exc_cause = _RAND_1532[63:0];
  _RAND_1533 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_bypassable = _RAND_1533[0:0];
  _RAND_1534 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_mem_cmd = _RAND_1534[4:0];
  _RAND_1535 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_mem_size = _RAND_1535[1:0];
  _RAND_1536 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_mem_signed = _RAND_1536[0:0];
  _RAND_1537 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_is_fence = _RAND_1537[0:0];
  _RAND_1538 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_is_fencei = _RAND_1538[0:0];
  _RAND_1539 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_is_amo = _RAND_1539[0:0];
  _RAND_1540 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_uses_ldq = _RAND_1540[0:0];
  _RAND_1541 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_uses_stq = _RAND_1541[0:0];
  _RAND_1542 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_is_sys_pc2epc = _RAND_1542[0:0];
  _RAND_1543 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_is_unique = _RAND_1543[0:0];
  _RAND_1544 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_flush_on_commit = _RAND_1544[0:0];
  _RAND_1545 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_ldst_is_rs1 = _RAND_1545[0:0];
  _RAND_1546 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_ldst = _RAND_1546[5:0];
  _RAND_1547 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_lrs1 = _RAND_1547[5:0];
  _RAND_1548 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_lrs2 = _RAND_1548[5:0];
  _RAND_1549 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_lrs3 = _RAND_1549[5:0];
  _RAND_1550 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_ldst_val = _RAND_1550[0:0];
  _RAND_1551 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_dst_rtype = _RAND_1551[1:0];
  _RAND_1552 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_lrs1_rtype = _RAND_1552[1:0];
  _RAND_1553 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_lrs2_rtype = _RAND_1553[1:0];
  _RAND_1554 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_frs3_en = _RAND_1554[0:0];
  _RAND_1555 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_fp_val = _RAND_1555[0:0];
  _RAND_1556 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_fp_single = _RAND_1556[0:0];
  _RAND_1557 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_xcpt_pf_if = _RAND_1557[0:0];
  _RAND_1558 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_xcpt_ae_if = _RAND_1558[0:0];
  _RAND_1559 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_xcpt_ma_if = _RAND_1559[0:0];
  _RAND_1560 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_bp_debug_if = _RAND_1560[0:0];
  _RAND_1561 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_bp_xcpt_if = _RAND_1561[0:0];
  _RAND_1562 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_debug_fsrc = _RAND_1562[1:0];
  _RAND_1563 = {1{`RANDOM}};
  enq_buffer_3_dec_uops_3_debug_tsrc = _RAND_1563[1:0];
  _RAND_1564 = {1{`RANDOM}};
  enq_buffer_3_val_mask_0 = _RAND_1564[0:0];
  _RAND_1565 = {1{`RANDOM}};
  enq_buffer_3_val_mask_1 = _RAND_1565[0:0];
  _RAND_1566 = {1{`RANDOM}};
  enq_buffer_3_val_mask_2 = _RAND_1566[0:0];
  _RAND_1567 = {1{`RANDOM}};
  enq_buffer_3_val_mask_3 = _RAND_1567[0:0];
  _RAND_1568 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_switch = _RAND_1568[0:0];
  _RAND_1569 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_switch_off = _RAND_1569[0:0];
  _RAND_1570 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_is_unicore = _RAND_1570[0:0];
  _RAND_1571 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_shift = _RAND_1571[2:0];
  _RAND_1572 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_lrs3_rtype = _RAND_1572[1:0];
  _RAND_1573 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_rflag = _RAND_1573[0:0];
  _RAND_1574 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_wflag = _RAND_1574[0:0];
  _RAND_1575 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_prflag = _RAND_1575[3:0];
  _RAND_1576 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_pwflag = _RAND_1576[3:0];
  _RAND_1577 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_pflag_busy = _RAND_1577[0:0];
  _RAND_1578 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_stale_pflag = _RAND_1578[3:0];
  _RAND_1579 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_op1_sel = _RAND_1579[3:0];
  _RAND_1580 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_op2_sel = _RAND_1580[3:0];
  _RAND_1581 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_split_num = _RAND_1581[5:0];
  _RAND_1582 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_self_index = _RAND_1582[5:0];
  _RAND_1583 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_rob_inst_idx = _RAND_1583[5:0];
  _RAND_1584 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_address_num = _RAND_1584[5:0];
  _RAND_1585 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_uopc = _RAND_1585[6:0];
  _RAND_1586 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_inst = _RAND_1586[31:0];
  _RAND_1587 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_debug_inst = _RAND_1587[31:0];
  _RAND_1588 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_is_rvc = _RAND_1588[0:0];
  _RAND_1589 = {2{`RANDOM}};
  enq_buffer_4_dec_uops_0_debug_pc = _RAND_1589[39:0];
  _RAND_1590 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_iq_type = _RAND_1590[2:0];
  _RAND_1591 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_fu_code = _RAND_1591[9:0];
  _RAND_1592 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_ctrl_br_type = _RAND_1592[3:0];
  _RAND_1593 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_ctrl_op1_sel = _RAND_1593[1:0];
  _RAND_1594 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_ctrl_op2_sel = _RAND_1594[2:0];
  _RAND_1595 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_ctrl_imm_sel = _RAND_1595[2:0];
  _RAND_1596 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_ctrl_op_fcn = _RAND_1596[3:0];
  _RAND_1597 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_ctrl_fcn_dw = _RAND_1597[0:0];
  _RAND_1598 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_ctrl_csr_cmd = _RAND_1598[2:0];
  _RAND_1599 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_ctrl_is_load = _RAND_1599[0:0];
  _RAND_1600 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_ctrl_is_sta = _RAND_1600[0:0];
  _RAND_1601 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_ctrl_is_std = _RAND_1601[0:0];
  _RAND_1602 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_ctrl_op3_sel = _RAND_1602[1:0];
  _RAND_1603 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_iw_state = _RAND_1603[1:0];
  _RAND_1604 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_iw_p1_poisoned = _RAND_1604[0:0];
  _RAND_1605 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_iw_p2_poisoned = _RAND_1605[0:0];
  _RAND_1606 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_is_br = _RAND_1606[0:0];
  _RAND_1607 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_is_jalr = _RAND_1607[0:0];
  _RAND_1608 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_is_jal = _RAND_1608[0:0];
  _RAND_1609 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_is_sfb = _RAND_1609[0:0];
  _RAND_1610 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_br_mask = _RAND_1610[11:0];
  _RAND_1611 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_br_tag = _RAND_1611[3:0];
  _RAND_1612 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_ftq_idx = _RAND_1612[4:0];
  _RAND_1613 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_edge_inst = _RAND_1613[0:0];
  _RAND_1614 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_pc_lob = _RAND_1614[5:0];
  _RAND_1615 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_taken = _RAND_1615[0:0];
  _RAND_1616 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_imm_packed = _RAND_1616[19:0];
  _RAND_1617 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_csr_addr = _RAND_1617[11:0];
  _RAND_1618 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_rob_idx = _RAND_1618[5:0];
  _RAND_1619 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_ldq_idx = _RAND_1619[4:0];
  _RAND_1620 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_stq_idx = _RAND_1620[4:0];
  _RAND_1621 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_rxq_idx = _RAND_1621[1:0];
  _RAND_1622 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_pdst = _RAND_1622[6:0];
  _RAND_1623 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_prs1 = _RAND_1623[6:0];
  _RAND_1624 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_prs2 = _RAND_1624[6:0];
  _RAND_1625 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_prs3 = _RAND_1625[6:0];
  _RAND_1626 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_ppred = _RAND_1626[4:0];
  _RAND_1627 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_prs1_busy = _RAND_1627[0:0];
  _RAND_1628 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_prs2_busy = _RAND_1628[0:0];
  _RAND_1629 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_prs3_busy = _RAND_1629[0:0];
  _RAND_1630 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_ppred_busy = _RAND_1630[0:0];
  _RAND_1631 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_stale_pdst = _RAND_1631[6:0];
  _RAND_1632 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_exception = _RAND_1632[0:0];
  _RAND_1633 = {2{`RANDOM}};
  enq_buffer_4_dec_uops_0_exc_cause = _RAND_1633[63:0];
  _RAND_1634 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_bypassable = _RAND_1634[0:0];
  _RAND_1635 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_mem_cmd = _RAND_1635[4:0];
  _RAND_1636 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_mem_size = _RAND_1636[1:0];
  _RAND_1637 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_mem_signed = _RAND_1637[0:0];
  _RAND_1638 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_is_fence = _RAND_1638[0:0];
  _RAND_1639 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_is_fencei = _RAND_1639[0:0];
  _RAND_1640 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_is_amo = _RAND_1640[0:0];
  _RAND_1641 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_uses_ldq = _RAND_1641[0:0];
  _RAND_1642 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_uses_stq = _RAND_1642[0:0];
  _RAND_1643 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_is_sys_pc2epc = _RAND_1643[0:0];
  _RAND_1644 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_is_unique = _RAND_1644[0:0];
  _RAND_1645 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_flush_on_commit = _RAND_1645[0:0];
  _RAND_1646 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_ldst_is_rs1 = _RAND_1646[0:0];
  _RAND_1647 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_ldst = _RAND_1647[5:0];
  _RAND_1648 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_lrs1 = _RAND_1648[5:0];
  _RAND_1649 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_lrs2 = _RAND_1649[5:0];
  _RAND_1650 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_lrs3 = _RAND_1650[5:0];
  _RAND_1651 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_ldst_val = _RAND_1651[0:0];
  _RAND_1652 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_dst_rtype = _RAND_1652[1:0];
  _RAND_1653 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_lrs1_rtype = _RAND_1653[1:0];
  _RAND_1654 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_lrs2_rtype = _RAND_1654[1:0];
  _RAND_1655 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_frs3_en = _RAND_1655[0:0];
  _RAND_1656 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_fp_val = _RAND_1656[0:0];
  _RAND_1657 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_fp_single = _RAND_1657[0:0];
  _RAND_1658 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_xcpt_pf_if = _RAND_1658[0:0];
  _RAND_1659 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_xcpt_ae_if = _RAND_1659[0:0];
  _RAND_1660 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_xcpt_ma_if = _RAND_1660[0:0];
  _RAND_1661 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_bp_debug_if = _RAND_1661[0:0];
  _RAND_1662 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_bp_xcpt_if = _RAND_1662[0:0];
  _RAND_1663 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_debug_fsrc = _RAND_1663[1:0];
  _RAND_1664 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_0_debug_tsrc = _RAND_1664[1:0];
  _RAND_1665 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_switch = _RAND_1665[0:0];
  _RAND_1666 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_switch_off = _RAND_1666[0:0];
  _RAND_1667 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_is_unicore = _RAND_1667[0:0];
  _RAND_1668 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_shift = _RAND_1668[2:0];
  _RAND_1669 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_lrs3_rtype = _RAND_1669[1:0];
  _RAND_1670 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_rflag = _RAND_1670[0:0];
  _RAND_1671 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_wflag = _RAND_1671[0:0];
  _RAND_1672 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_prflag = _RAND_1672[3:0];
  _RAND_1673 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_pwflag = _RAND_1673[3:0];
  _RAND_1674 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_pflag_busy = _RAND_1674[0:0];
  _RAND_1675 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_stale_pflag = _RAND_1675[3:0];
  _RAND_1676 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_op1_sel = _RAND_1676[3:0];
  _RAND_1677 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_op2_sel = _RAND_1677[3:0];
  _RAND_1678 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_split_num = _RAND_1678[5:0];
  _RAND_1679 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_self_index = _RAND_1679[5:0];
  _RAND_1680 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_rob_inst_idx = _RAND_1680[5:0];
  _RAND_1681 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_address_num = _RAND_1681[5:0];
  _RAND_1682 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_uopc = _RAND_1682[6:0];
  _RAND_1683 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_inst = _RAND_1683[31:0];
  _RAND_1684 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_debug_inst = _RAND_1684[31:0];
  _RAND_1685 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_is_rvc = _RAND_1685[0:0];
  _RAND_1686 = {2{`RANDOM}};
  enq_buffer_4_dec_uops_1_debug_pc = _RAND_1686[39:0];
  _RAND_1687 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_iq_type = _RAND_1687[2:0];
  _RAND_1688 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_fu_code = _RAND_1688[9:0];
  _RAND_1689 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_ctrl_br_type = _RAND_1689[3:0];
  _RAND_1690 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_ctrl_op1_sel = _RAND_1690[1:0];
  _RAND_1691 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_ctrl_op2_sel = _RAND_1691[2:0];
  _RAND_1692 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_ctrl_imm_sel = _RAND_1692[2:0];
  _RAND_1693 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_ctrl_op_fcn = _RAND_1693[3:0];
  _RAND_1694 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_ctrl_fcn_dw = _RAND_1694[0:0];
  _RAND_1695 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_ctrl_csr_cmd = _RAND_1695[2:0];
  _RAND_1696 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_ctrl_is_load = _RAND_1696[0:0];
  _RAND_1697 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_ctrl_is_sta = _RAND_1697[0:0];
  _RAND_1698 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_ctrl_is_std = _RAND_1698[0:0];
  _RAND_1699 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_ctrl_op3_sel = _RAND_1699[1:0];
  _RAND_1700 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_iw_state = _RAND_1700[1:0];
  _RAND_1701 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_iw_p1_poisoned = _RAND_1701[0:0];
  _RAND_1702 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_iw_p2_poisoned = _RAND_1702[0:0];
  _RAND_1703 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_is_br = _RAND_1703[0:0];
  _RAND_1704 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_is_jalr = _RAND_1704[0:0];
  _RAND_1705 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_is_jal = _RAND_1705[0:0];
  _RAND_1706 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_is_sfb = _RAND_1706[0:0];
  _RAND_1707 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_br_mask = _RAND_1707[11:0];
  _RAND_1708 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_br_tag = _RAND_1708[3:0];
  _RAND_1709 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_ftq_idx = _RAND_1709[4:0];
  _RAND_1710 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_edge_inst = _RAND_1710[0:0];
  _RAND_1711 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_pc_lob = _RAND_1711[5:0];
  _RAND_1712 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_taken = _RAND_1712[0:0];
  _RAND_1713 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_imm_packed = _RAND_1713[19:0];
  _RAND_1714 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_csr_addr = _RAND_1714[11:0];
  _RAND_1715 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_rob_idx = _RAND_1715[5:0];
  _RAND_1716 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_ldq_idx = _RAND_1716[4:0];
  _RAND_1717 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_stq_idx = _RAND_1717[4:0];
  _RAND_1718 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_rxq_idx = _RAND_1718[1:0];
  _RAND_1719 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_pdst = _RAND_1719[6:0];
  _RAND_1720 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_prs1 = _RAND_1720[6:0];
  _RAND_1721 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_prs2 = _RAND_1721[6:0];
  _RAND_1722 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_prs3 = _RAND_1722[6:0];
  _RAND_1723 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_ppred = _RAND_1723[4:0];
  _RAND_1724 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_prs1_busy = _RAND_1724[0:0];
  _RAND_1725 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_prs2_busy = _RAND_1725[0:0];
  _RAND_1726 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_prs3_busy = _RAND_1726[0:0];
  _RAND_1727 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_ppred_busy = _RAND_1727[0:0];
  _RAND_1728 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_stale_pdst = _RAND_1728[6:0];
  _RAND_1729 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_exception = _RAND_1729[0:0];
  _RAND_1730 = {2{`RANDOM}};
  enq_buffer_4_dec_uops_1_exc_cause = _RAND_1730[63:0];
  _RAND_1731 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_bypassable = _RAND_1731[0:0];
  _RAND_1732 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_mem_cmd = _RAND_1732[4:0];
  _RAND_1733 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_mem_size = _RAND_1733[1:0];
  _RAND_1734 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_mem_signed = _RAND_1734[0:0];
  _RAND_1735 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_is_fence = _RAND_1735[0:0];
  _RAND_1736 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_is_fencei = _RAND_1736[0:0];
  _RAND_1737 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_is_amo = _RAND_1737[0:0];
  _RAND_1738 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_uses_ldq = _RAND_1738[0:0];
  _RAND_1739 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_uses_stq = _RAND_1739[0:0];
  _RAND_1740 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_is_sys_pc2epc = _RAND_1740[0:0];
  _RAND_1741 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_is_unique = _RAND_1741[0:0];
  _RAND_1742 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_flush_on_commit = _RAND_1742[0:0];
  _RAND_1743 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_ldst_is_rs1 = _RAND_1743[0:0];
  _RAND_1744 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_ldst = _RAND_1744[5:0];
  _RAND_1745 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_lrs1 = _RAND_1745[5:0];
  _RAND_1746 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_lrs2 = _RAND_1746[5:0];
  _RAND_1747 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_lrs3 = _RAND_1747[5:0];
  _RAND_1748 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_ldst_val = _RAND_1748[0:0];
  _RAND_1749 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_dst_rtype = _RAND_1749[1:0];
  _RAND_1750 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_lrs1_rtype = _RAND_1750[1:0];
  _RAND_1751 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_lrs2_rtype = _RAND_1751[1:0];
  _RAND_1752 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_frs3_en = _RAND_1752[0:0];
  _RAND_1753 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_fp_val = _RAND_1753[0:0];
  _RAND_1754 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_fp_single = _RAND_1754[0:0];
  _RAND_1755 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_xcpt_pf_if = _RAND_1755[0:0];
  _RAND_1756 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_xcpt_ae_if = _RAND_1756[0:0];
  _RAND_1757 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_xcpt_ma_if = _RAND_1757[0:0];
  _RAND_1758 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_bp_debug_if = _RAND_1758[0:0];
  _RAND_1759 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_bp_xcpt_if = _RAND_1759[0:0];
  _RAND_1760 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_debug_fsrc = _RAND_1760[1:0];
  _RAND_1761 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_1_debug_tsrc = _RAND_1761[1:0];
  _RAND_1762 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_switch = _RAND_1762[0:0];
  _RAND_1763 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_switch_off = _RAND_1763[0:0];
  _RAND_1764 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_is_unicore = _RAND_1764[0:0];
  _RAND_1765 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_shift = _RAND_1765[2:0];
  _RAND_1766 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_lrs3_rtype = _RAND_1766[1:0];
  _RAND_1767 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_rflag = _RAND_1767[0:0];
  _RAND_1768 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_wflag = _RAND_1768[0:0];
  _RAND_1769 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_prflag = _RAND_1769[3:0];
  _RAND_1770 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_pwflag = _RAND_1770[3:0];
  _RAND_1771 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_pflag_busy = _RAND_1771[0:0];
  _RAND_1772 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_stale_pflag = _RAND_1772[3:0];
  _RAND_1773 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_op1_sel = _RAND_1773[3:0];
  _RAND_1774 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_op2_sel = _RAND_1774[3:0];
  _RAND_1775 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_split_num = _RAND_1775[5:0];
  _RAND_1776 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_self_index = _RAND_1776[5:0];
  _RAND_1777 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_rob_inst_idx = _RAND_1777[5:0];
  _RAND_1778 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_address_num = _RAND_1778[5:0];
  _RAND_1779 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_uopc = _RAND_1779[6:0];
  _RAND_1780 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_inst = _RAND_1780[31:0];
  _RAND_1781 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_debug_inst = _RAND_1781[31:0];
  _RAND_1782 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_is_rvc = _RAND_1782[0:0];
  _RAND_1783 = {2{`RANDOM}};
  enq_buffer_4_dec_uops_2_debug_pc = _RAND_1783[39:0];
  _RAND_1784 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_iq_type = _RAND_1784[2:0];
  _RAND_1785 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_fu_code = _RAND_1785[9:0];
  _RAND_1786 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_ctrl_br_type = _RAND_1786[3:0];
  _RAND_1787 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_ctrl_op1_sel = _RAND_1787[1:0];
  _RAND_1788 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_ctrl_op2_sel = _RAND_1788[2:0];
  _RAND_1789 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_ctrl_imm_sel = _RAND_1789[2:0];
  _RAND_1790 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_ctrl_op_fcn = _RAND_1790[3:0];
  _RAND_1791 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_ctrl_fcn_dw = _RAND_1791[0:0];
  _RAND_1792 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_ctrl_csr_cmd = _RAND_1792[2:0];
  _RAND_1793 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_ctrl_is_load = _RAND_1793[0:0];
  _RAND_1794 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_ctrl_is_sta = _RAND_1794[0:0];
  _RAND_1795 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_ctrl_is_std = _RAND_1795[0:0];
  _RAND_1796 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_ctrl_op3_sel = _RAND_1796[1:0];
  _RAND_1797 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_iw_state = _RAND_1797[1:0];
  _RAND_1798 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_iw_p1_poisoned = _RAND_1798[0:0];
  _RAND_1799 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_iw_p2_poisoned = _RAND_1799[0:0];
  _RAND_1800 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_is_br = _RAND_1800[0:0];
  _RAND_1801 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_is_jalr = _RAND_1801[0:0];
  _RAND_1802 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_is_jal = _RAND_1802[0:0];
  _RAND_1803 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_is_sfb = _RAND_1803[0:0];
  _RAND_1804 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_br_mask = _RAND_1804[11:0];
  _RAND_1805 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_br_tag = _RAND_1805[3:0];
  _RAND_1806 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_ftq_idx = _RAND_1806[4:0];
  _RAND_1807 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_edge_inst = _RAND_1807[0:0];
  _RAND_1808 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_pc_lob = _RAND_1808[5:0];
  _RAND_1809 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_taken = _RAND_1809[0:0];
  _RAND_1810 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_imm_packed = _RAND_1810[19:0];
  _RAND_1811 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_csr_addr = _RAND_1811[11:0];
  _RAND_1812 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_rob_idx = _RAND_1812[5:0];
  _RAND_1813 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_ldq_idx = _RAND_1813[4:0];
  _RAND_1814 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_stq_idx = _RAND_1814[4:0];
  _RAND_1815 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_rxq_idx = _RAND_1815[1:0];
  _RAND_1816 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_pdst = _RAND_1816[6:0];
  _RAND_1817 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_prs1 = _RAND_1817[6:0];
  _RAND_1818 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_prs2 = _RAND_1818[6:0];
  _RAND_1819 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_prs3 = _RAND_1819[6:0];
  _RAND_1820 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_ppred = _RAND_1820[4:0];
  _RAND_1821 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_prs1_busy = _RAND_1821[0:0];
  _RAND_1822 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_prs2_busy = _RAND_1822[0:0];
  _RAND_1823 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_prs3_busy = _RAND_1823[0:0];
  _RAND_1824 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_ppred_busy = _RAND_1824[0:0];
  _RAND_1825 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_stale_pdst = _RAND_1825[6:0];
  _RAND_1826 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_exception = _RAND_1826[0:0];
  _RAND_1827 = {2{`RANDOM}};
  enq_buffer_4_dec_uops_2_exc_cause = _RAND_1827[63:0];
  _RAND_1828 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_bypassable = _RAND_1828[0:0];
  _RAND_1829 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_mem_cmd = _RAND_1829[4:0];
  _RAND_1830 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_mem_size = _RAND_1830[1:0];
  _RAND_1831 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_mem_signed = _RAND_1831[0:0];
  _RAND_1832 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_is_fence = _RAND_1832[0:0];
  _RAND_1833 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_is_fencei = _RAND_1833[0:0];
  _RAND_1834 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_is_amo = _RAND_1834[0:0];
  _RAND_1835 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_uses_ldq = _RAND_1835[0:0];
  _RAND_1836 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_uses_stq = _RAND_1836[0:0];
  _RAND_1837 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_is_sys_pc2epc = _RAND_1837[0:0];
  _RAND_1838 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_is_unique = _RAND_1838[0:0];
  _RAND_1839 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_flush_on_commit = _RAND_1839[0:0];
  _RAND_1840 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_ldst_is_rs1 = _RAND_1840[0:0];
  _RAND_1841 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_ldst = _RAND_1841[5:0];
  _RAND_1842 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_lrs1 = _RAND_1842[5:0];
  _RAND_1843 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_lrs2 = _RAND_1843[5:0];
  _RAND_1844 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_lrs3 = _RAND_1844[5:0];
  _RAND_1845 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_ldst_val = _RAND_1845[0:0];
  _RAND_1846 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_dst_rtype = _RAND_1846[1:0];
  _RAND_1847 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_lrs1_rtype = _RAND_1847[1:0];
  _RAND_1848 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_lrs2_rtype = _RAND_1848[1:0];
  _RAND_1849 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_frs3_en = _RAND_1849[0:0];
  _RAND_1850 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_fp_val = _RAND_1850[0:0];
  _RAND_1851 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_fp_single = _RAND_1851[0:0];
  _RAND_1852 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_xcpt_pf_if = _RAND_1852[0:0];
  _RAND_1853 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_xcpt_ae_if = _RAND_1853[0:0];
  _RAND_1854 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_xcpt_ma_if = _RAND_1854[0:0];
  _RAND_1855 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_bp_debug_if = _RAND_1855[0:0];
  _RAND_1856 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_bp_xcpt_if = _RAND_1856[0:0];
  _RAND_1857 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_debug_fsrc = _RAND_1857[1:0];
  _RAND_1858 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_2_debug_tsrc = _RAND_1858[1:0];
  _RAND_1859 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_switch = _RAND_1859[0:0];
  _RAND_1860 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_switch_off = _RAND_1860[0:0];
  _RAND_1861 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_is_unicore = _RAND_1861[0:0];
  _RAND_1862 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_shift = _RAND_1862[2:0];
  _RAND_1863 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_lrs3_rtype = _RAND_1863[1:0];
  _RAND_1864 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_rflag = _RAND_1864[0:0];
  _RAND_1865 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_wflag = _RAND_1865[0:0];
  _RAND_1866 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_prflag = _RAND_1866[3:0];
  _RAND_1867 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_pwflag = _RAND_1867[3:0];
  _RAND_1868 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_pflag_busy = _RAND_1868[0:0];
  _RAND_1869 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_stale_pflag = _RAND_1869[3:0];
  _RAND_1870 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_op1_sel = _RAND_1870[3:0];
  _RAND_1871 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_op2_sel = _RAND_1871[3:0];
  _RAND_1872 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_split_num = _RAND_1872[5:0];
  _RAND_1873 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_self_index = _RAND_1873[5:0];
  _RAND_1874 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_rob_inst_idx = _RAND_1874[5:0];
  _RAND_1875 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_address_num = _RAND_1875[5:0];
  _RAND_1876 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_uopc = _RAND_1876[6:0];
  _RAND_1877 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_inst = _RAND_1877[31:0];
  _RAND_1878 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_debug_inst = _RAND_1878[31:0];
  _RAND_1879 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_is_rvc = _RAND_1879[0:0];
  _RAND_1880 = {2{`RANDOM}};
  enq_buffer_4_dec_uops_3_debug_pc = _RAND_1880[39:0];
  _RAND_1881 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_iq_type = _RAND_1881[2:0];
  _RAND_1882 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_fu_code = _RAND_1882[9:0];
  _RAND_1883 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_ctrl_br_type = _RAND_1883[3:0];
  _RAND_1884 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_ctrl_op1_sel = _RAND_1884[1:0];
  _RAND_1885 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_ctrl_op2_sel = _RAND_1885[2:0];
  _RAND_1886 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_ctrl_imm_sel = _RAND_1886[2:0];
  _RAND_1887 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_ctrl_op_fcn = _RAND_1887[3:0];
  _RAND_1888 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_ctrl_fcn_dw = _RAND_1888[0:0];
  _RAND_1889 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_ctrl_csr_cmd = _RAND_1889[2:0];
  _RAND_1890 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_ctrl_is_load = _RAND_1890[0:0];
  _RAND_1891 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_ctrl_is_sta = _RAND_1891[0:0];
  _RAND_1892 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_ctrl_is_std = _RAND_1892[0:0];
  _RAND_1893 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_ctrl_op3_sel = _RAND_1893[1:0];
  _RAND_1894 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_iw_state = _RAND_1894[1:0];
  _RAND_1895 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_iw_p1_poisoned = _RAND_1895[0:0];
  _RAND_1896 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_iw_p2_poisoned = _RAND_1896[0:0];
  _RAND_1897 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_is_br = _RAND_1897[0:0];
  _RAND_1898 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_is_jalr = _RAND_1898[0:0];
  _RAND_1899 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_is_jal = _RAND_1899[0:0];
  _RAND_1900 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_is_sfb = _RAND_1900[0:0];
  _RAND_1901 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_br_mask = _RAND_1901[11:0];
  _RAND_1902 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_br_tag = _RAND_1902[3:0];
  _RAND_1903 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_ftq_idx = _RAND_1903[4:0];
  _RAND_1904 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_edge_inst = _RAND_1904[0:0];
  _RAND_1905 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_pc_lob = _RAND_1905[5:0];
  _RAND_1906 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_taken = _RAND_1906[0:0];
  _RAND_1907 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_imm_packed = _RAND_1907[19:0];
  _RAND_1908 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_csr_addr = _RAND_1908[11:0];
  _RAND_1909 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_rob_idx = _RAND_1909[5:0];
  _RAND_1910 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_ldq_idx = _RAND_1910[4:0];
  _RAND_1911 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_stq_idx = _RAND_1911[4:0];
  _RAND_1912 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_rxq_idx = _RAND_1912[1:0];
  _RAND_1913 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_pdst = _RAND_1913[6:0];
  _RAND_1914 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_prs1 = _RAND_1914[6:0];
  _RAND_1915 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_prs2 = _RAND_1915[6:0];
  _RAND_1916 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_prs3 = _RAND_1916[6:0];
  _RAND_1917 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_ppred = _RAND_1917[4:0];
  _RAND_1918 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_prs1_busy = _RAND_1918[0:0];
  _RAND_1919 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_prs2_busy = _RAND_1919[0:0];
  _RAND_1920 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_prs3_busy = _RAND_1920[0:0];
  _RAND_1921 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_ppred_busy = _RAND_1921[0:0];
  _RAND_1922 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_stale_pdst = _RAND_1922[6:0];
  _RAND_1923 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_exception = _RAND_1923[0:0];
  _RAND_1924 = {2{`RANDOM}};
  enq_buffer_4_dec_uops_3_exc_cause = _RAND_1924[63:0];
  _RAND_1925 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_bypassable = _RAND_1925[0:0];
  _RAND_1926 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_mem_cmd = _RAND_1926[4:0];
  _RAND_1927 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_mem_size = _RAND_1927[1:0];
  _RAND_1928 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_mem_signed = _RAND_1928[0:0];
  _RAND_1929 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_is_fence = _RAND_1929[0:0];
  _RAND_1930 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_is_fencei = _RAND_1930[0:0];
  _RAND_1931 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_is_amo = _RAND_1931[0:0];
  _RAND_1932 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_uses_ldq = _RAND_1932[0:0];
  _RAND_1933 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_uses_stq = _RAND_1933[0:0];
  _RAND_1934 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_is_sys_pc2epc = _RAND_1934[0:0];
  _RAND_1935 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_is_unique = _RAND_1935[0:0];
  _RAND_1936 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_flush_on_commit = _RAND_1936[0:0];
  _RAND_1937 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_ldst_is_rs1 = _RAND_1937[0:0];
  _RAND_1938 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_ldst = _RAND_1938[5:0];
  _RAND_1939 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_lrs1 = _RAND_1939[5:0];
  _RAND_1940 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_lrs2 = _RAND_1940[5:0];
  _RAND_1941 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_lrs3 = _RAND_1941[5:0];
  _RAND_1942 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_ldst_val = _RAND_1942[0:0];
  _RAND_1943 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_dst_rtype = _RAND_1943[1:0];
  _RAND_1944 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_lrs1_rtype = _RAND_1944[1:0];
  _RAND_1945 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_lrs2_rtype = _RAND_1945[1:0];
  _RAND_1946 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_frs3_en = _RAND_1946[0:0];
  _RAND_1947 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_fp_val = _RAND_1947[0:0];
  _RAND_1948 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_fp_single = _RAND_1948[0:0];
  _RAND_1949 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_xcpt_pf_if = _RAND_1949[0:0];
  _RAND_1950 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_xcpt_ae_if = _RAND_1950[0:0];
  _RAND_1951 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_xcpt_ma_if = _RAND_1951[0:0];
  _RAND_1952 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_bp_debug_if = _RAND_1952[0:0];
  _RAND_1953 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_bp_xcpt_if = _RAND_1953[0:0];
  _RAND_1954 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_debug_fsrc = _RAND_1954[1:0];
  _RAND_1955 = {1{`RANDOM}};
  enq_buffer_4_dec_uops_3_debug_tsrc = _RAND_1955[1:0];
  _RAND_1956 = {1{`RANDOM}};
  enq_buffer_4_val_mask_0 = _RAND_1956[0:0];
  _RAND_1957 = {1{`RANDOM}};
  enq_buffer_4_val_mask_1 = _RAND_1957[0:0];
  _RAND_1958 = {1{`RANDOM}};
  enq_buffer_4_val_mask_2 = _RAND_1958[0:0];
  _RAND_1959 = {1{`RANDOM}};
  enq_buffer_4_val_mask_3 = _RAND_1959[0:0];
  _RAND_1960 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_switch = _RAND_1960[0:0];
  _RAND_1961 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_switch_off = _RAND_1961[0:0];
  _RAND_1962 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_is_unicore = _RAND_1962[0:0];
  _RAND_1963 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_shift = _RAND_1963[2:0];
  _RAND_1964 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_lrs3_rtype = _RAND_1964[1:0];
  _RAND_1965 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_rflag = _RAND_1965[0:0];
  _RAND_1966 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_wflag = _RAND_1966[0:0];
  _RAND_1967 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_prflag = _RAND_1967[3:0];
  _RAND_1968 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_pwflag = _RAND_1968[3:0];
  _RAND_1969 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_pflag_busy = _RAND_1969[0:0];
  _RAND_1970 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_stale_pflag = _RAND_1970[3:0];
  _RAND_1971 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_op1_sel = _RAND_1971[3:0];
  _RAND_1972 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_op2_sel = _RAND_1972[3:0];
  _RAND_1973 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_split_num = _RAND_1973[5:0];
  _RAND_1974 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_self_index = _RAND_1974[5:0];
  _RAND_1975 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_rob_inst_idx = _RAND_1975[5:0];
  _RAND_1976 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_address_num = _RAND_1976[5:0];
  _RAND_1977 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_uopc = _RAND_1977[6:0];
  _RAND_1978 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_inst = _RAND_1978[31:0];
  _RAND_1979 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_debug_inst = _RAND_1979[31:0];
  _RAND_1980 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_is_rvc = _RAND_1980[0:0];
  _RAND_1981 = {2{`RANDOM}};
  enq_buffer_5_dec_uops_0_debug_pc = _RAND_1981[39:0];
  _RAND_1982 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_iq_type = _RAND_1982[2:0];
  _RAND_1983 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_fu_code = _RAND_1983[9:0];
  _RAND_1984 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_ctrl_br_type = _RAND_1984[3:0];
  _RAND_1985 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_ctrl_op1_sel = _RAND_1985[1:0];
  _RAND_1986 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_ctrl_op2_sel = _RAND_1986[2:0];
  _RAND_1987 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_ctrl_imm_sel = _RAND_1987[2:0];
  _RAND_1988 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_ctrl_op_fcn = _RAND_1988[3:0];
  _RAND_1989 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_ctrl_fcn_dw = _RAND_1989[0:0];
  _RAND_1990 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_ctrl_csr_cmd = _RAND_1990[2:0];
  _RAND_1991 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_ctrl_is_load = _RAND_1991[0:0];
  _RAND_1992 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_ctrl_is_sta = _RAND_1992[0:0];
  _RAND_1993 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_ctrl_is_std = _RAND_1993[0:0];
  _RAND_1994 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_ctrl_op3_sel = _RAND_1994[1:0];
  _RAND_1995 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_iw_state = _RAND_1995[1:0];
  _RAND_1996 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_iw_p1_poisoned = _RAND_1996[0:0];
  _RAND_1997 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_iw_p2_poisoned = _RAND_1997[0:0];
  _RAND_1998 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_is_br = _RAND_1998[0:0];
  _RAND_1999 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_is_jalr = _RAND_1999[0:0];
  _RAND_2000 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_is_jal = _RAND_2000[0:0];
  _RAND_2001 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_is_sfb = _RAND_2001[0:0];
  _RAND_2002 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_br_mask = _RAND_2002[11:0];
  _RAND_2003 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_br_tag = _RAND_2003[3:0];
  _RAND_2004 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_ftq_idx = _RAND_2004[4:0];
  _RAND_2005 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_edge_inst = _RAND_2005[0:0];
  _RAND_2006 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_pc_lob = _RAND_2006[5:0];
  _RAND_2007 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_taken = _RAND_2007[0:0];
  _RAND_2008 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_imm_packed = _RAND_2008[19:0];
  _RAND_2009 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_csr_addr = _RAND_2009[11:0];
  _RAND_2010 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_rob_idx = _RAND_2010[5:0];
  _RAND_2011 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_ldq_idx = _RAND_2011[4:0];
  _RAND_2012 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_stq_idx = _RAND_2012[4:0];
  _RAND_2013 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_rxq_idx = _RAND_2013[1:0];
  _RAND_2014 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_pdst = _RAND_2014[6:0];
  _RAND_2015 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_prs1 = _RAND_2015[6:0];
  _RAND_2016 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_prs2 = _RAND_2016[6:0];
  _RAND_2017 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_prs3 = _RAND_2017[6:0];
  _RAND_2018 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_ppred = _RAND_2018[4:0];
  _RAND_2019 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_prs1_busy = _RAND_2019[0:0];
  _RAND_2020 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_prs2_busy = _RAND_2020[0:0];
  _RAND_2021 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_prs3_busy = _RAND_2021[0:0];
  _RAND_2022 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_ppred_busy = _RAND_2022[0:0];
  _RAND_2023 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_stale_pdst = _RAND_2023[6:0];
  _RAND_2024 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_exception = _RAND_2024[0:0];
  _RAND_2025 = {2{`RANDOM}};
  enq_buffer_5_dec_uops_0_exc_cause = _RAND_2025[63:0];
  _RAND_2026 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_bypassable = _RAND_2026[0:0];
  _RAND_2027 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_mem_cmd = _RAND_2027[4:0];
  _RAND_2028 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_mem_size = _RAND_2028[1:0];
  _RAND_2029 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_mem_signed = _RAND_2029[0:0];
  _RAND_2030 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_is_fence = _RAND_2030[0:0];
  _RAND_2031 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_is_fencei = _RAND_2031[0:0];
  _RAND_2032 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_is_amo = _RAND_2032[0:0];
  _RAND_2033 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_uses_ldq = _RAND_2033[0:0];
  _RAND_2034 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_uses_stq = _RAND_2034[0:0];
  _RAND_2035 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_is_sys_pc2epc = _RAND_2035[0:0];
  _RAND_2036 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_is_unique = _RAND_2036[0:0];
  _RAND_2037 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_flush_on_commit = _RAND_2037[0:0];
  _RAND_2038 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_ldst_is_rs1 = _RAND_2038[0:0];
  _RAND_2039 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_ldst = _RAND_2039[5:0];
  _RAND_2040 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_lrs1 = _RAND_2040[5:0];
  _RAND_2041 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_lrs2 = _RAND_2041[5:0];
  _RAND_2042 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_lrs3 = _RAND_2042[5:0];
  _RAND_2043 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_ldst_val = _RAND_2043[0:0];
  _RAND_2044 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_dst_rtype = _RAND_2044[1:0];
  _RAND_2045 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_lrs1_rtype = _RAND_2045[1:0];
  _RAND_2046 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_lrs2_rtype = _RAND_2046[1:0];
  _RAND_2047 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_frs3_en = _RAND_2047[0:0];
  _RAND_2048 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_fp_val = _RAND_2048[0:0];
  _RAND_2049 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_fp_single = _RAND_2049[0:0];
  _RAND_2050 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_xcpt_pf_if = _RAND_2050[0:0];
  _RAND_2051 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_xcpt_ae_if = _RAND_2051[0:0];
  _RAND_2052 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_xcpt_ma_if = _RAND_2052[0:0];
  _RAND_2053 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_bp_debug_if = _RAND_2053[0:0];
  _RAND_2054 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_bp_xcpt_if = _RAND_2054[0:0];
  _RAND_2055 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_debug_fsrc = _RAND_2055[1:0];
  _RAND_2056 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_0_debug_tsrc = _RAND_2056[1:0];
  _RAND_2057 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_switch = _RAND_2057[0:0];
  _RAND_2058 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_switch_off = _RAND_2058[0:0];
  _RAND_2059 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_is_unicore = _RAND_2059[0:0];
  _RAND_2060 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_shift = _RAND_2060[2:0];
  _RAND_2061 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_lrs3_rtype = _RAND_2061[1:0];
  _RAND_2062 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_rflag = _RAND_2062[0:0];
  _RAND_2063 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_wflag = _RAND_2063[0:0];
  _RAND_2064 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_prflag = _RAND_2064[3:0];
  _RAND_2065 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_pwflag = _RAND_2065[3:0];
  _RAND_2066 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_pflag_busy = _RAND_2066[0:0];
  _RAND_2067 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_stale_pflag = _RAND_2067[3:0];
  _RAND_2068 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_op1_sel = _RAND_2068[3:0];
  _RAND_2069 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_op2_sel = _RAND_2069[3:0];
  _RAND_2070 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_split_num = _RAND_2070[5:0];
  _RAND_2071 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_self_index = _RAND_2071[5:0];
  _RAND_2072 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_rob_inst_idx = _RAND_2072[5:0];
  _RAND_2073 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_address_num = _RAND_2073[5:0];
  _RAND_2074 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_uopc = _RAND_2074[6:0];
  _RAND_2075 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_inst = _RAND_2075[31:0];
  _RAND_2076 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_debug_inst = _RAND_2076[31:0];
  _RAND_2077 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_is_rvc = _RAND_2077[0:0];
  _RAND_2078 = {2{`RANDOM}};
  enq_buffer_5_dec_uops_1_debug_pc = _RAND_2078[39:0];
  _RAND_2079 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_iq_type = _RAND_2079[2:0];
  _RAND_2080 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_fu_code = _RAND_2080[9:0];
  _RAND_2081 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_ctrl_br_type = _RAND_2081[3:0];
  _RAND_2082 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_ctrl_op1_sel = _RAND_2082[1:0];
  _RAND_2083 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_ctrl_op2_sel = _RAND_2083[2:0];
  _RAND_2084 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_ctrl_imm_sel = _RAND_2084[2:0];
  _RAND_2085 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_ctrl_op_fcn = _RAND_2085[3:0];
  _RAND_2086 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_ctrl_fcn_dw = _RAND_2086[0:0];
  _RAND_2087 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_ctrl_csr_cmd = _RAND_2087[2:0];
  _RAND_2088 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_ctrl_is_load = _RAND_2088[0:0];
  _RAND_2089 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_ctrl_is_sta = _RAND_2089[0:0];
  _RAND_2090 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_ctrl_is_std = _RAND_2090[0:0];
  _RAND_2091 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_ctrl_op3_sel = _RAND_2091[1:0];
  _RAND_2092 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_iw_state = _RAND_2092[1:0];
  _RAND_2093 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_iw_p1_poisoned = _RAND_2093[0:0];
  _RAND_2094 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_iw_p2_poisoned = _RAND_2094[0:0];
  _RAND_2095 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_is_br = _RAND_2095[0:0];
  _RAND_2096 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_is_jalr = _RAND_2096[0:0];
  _RAND_2097 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_is_jal = _RAND_2097[0:0];
  _RAND_2098 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_is_sfb = _RAND_2098[0:0];
  _RAND_2099 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_br_mask = _RAND_2099[11:0];
  _RAND_2100 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_br_tag = _RAND_2100[3:0];
  _RAND_2101 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_ftq_idx = _RAND_2101[4:0];
  _RAND_2102 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_edge_inst = _RAND_2102[0:0];
  _RAND_2103 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_pc_lob = _RAND_2103[5:0];
  _RAND_2104 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_taken = _RAND_2104[0:0];
  _RAND_2105 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_imm_packed = _RAND_2105[19:0];
  _RAND_2106 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_csr_addr = _RAND_2106[11:0];
  _RAND_2107 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_rob_idx = _RAND_2107[5:0];
  _RAND_2108 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_ldq_idx = _RAND_2108[4:0];
  _RAND_2109 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_stq_idx = _RAND_2109[4:0];
  _RAND_2110 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_rxq_idx = _RAND_2110[1:0];
  _RAND_2111 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_pdst = _RAND_2111[6:0];
  _RAND_2112 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_prs1 = _RAND_2112[6:0];
  _RAND_2113 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_prs2 = _RAND_2113[6:0];
  _RAND_2114 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_prs3 = _RAND_2114[6:0];
  _RAND_2115 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_ppred = _RAND_2115[4:0];
  _RAND_2116 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_prs1_busy = _RAND_2116[0:0];
  _RAND_2117 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_prs2_busy = _RAND_2117[0:0];
  _RAND_2118 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_prs3_busy = _RAND_2118[0:0];
  _RAND_2119 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_ppred_busy = _RAND_2119[0:0];
  _RAND_2120 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_stale_pdst = _RAND_2120[6:0];
  _RAND_2121 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_exception = _RAND_2121[0:0];
  _RAND_2122 = {2{`RANDOM}};
  enq_buffer_5_dec_uops_1_exc_cause = _RAND_2122[63:0];
  _RAND_2123 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_bypassable = _RAND_2123[0:0];
  _RAND_2124 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_mem_cmd = _RAND_2124[4:0];
  _RAND_2125 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_mem_size = _RAND_2125[1:0];
  _RAND_2126 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_mem_signed = _RAND_2126[0:0];
  _RAND_2127 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_is_fence = _RAND_2127[0:0];
  _RAND_2128 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_is_fencei = _RAND_2128[0:0];
  _RAND_2129 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_is_amo = _RAND_2129[0:0];
  _RAND_2130 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_uses_ldq = _RAND_2130[0:0];
  _RAND_2131 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_uses_stq = _RAND_2131[0:0];
  _RAND_2132 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_is_sys_pc2epc = _RAND_2132[0:0];
  _RAND_2133 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_is_unique = _RAND_2133[0:0];
  _RAND_2134 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_flush_on_commit = _RAND_2134[0:0];
  _RAND_2135 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_ldst_is_rs1 = _RAND_2135[0:0];
  _RAND_2136 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_ldst = _RAND_2136[5:0];
  _RAND_2137 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_lrs1 = _RAND_2137[5:0];
  _RAND_2138 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_lrs2 = _RAND_2138[5:0];
  _RAND_2139 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_lrs3 = _RAND_2139[5:0];
  _RAND_2140 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_ldst_val = _RAND_2140[0:0];
  _RAND_2141 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_dst_rtype = _RAND_2141[1:0];
  _RAND_2142 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_lrs1_rtype = _RAND_2142[1:0];
  _RAND_2143 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_lrs2_rtype = _RAND_2143[1:0];
  _RAND_2144 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_frs3_en = _RAND_2144[0:0];
  _RAND_2145 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_fp_val = _RAND_2145[0:0];
  _RAND_2146 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_fp_single = _RAND_2146[0:0];
  _RAND_2147 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_xcpt_pf_if = _RAND_2147[0:0];
  _RAND_2148 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_xcpt_ae_if = _RAND_2148[0:0];
  _RAND_2149 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_xcpt_ma_if = _RAND_2149[0:0];
  _RAND_2150 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_bp_debug_if = _RAND_2150[0:0];
  _RAND_2151 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_bp_xcpt_if = _RAND_2151[0:0];
  _RAND_2152 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_debug_fsrc = _RAND_2152[1:0];
  _RAND_2153 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_1_debug_tsrc = _RAND_2153[1:0];
  _RAND_2154 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_switch = _RAND_2154[0:0];
  _RAND_2155 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_switch_off = _RAND_2155[0:0];
  _RAND_2156 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_is_unicore = _RAND_2156[0:0];
  _RAND_2157 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_shift = _RAND_2157[2:0];
  _RAND_2158 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_lrs3_rtype = _RAND_2158[1:0];
  _RAND_2159 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_rflag = _RAND_2159[0:0];
  _RAND_2160 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_wflag = _RAND_2160[0:0];
  _RAND_2161 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_prflag = _RAND_2161[3:0];
  _RAND_2162 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_pwflag = _RAND_2162[3:0];
  _RAND_2163 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_pflag_busy = _RAND_2163[0:0];
  _RAND_2164 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_stale_pflag = _RAND_2164[3:0];
  _RAND_2165 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_op1_sel = _RAND_2165[3:0];
  _RAND_2166 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_op2_sel = _RAND_2166[3:0];
  _RAND_2167 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_split_num = _RAND_2167[5:0];
  _RAND_2168 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_self_index = _RAND_2168[5:0];
  _RAND_2169 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_rob_inst_idx = _RAND_2169[5:0];
  _RAND_2170 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_address_num = _RAND_2170[5:0];
  _RAND_2171 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_uopc = _RAND_2171[6:0];
  _RAND_2172 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_inst = _RAND_2172[31:0];
  _RAND_2173 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_debug_inst = _RAND_2173[31:0];
  _RAND_2174 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_is_rvc = _RAND_2174[0:0];
  _RAND_2175 = {2{`RANDOM}};
  enq_buffer_5_dec_uops_2_debug_pc = _RAND_2175[39:0];
  _RAND_2176 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_iq_type = _RAND_2176[2:0];
  _RAND_2177 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_fu_code = _RAND_2177[9:0];
  _RAND_2178 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_ctrl_br_type = _RAND_2178[3:0];
  _RAND_2179 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_ctrl_op1_sel = _RAND_2179[1:0];
  _RAND_2180 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_ctrl_op2_sel = _RAND_2180[2:0];
  _RAND_2181 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_ctrl_imm_sel = _RAND_2181[2:0];
  _RAND_2182 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_ctrl_op_fcn = _RAND_2182[3:0];
  _RAND_2183 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_ctrl_fcn_dw = _RAND_2183[0:0];
  _RAND_2184 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_ctrl_csr_cmd = _RAND_2184[2:0];
  _RAND_2185 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_ctrl_is_load = _RAND_2185[0:0];
  _RAND_2186 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_ctrl_is_sta = _RAND_2186[0:0];
  _RAND_2187 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_ctrl_is_std = _RAND_2187[0:0];
  _RAND_2188 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_ctrl_op3_sel = _RAND_2188[1:0];
  _RAND_2189 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_iw_state = _RAND_2189[1:0];
  _RAND_2190 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_iw_p1_poisoned = _RAND_2190[0:0];
  _RAND_2191 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_iw_p2_poisoned = _RAND_2191[0:0];
  _RAND_2192 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_is_br = _RAND_2192[0:0];
  _RAND_2193 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_is_jalr = _RAND_2193[0:0];
  _RAND_2194 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_is_jal = _RAND_2194[0:0];
  _RAND_2195 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_is_sfb = _RAND_2195[0:0];
  _RAND_2196 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_br_mask = _RAND_2196[11:0];
  _RAND_2197 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_br_tag = _RAND_2197[3:0];
  _RAND_2198 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_ftq_idx = _RAND_2198[4:0];
  _RAND_2199 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_edge_inst = _RAND_2199[0:0];
  _RAND_2200 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_pc_lob = _RAND_2200[5:0];
  _RAND_2201 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_taken = _RAND_2201[0:0];
  _RAND_2202 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_imm_packed = _RAND_2202[19:0];
  _RAND_2203 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_csr_addr = _RAND_2203[11:0];
  _RAND_2204 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_rob_idx = _RAND_2204[5:0];
  _RAND_2205 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_ldq_idx = _RAND_2205[4:0];
  _RAND_2206 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_stq_idx = _RAND_2206[4:0];
  _RAND_2207 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_rxq_idx = _RAND_2207[1:0];
  _RAND_2208 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_pdst = _RAND_2208[6:0];
  _RAND_2209 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_prs1 = _RAND_2209[6:0];
  _RAND_2210 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_prs2 = _RAND_2210[6:0];
  _RAND_2211 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_prs3 = _RAND_2211[6:0];
  _RAND_2212 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_ppred = _RAND_2212[4:0];
  _RAND_2213 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_prs1_busy = _RAND_2213[0:0];
  _RAND_2214 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_prs2_busy = _RAND_2214[0:0];
  _RAND_2215 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_prs3_busy = _RAND_2215[0:0];
  _RAND_2216 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_ppred_busy = _RAND_2216[0:0];
  _RAND_2217 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_stale_pdst = _RAND_2217[6:0];
  _RAND_2218 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_exception = _RAND_2218[0:0];
  _RAND_2219 = {2{`RANDOM}};
  enq_buffer_5_dec_uops_2_exc_cause = _RAND_2219[63:0];
  _RAND_2220 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_bypassable = _RAND_2220[0:0];
  _RAND_2221 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_mem_cmd = _RAND_2221[4:0];
  _RAND_2222 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_mem_size = _RAND_2222[1:0];
  _RAND_2223 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_mem_signed = _RAND_2223[0:0];
  _RAND_2224 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_is_fence = _RAND_2224[0:0];
  _RAND_2225 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_is_fencei = _RAND_2225[0:0];
  _RAND_2226 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_is_amo = _RAND_2226[0:0];
  _RAND_2227 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_uses_ldq = _RAND_2227[0:0];
  _RAND_2228 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_uses_stq = _RAND_2228[0:0];
  _RAND_2229 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_is_sys_pc2epc = _RAND_2229[0:0];
  _RAND_2230 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_is_unique = _RAND_2230[0:0];
  _RAND_2231 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_flush_on_commit = _RAND_2231[0:0];
  _RAND_2232 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_ldst_is_rs1 = _RAND_2232[0:0];
  _RAND_2233 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_ldst = _RAND_2233[5:0];
  _RAND_2234 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_lrs1 = _RAND_2234[5:0];
  _RAND_2235 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_lrs2 = _RAND_2235[5:0];
  _RAND_2236 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_lrs3 = _RAND_2236[5:0];
  _RAND_2237 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_ldst_val = _RAND_2237[0:0];
  _RAND_2238 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_dst_rtype = _RAND_2238[1:0];
  _RAND_2239 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_lrs1_rtype = _RAND_2239[1:0];
  _RAND_2240 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_lrs2_rtype = _RAND_2240[1:0];
  _RAND_2241 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_frs3_en = _RAND_2241[0:0];
  _RAND_2242 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_fp_val = _RAND_2242[0:0];
  _RAND_2243 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_fp_single = _RAND_2243[0:0];
  _RAND_2244 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_xcpt_pf_if = _RAND_2244[0:0];
  _RAND_2245 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_xcpt_ae_if = _RAND_2245[0:0];
  _RAND_2246 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_xcpt_ma_if = _RAND_2246[0:0];
  _RAND_2247 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_bp_debug_if = _RAND_2247[0:0];
  _RAND_2248 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_bp_xcpt_if = _RAND_2248[0:0];
  _RAND_2249 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_debug_fsrc = _RAND_2249[1:0];
  _RAND_2250 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_2_debug_tsrc = _RAND_2250[1:0];
  _RAND_2251 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_switch = _RAND_2251[0:0];
  _RAND_2252 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_switch_off = _RAND_2252[0:0];
  _RAND_2253 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_is_unicore = _RAND_2253[0:0];
  _RAND_2254 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_shift = _RAND_2254[2:0];
  _RAND_2255 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_lrs3_rtype = _RAND_2255[1:0];
  _RAND_2256 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_rflag = _RAND_2256[0:0];
  _RAND_2257 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_wflag = _RAND_2257[0:0];
  _RAND_2258 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_prflag = _RAND_2258[3:0];
  _RAND_2259 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_pwflag = _RAND_2259[3:0];
  _RAND_2260 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_pflag_busy = _RAND_2260[0:0];
  _RAND_2261 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_stale_pflag = _RAND_2261[3:0];
  _RAND_2262 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_op1_sel = _RAND_2262[3:0];
  _RAND_2263 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_op2_sel = _RAND_2263[3:0];
  _RAND_2264 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_split_num = _RAND_2264[5:0];
  _RAND_2265 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_self_index = _RAND_2265[5:0];
  _RAND_2266 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_rob_inst_idx = _RAND_2266[5:0];
  _RAND_2267 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_address_num = _RAND_2267[5:0];
  _RAND_2268 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_uopc = _RAND_2268[6:0];
  _RAND_2269 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_inst = _RAND_2269[31:0];
  _RAND_2270 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_debug_inst = _RAND_2270[31:0];
  _RAND_2271 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_is_rvc = _RAND_2271[0:0];
  _RAND_2272 = {2{`RANDOM}};
  enq_buffer_5_dec_uops_3_debug_pc = _RAND_2272[39:0];
  _RAND_2273 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_iq_type = _RAND_2273[2:0];
  _RAND_2274 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_fu_code = _RAND_2274[9:0];
  _RAND_2275 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_ctrl_br_type = _RAND_2275[3:0];
  _RAND_2276 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_ctrl_op1_sel = _RAND_2276[1:0];
  _RAND_2277 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_ctrl_op2_sel = _RAND_2277[2:0];
  _RAND_2278 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_ctrl_imm_sel = _RAND_2278[2:0];
  _RAND_2279 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_ctrl_op_fcn = _RAND_2279[3:0];
  _RAND_2280 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_ctrl_fcn_dw = _RAND_2280[0:0];
  _RAND_2281 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_ctrl_csr_cmd = _RAND_2281[2:0];
  _RAND_2282 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_ctrl_is_load = _RAND_2282[0:0];
  _RAND_2283 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_ctrl_is_sta = _RAND_2283[0:0];
  _RAND_2284 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_ctrl_is_std = _RAND_2284[0:0];
  _RAND_2285 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_ctrl_op3_sel = _RAND_2285[1:0];
  _RAND_2286 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_iw_state = _RAND_2286[1:0];
  _RAND_2287 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_iw_p1_poisoned = _RAND_2287[0:0];
  _RAND_2288 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_iw_p2_poisoned = _RAND_2288[0:0];
  _RAND_2289 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_is_br = _RAND_2289[0:0];
  _RAND_2290 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_is_jalr = _RAND_2290[0:0];
  _RAND_2291 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_is_jal = _RAND_2291[0:0];
  _RAND_2292 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_is_sfb = _RAND_2292[0:0];
  _RAND_2293 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_br_mask = _RAND_2293[11:0];
  _RAND_2294 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_br_tag = _RAND_2294[3:0];
  _RAND_2295 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_ftq_idx = _RAND_2295[4:0];
  _RAND_2296 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_edge_inst = _RAND_2296[0:0];
  _RAND_2297 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_pc_lob = _RAND_2297[5:0];
  _RAND_2298 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_taken = _RAND_2298[0:0];
  _RAND_2299 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_imm_packed = _RAND_2299[19:0];
  _RAND_2300 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_csr_addr = _RAND_2300[11:0];
  _RAND_2301 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_rob_idx = _RAND_2301[5:0];
  _RAND_2302 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_ldq_idx = _RAND_2302[4:0];
  _RAND_2303 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_stq_idx = _RAND_2303[4:0];
  _RAND_2304 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_rxq_idx = _RAND_2304[1:0];
  _RAND_2305 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_pdst = _RAND_2305[6:0];
  _RAND_2306 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_prs1 = _RAND_2306[6:0];
  _RAND_2307 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_prs2 = _RAND_2307[6:0];
  _RAND_2308 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_prs3 = _RAND_2308[6:0];
  _RAND_2309 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_ppred = _RAND_2309[4:0];
  _RAND_2310 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_prs1_busy = _RAND_2310[0:0];
  _RAND_2311 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_prs2_busy = _RAND_2311[0:0];
  _RAND_2312 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_prs3_busy = _RAND_2312[0:0];
  _RAND_2313 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_ppred_busy = _RAND_2313[0:0];
  _RAND_2314 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_stale_pdst = _RAND_2314[6:0];
  _RAND_2315 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_exception = _RAND_2315[0:0];
  _RAND_2316 = {2{`RANDOM}};
  enq_buffer_5_dec_uops_3_exc_cause = _RAND_2316[63:0];
  _RAND_2317 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_bypassable = _RAND_2317[0:0];
  _RAND_2318 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_mem_cmd = _RAND_2318[4:0];
  _RAND_2319 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_mem_size = _RAND_2319[1:0];
  _RAND_2320 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_mem_signed = _RAND_2320[0:0];
  _RAND_2321 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_is_fence = _RAND_2321[0:0];
  _RAND_2322 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_is_fencei = _RAND_2322[0:0];
  _RAND_2323 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_is_amo = _RAND_2323[0:0];
  _RAND_2324 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_uses_ldq = _RAND_2324[0:0];
  _RAND_2325 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_uses_stq = _RAND_2325[0:0];
  _RAND_2326 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_is_sys_pc2epc = _RAND_2326[0:0];
  _RAND_2327 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_is_unique = _RAND_2327[0:0];
  _RAND_2328 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_flush_on_commit = _RAND_2328[0:0];
  _RAND_2329 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_ldst_is_rs1 = _RAND_2329[0:0];
  _RAND_2330 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_ldst = _RAND_2330[5:0];
  _RAND_2331 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_lrs1 = _RAND_2331[5:0];
  _RAND_2332 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_lrs2 = _RAND_2332[5:0];
  _RAND_2333 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_lrs3 = _RAND_2333[5:0];
  _RAND_2334 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_ldst_val = _RAND_2334[0:0];
  _RAND_2335 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_dst_rtype = _RAND_2335[1:0];
  _RAND_2336 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_lrs1_rtype = _RAND_2336[1:0];
  _RAND_2337 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_lrs2_rtype = _RAND_2337[1:0];
  _RAND_2338 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_frs3_en = _RAND_2338[0:0];
  _RAND_2339 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_fp_val = _RAND_2339[0:0];
  _RAND_2340 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_fp_single = _RAND_2340[0:0];
  _RAND_2341 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_xcpt_pf_if = _RAND_2341[0:0];
  _RAND_2342 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_xcpt_ae_if = _RAND_2342[0:0];
  _RAND_2343 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_xcpt_ma_if = _RAND_2343[0:0];
  _RAND_2344 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_bp_debug_if = _RAND_2344[0:0];
  _RAND_2345 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_bp_xcpt_if = _RAND_2345[0:0];
  _RAND_2346 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_debug_fsrc = _RAND_2346[1:0];
  _RAND_2347 = {1{`RANDOM}};
  enq_buffer_5_dec_uops_3_debug_tsrc = _RAND_2347[1:0];
  _RAND_2348 = {1{`RANDOM}};
  enq_buffer_5_val_mask_0 = _RAND_2348[0:0];
  _RAND_2349 = {1{`RANDOM}};
  enq_buffer_5_val_mask_1 = _RAND_2349[0:0];
  _RAND_2350 = {1{`RANDOM}};
  enq_buffer_5_val_mask_2 = _RAND_2350[0:0];
  _RAND_2351 = {1{`RANDOM}};
  enq_buffer_5_val_mask_3 = _RAND_2351[0:0];
  _RAND_2352 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_switch = _RAND_2352[0:0];
  _RAND_2353 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_switch_off = _RAND_2353[0:0];
  _RAND_2354 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_is_unicore = _RAND_2354[0:0];
  _RAND_2355 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_shift = _RAND_2355[2:0];
  _RAND_2356 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_lrs3_rtype = _RAND_2356[1:0];
  _RAND_2357 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_rflag = _RAND_2357[0:0];
  _RAND_2358 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_wflag = _RAND_2358[0:0];
  _RAND_2359 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_prflag = _RAND_2359[3:0];
  _RAND_2360 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_pwflag = _RAND_2360[3:0];
  _RAND_2361 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_pflag_busy = _RAND_2361[0:0];
  _RAND_2362 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_stale_pflag = _RAND_2362[3:0];
  _RAND_2363 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_op1_sel = _RAND_2363[3:0];
  _RAND_2364 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_op2_sel = _RAND_2364[3:0];
  _RAND_2365 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_split_num = _RAND_2365[5:0];
  _RAND_2366 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_self_index = _RAND_2366[5:0];
  _RAND_2367 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_rob_inst_idx = _RAND_2367[5:0];
  _RAND_2368 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_address_num = _RAND_2368[5:0];
  _RAND_2369 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_uopc = _RAND_2369[6:0];
  _RAND_2370 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_inst = _RAND_2370[31:0];
  _RAND_2371 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_debug_inst = _RAND_2371[31:0];
  _RAND_2372 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_is_rvc = _RAND_2372[0:0];
  _RAND_2373 = {2{`RANDOM}};
  enq_buffer_6_dec_uops_0_debug_pc = _RAND_2373[39:0];
  _RAND_2374 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_iq_type = _RAND_2374[2:0];
  _RAND_2375 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_fu_code = _RAND_2375[9:0];
  _RAND_2376 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_ctrl_br_type = _RAND_2376[3:0];
  _RAND_2377 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_ctrl_op1_sel = _RAND_2377[1:0];
  _RAND_2378 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_ctrl_op2_sel = _RAND_2378[2:0];
  _RAND_2379 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_ctrl_imm_sel = _RAND_2379[2:0];
  _RAND_2380 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_ctrl_op_fcn = _RAND_2380[3:0];
  _RAND_2381 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_ctrl_fcn_dw = _RAND_2381[0:0];
  _RAND_2382 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_ctrl_csr_cmd = _RAND_2382[2:0];
  _RAND_2383 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_ctrl_is_load = _RAND_2383[0:0];
  _RAND_2384 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_ctrl_is_sta = _RAND_2384[0:0];
  _RAND_2385 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_ctrl_is_std = _RAND_2385[0:0];
  _RAND_2386 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_ctrl_op3_sel = _RAND_2386[1:0];
  _RAND_2387 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_iw_state = _RAND_2387[1:0];
  _RAND_2388 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_iw_p1_poisoned = _RAND_2388[0:0];
  _RAND_2389 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_iw_p2_poisoned = _RAND_2389[0:0];
  _RAND_2390 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_is_br = _RAND_2390[0:0];
  _RAND_2391 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_is_jalr = _RAND_2391[0:0];
  _RAND_2392 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_is_jal = _RAND_2392[0:0];
  _RAND_2393 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_is_sfb = _RAND_2393[0:0];
  _RAND_2394 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_br_mask = _RAND_2394[11:0];
  _RAND_2395 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_br_tag = _RAND_2395[3:0];
  _RAND_2396 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_ftq_idx = _RAND_2396[4:0];
  _RAND_2397 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_edge_inst = _RAND_2397[0:0];
  _RAND_2398 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_pc_lob = _RAND_2398[5:0];
  _RAND_2399 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_taken = _RAND_2399[0:0];
  _RAND_2400 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_imm_packed = _RAND_2400[19:0];
  _RAND_2401 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_csr_addr = _RAND_2401[11:0];
  _RAND_2402 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_rob_idx = _RAND_2402[5:0];
  _RAND_2403 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_ldq_idx = _RAND_2403[4:0];
  _RAND_2404 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_stq_idx = _RAND_2404[4:0];
  _RAND_2405 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_rxq_idx = _RAND_2405[1:0];
  _RAND_2406 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_pdst = _RAND_2406[6:0];
  _RAND_2407 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_prs1 = _RAND_2407[6:0];
  _RAND_2408 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_prs2 = _RAND_2408[6:0];
  _RAND_2409 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_prs3 = _RAND_2409[6:0];
  _RAND_2410 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_ppred = _RAND_2410[4:0];
  _RAND_2411 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_prs1_busy = _RAND_2411[0:0];
  _RAND_2412 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_prs2_busy = _RAND_2412[0:0];
  _RAND_2413 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_prs3_busy = _RAND_2413[0:0];
  _RAND_2414 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_ppred_busy = _RAND_2414[0:0];
  _RAND_2415 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_stale_pdst = _RAND_2415[6:0];
  _RAND_2416 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_exception = _RAND_2416[0:0];
  _RAND_2417 = {2{`RANDOM}};
  enq_buffer_6_dec_uops_0_exc_cause = _RAND_2417[63:0];
  _RAND_2418 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_bypassable = _RAND_2418[0:0];
  _RAND_2419 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_mem_cmd = _RAND_2419[4:0];
  _RAND_2420 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_mem_size = _RAND_2420[1:0];
  _RAND_2421 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_mem_signed = _RAND_2421[0:0];
  _RAND_2422 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_is_fence = _RAND_2422[0:0];
  _RAND_2423 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_is_fencei = _RAND_2423[0:0];
  _RAND_2424 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_is_amo = _RAND_2424[0:0];
  _RAND_2425 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_uses_ldq = _RAND_2425[0:0];
  _RAND_2426 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_uses_stq = _RAND_2426[0:0];
  _RAND_2427 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_is_sys_pc2epc = _RAND_2427[0:0];
  _RAND_2428 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_is_unique = _RAND_2428[0:0];
  _RAND_2429 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_flush_on_commit = _RAND_2429[0:0];
  _RAND_2430 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_ldst_is_rs1 = _RAND_2430[0:0];
  _RAND_2431 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_ldst = _RAND_2431[5:0];
  _RAND_2432 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_lrs1 = _RAND_2432[5:0];
  _RAND_2433 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_lrs2 = _RAND_2433[5:0];
  _RAND_2434 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_lrs3 = _RAND_2434[5:0];
  _RAND_2435 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_ldst_val = _RAND_2435[0:0];
  _RAND_2436 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_dst_rtype = _RAND_2436[1:0];
  _RAND_2437 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_lrs1_rtype = _RAND_2437[1:0];
  _RAND_2438 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_lrs2_rtype = _RAND_2438[1:0];
  _RAND_2439 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_frs3_en = _RAND_2439[0:0];
  _RAND_2440 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_fp_val = _RAND_2440[0:0];
  _RAND_2441 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_fp_single = _RAND_2441[0:0];
  _RAND_2442 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_xcpt_pf_if = _RAND_2442[0:0];
  _RAND_2443 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_xcpt_ae_if = _RAND_2443[0:0];
  _RAND_2444 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_xcpt_ma_if = _RAND_2444[0:0];
  _RAND_2445 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_bp_debug_if = _RAND_2445[0:0];
  _RAND_2446 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_bp_xcpt_if = _RAND_2446[0:0];
  _RAND_2447 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_debug_fsrc = _RAND_2447[1:0];
  _RAND_2448 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_0_debug_tsrc = _RAND_2448[1:0];
  _RAND_2449 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_switch = _RAND_2449[0:0];
  _RAND_2450 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_switch_off = _RAND_2450[0:0];
  _RAND_2451 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_is_unicore = _RAND_2451[0:0];
  _RAND_2452 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_shift = _RAND_2452[2:0];
  _RAND_2453 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_lrs3_rtype = _RAND_2453[1:0];
  _RAND_2454 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_rflag = _RAND_2454[0:0];
  _RAND_2455 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_wflag = _RAND_2455[0:0];
  _RAND_2456 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_prflag = _RAND_2456[3:0];
  _RAND_2457 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_pwflag = _RAND_2457[3:0];
  _RAND_2458 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_pflag_busy = _RAND_2458[0:0];
  _RAND_2459 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_stale_pflag = _RAND_2459[3:0];
  _RAND_2460 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_op1_sel = _RAND_2460[3:0];
  _RAND_2461 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_op2_sel = _RAND_2461[3:0];
  _RAND_2462 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_split_num = _RAND_2462[5:0];
  _RAND_2463 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_self_index = _RAND_2463[5:0];
  _RAND_2464 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_rob_inst_idx = _RAND_2464[5:0];
  _RAND_2465 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_address_num = _RAND_2465[5:0];
  _RAND_2466 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_uopc = _RAND_2466[6:0];
  _RAND_2467 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_inst = _RAND_2467[31:0];
  _RAND_2468 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_debug_inst = _RAND_2468[31:0];
  _RAND_2469 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_is_rvc = _RAND_2469[0:0];
  _RAND_2470 = {2{`RANDOM}};
  enq_buffer_6_dec_uops_1_debug_pc = _RAND_2470[39:0];
  _RAND_2471 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_iq_type = _RAND_2471[2:0];
  _RAND_2472 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_fu_code = _RAND_2472[9:0];
  _RAND_2473 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_ctrl_br_type = _RAND_2473[3:0];
  _RAND_2474 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_ctrl_op1_sel = _RAND_2474[1:0];
  _RAND_2475 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_ctrl_op2_sel = _RAND_2475[2:0];
  _RAND_2476 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_ctrl_imm_sel = _RAND_2476[2:0];
  _RAND_2477 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_ctrl_op_fcn = _RAND_2477[3:0];
  _RAND_2478 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_ctrl_fcn_dw = _RAND_2478[0:0];
  _RAND_2479 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_ctrl_csr_cmd = _RAND_2479[2:0];
  _RAND_2480 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_ctrl_is_load = _RAND_2480[0:0];
  _RAND_2481 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_ctrl_is_sta = _RAND_2481[0:0];
  _RAND_2482 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_ctrl_is_std = _RAND_2482[0:0];
  _RAND_2483 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_ctrl_op3_sel = _RAND_2483[1:0];
  _RAND_2484 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_iw_state = _RAND_2484[1:0];
  _RAND_2485 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_iw_p1_poisoned = _RAND_2485[0:0];
  _RAND_2486 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_iw_p2_poisoned = _RAND_2486[0:0];
  _RAND_2487 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_is_br = _RAND_2487[0:0];
  _RAND_2488 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_is_jalr = _RAND_2488[0:0];
  _RAND_2489 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_is_jal = _RAND_2489[0:0];
  _RAND_2490 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_is_sfb = _RAND_2490[0:0];
  _RAND_2491 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_br_mask = _RAND_2491[11:0];
  _RAND_2492 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_br_tag = _RAND_2492[3:0];
  _RAND_2493 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_ftq_idx = _RAND_2493[4:0];
  _RAND_2494 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_edge_inst = _RAND_2494[0:0];
  _RAND_2495 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_pc_lob = _RAND_2495[5:0];
  _RAND_2496 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_taken = _RAND_2496[0:0];
  _RAND_2497 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_imm_packed = _RAND_2497[19:0];
  _RAND_2498 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_csr_addr = _RAND_2498[11:0];
  _RAND_2499 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_rob_idx = _RAND_2499[5:0];
  _RAND_2500 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_ldq_idx = _RAND_2500[4:0];
  _RAND_2501 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_stq_idx = _RAND_2501[4:0];
  _RAND_2502 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_rxq_idx = _RAND_2502[1:0];
  _RAND_2503 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_pdst = _RAND_2503[6:0];
  _RAND_2504 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_prs1 = _RAND_2504[6:0];
  _RAND_2505 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_prs2 = _RAND_2505[6:0];
  _RAND_2506 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_prs3 = _RAND_2506[6:0];
  _RAND_2507 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_ppred = _RAND_2507[4:0];
  _RAND_2508 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_prs1_busy = _RAND_2508[0:0];
  _RAND_2509 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_prs2_busy = _RAND_2509[0:0];
  _RAND_2510 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_prs3_busy = _RAND_2510[0:0];
  _RAND_2511 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_ppred_busy = _RAND_2511[0:0];
  _RAND_2512 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_stale_pdst = _RAND_2512[6:0];
  _RAND_2513 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_exception = _RAND_2513[0:0];
  _RAND_2514 = {2{`RANDOM}};
  enq_buffer_6_dec_uops_1_exc_cause = _RAND_2514[63:0];
  _RAND_2515 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_bypassable = _RAND_2515[0:0];
  _RAND_2516 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_mem_cmd = _RAND_2516[4:0];
  _RAND_2517 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_mem_size = _RAND_2517[1:0];
  _RAND_2518 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_mem_signed = _RAND_2518[0:0];
  _RAND_2519 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_is_fence = _RAND_2519[0:0];
  _RAND_2520 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_is_fencei = _RAND_2520[0:0];
  _RAND_2521 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_is_amo = _RAND_2521[0:0];
  _RAND_2522 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_uses_ldq = _RAND_2522[0:0];
  _RAND_2523 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_uses_stq = _RAND_2523[0:0];
  _RAND_2524 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_is_sys_pc2epc = _RAND_2524[0:0];
  _RAND_2525 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_is_unique = _RAND_2525[0:0];
  _RAND_2526 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_flush_on_commit = _RAND_2526[0:0];
  _RAND_2527 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_ldst_is_rs1 = _RAND_2527[0:0];
  _RAND_2528 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_ldst = _RAND_2528[5:0];
  _RAND_2529 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_lrs1 = _RAND_2529[5:0];
  _RAND_2530 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_lrs2 = _RAND_2530[5:0];
  _RAND_2531 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_lrs3 = _RAND_2531[5:0];
  _RAND_2532 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_ldst_val = _RAND_2532[0:0];
  _RAND_2533 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_dst_rtype = _RAND_2533[1:0];
  _RAND_2534 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_lrs1_rtype = _RAND_2534[1:0];
  _RAND_2535 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_lrs2_rtype = _RAND_2535[1:0];
  _RAND_2536 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_frs3_en = _RAND_2536[0:0];
  _RAND_2537 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_fp_val = _RAND_2537[0:0];
  _RAND_2538 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_fp_single = _RAND_2538[0:0];
  _RAND_2539 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_xcpt_pf_if = _RAND_2539[0:0];
  _RAND_2540 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_xcpt_ae_if = _RAND_2540[0:0];
  _RAND_2541 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_xcpt_ma_if = _RAND_2541[0:0];
  _RAND_2542 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_bp_debug_if = _RAND_2542[0:0];
  _RAND_2543 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_bp_xcpt_if = _RAND_2543[0:0];
  _RAND_2544 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_debug_fsrc = _RAND_2544[1:0];
  _RAND_2545 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_1_debug_tsrc = _RAND_2545[1:0];
  _RAND_2546 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_switch = _RAND_2546[0:0];
  _RAND_2547 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_switch_off = _RAND_2547[0:0];
  _RAND_2548 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_is_unicore = _RAND_2548[0:0];
  _RAND_2549 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_shift = _RAND_2549[2:0];
  _RAND_2550 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_lrs3_rtype = _RAND_2550[1:0];
  _RAND_2551 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_rflag = _RAND_2551[0:0];
  _RAND_2552 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_wflag = _RAND_2552[0:0];
  _RAND_2553 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_prflag = _RAND_2553[3:0];
  _RAND_2554 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_pwflag = _RAND_2554[3:0];
  _RAND_2555 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_pflag_busy = _RAND_2555[0:0];
  _RAND_2556 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_stale_pflag = _RAND_2556[3:0];
  _RAND_2557 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_op1_sel = _RAND_2557[3:0];
  _RAND_2558 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_op2_sel = _RAND_2558[3:0];
  _RAND_2559 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_split_num = _RAND_2559[5:0];
  _RAND_2560 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_self_index = _RAND_2560[5:0];
  _RAND_2561 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_rob_inst_idx = _RAND_2561[5:0];
  _RAND_2562 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_address_num = _RAND_2562[5:0];
  _RAND_2563 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_uopc = _RAND_2563[6:0];
  _RAND_2564 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_inst = _RAND_2564[31:0];
  _RAND_2565 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_debug_inst = _RAND_2565[31:0];
  _RAND_2566 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_is_rvc = _RAND_2566[0:0];
  _RAND_2567 = {2{`RANDOM}};
  enq_buffer_6_dec_uops_2_debug_pc = _RAND_2567[39:0];
  _RAND_2568 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_iq_type = _RAND_2568[2:0];
  _RAND_2569 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_fu_code = _RAND_2569[9:0];
  _RAND_2570 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_ctrl_br_type = _RAND_2570[3:0];
  _RAND_2571 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_ctrl_op1_sel = _RAND_2571[1:0];
  _RAND_2572 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_ctrl_op2_sel = _RAND_2572[2:0];
  _RAND_2573 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_ctrl_imm_sel = _RAND_2573[2:0];
  _RAND_2574 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_ctrl_op_fcn = _RAND_2574[3:0];
  _RAND_2575 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_ctrl_fcn_dw = _RAND_2575[0:0];
  _RAND_2576 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_ctrl_csr_cmd = _RAND_2576[2:0];
  _RAND_2577 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_ctrl_is_load = _RAND_2577[0:0];
  _RAND_2578 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_ctrl_is_sta = _RAND_2578[0:0];
  _RAND_2579 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_ctrl_is_std = _RAND_2579[0:0];
  _RAND_2580 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_ctrl_op3_sel = _RAND_2580[1:0];
  _RAND_2581 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_iw_state = _RAND_2581[1:0];
  _RAND_2582 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_iw_p1_poisoned = _RAND_2582[0:0];
  _RAND_2583 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_iw_p2_poisoned = _RAND_2583[0:0];
  _RAND_2584 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_is_br = _RAND_2584[0:0];
  _RAND_2585 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_is_jalr = _RAND_2585[0:0];
  _RAND_2586 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_is_jal = _RAND_2586[0:0];
  _RAND_2587 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_is_sfb = _RAND_2587[0:0];
  _RAND_2588 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_br_mask = _RAND_2588[11:0];
  _RAND_2589 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_br_tag = _RAND_2589[3:0];
  _RAND_2590 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_ftq_idx = _RAND_2590[4:0];
  _RAND_2591 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_edge_inst = _RAND_2591[0:0];
  _RAND_2592 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_pc_lob = _RAND_2592[5:0];
  _RAND_2593 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_taken = _RAND_2593[0:0];
  _RAND_2594 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_imm_packed = _RAND_2594[19:0];
  _RAND_2595 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_csr_addr = _RAND_2595[11:0];
  _RAND_2596 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_rob_idx = _RAND_2596[5:0];
  _RAND_2597 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_ldq_idx = _RAND_2597[4:0];
  _RAND_2598 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_stq_idx = _RAND_2598[4:0];
  _RAND_2599 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_rxq_idx = _RAND_2599[1:0];
  _RAND_2600 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_pdst = _RAND_2600[6:0];
  _RAND_2601 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_prs1 = _RAND_2601[6:0];
  _RAND_2602 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_prs2 = _RAND_2602[6:0];
  _RAND_2603 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_prs3 = _RAND_2603[6:0];
  _RAND_2604 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_ppred = _RAND_2604[4:0];
  _RAND_2605 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_prs1_busy = _RAND_2605[0:0];
  _RAND_2606 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_prs2_busy = _RAND_2606[0:0];
  _RAND_2607 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_prs3_busy = _RAND_2607[0:0];
  _RAND_2608 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_ppred_busy = _RAND_2608[0:0];
  _RAND_2609 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_stale_pdst = _RAND_2609[6:0];
  _RAND_2610 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_exception = _RAND_2610[0:0];
  _RAND_2611 = {2{`RANDOM}};
  enq_buffer_6_dec_uops_2_exc_cause = _RAND_2611[63:0];
  _RAND_2612 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_bypassable = _RAND_2612[0:0];
  _RAND_2613 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_mem_cmd = _RAND_2613[4:0];
  _RAND_2614 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_mem_size = _RAND_2614[1:0];
  _RAND_2615 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_mem_signed = _RAND_2615[0:0];
  _RAND_2616 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_is_fence = _RAND_2616[0:0];
  _RAND_2617 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_is_fencei = _RAND_2617[0:0];
  _RAND_2618 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_is_amo = _RAND_2618[0:0];
  _RAND_2619 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_uses_ldq = _RAND_2619[0:0];
  _RAND_2620 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_uses_stq = _RAND_2620[0:0];
  _RAND_2621 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_is_sys_pc2epc = _RAND_2621[0:0];
  _RAND_2622 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_is_unique = _RAND_2622[0:0];
  _RAND_2623 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_flush_on_commit = _RAND_2623[0:0];
  _RAND_2624 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_ldst_is_rs1 = _RAND_2624[0:0];
  _RAND_2625 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_ldst = _RAND_2625[5:0];
  _RAND_2626 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_lrs1 = _RAND_2626[5:0];
  _RAND_2627 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_lrs2 = _RAND_2627[5:0];
  _RAND_2628 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_lrs3 = _RAND_2628[5:0];
  _RAND_2629 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_ldst_val = _RAND_2629[0:0];
  _RAND_2630 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_dst_rtype = _RAND_2630[1:0];
  _RAND_2631 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_lrs1_rtype = _RAND_2631[1:0];
  _RAND_2632 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_lrs2_rtype = _RAND_2632[1:0];
  _RAND_2633 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_frs3_en = _RAND_2633[0:0];
  _RAND_2634 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_fp_val = _RAND_2634[0:0];
  _RAND_2635 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_fp_single = _RAND_2635[0:0];
  _RAND_2636 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_xcpt_pf_if = _RAND_2636[0:0];
  _RAND_2637 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_xcpt_ae_if = _RAND_2637[0:0];
  _RAND_2638 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_xcpt_ma_if = _RAND_2638[0:0];
  _RAND_2639 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_bp_debug_if = _RAND_2639[0:0];
  _RAND_2640 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_bp_xcpt_if = _RAND_2640[0:0];
  _RAND_2641 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_debug_fsrc = _RAND_2641[1:0];
  _RAND_2642 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_2_debug_tsrc = _RAND_2642[1:0];
  _RAND_2643 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_switch = _RAND_2643[0:0];
  _RAND_2644 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_switch_off = _RAND_2644[0:0];
  _RAND_2645 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_is_unicore = _RAND_2645[0:0];
  _RAND_2646 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_shift = _RAND_2646[2:0];
  _RAND_2647 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_lrs3_rtype = _RAND_2647[1:0];
  _RAND_2648 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_rflag = _RAND_2648[0:0];
  _RAND_2649 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_wflag = _RAND_2649[0:0];
  _RAND_2650 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_prflag = _RAND_2650[3:0];
  _RAND_2651 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_pwflag = _RAND_2651[3:0];
  _RAND_2652 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_pflag_busy = _RAND_2652[0:0];
  _RAND_2653 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_stale_pflag = _RAND_2653[3:0];
  _RAND_2654 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_op1_sel = _RAND_2654[3:0];
  _RAND_2655 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_op2_sel = _RAND_2655[3:0];
  _RAND_2656 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_split_num = _RAND_2656[5:0];
  _RAND_2657 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_self_index = _RAND_2657[5:0];
  _RAND_2658 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_rob_inst_idx = _RAND_2658[5:0];
  _RAND_2659 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_address_num = _RAND_2659[5:0];
  _RAND_2660 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_uopc = _RAND_2660[6:0];
  _RAND_2661 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_inst = _RAND_2661[31:0];
  _RAND_2662 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_debug_inst = _RAND_2662[31:0];
  _RAND_2663 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_is_rvc = _RAND_2663[0:0];
  _RAND_2664 = {2{`RANDOM}};
  enq_buffer_6_dec_uops_3_debug_pc = _RAND_2664[39:0];
  _RAND_2665 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_iq_type = _RAND_2665[2:0];
  _RAND_2666 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_fu_code = _RAND_2666[9:0];
  _RAND_2667 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_ctrl_br_type = _RAND_2667[3:0];
  _RAND_2668 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_ctrl_op1_sel = _RAND_2668[1:0];
  _RAND_2669 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_ctrl_op2_sel = _RAND_2669[2:0];
  _RAND_2670 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_ctrl_imm_sel = _RAND_2670[2:0];
  _RAND_2671 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_ctrl_op_fcn = _RAND_2671[3:0];
  _RAND_2672 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_ctrl_fcn_dw = _RAND_2672[0:0];
  _RAND_2673 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_ctrl_csr_cmd = _RAND_2673[2:0];
  _RAND_2674 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_ctrl_is_load = _RAND_2674[0:0];
  _RAND_2675 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_ctrl_is_sta = _RAND_2675[0:0];
  _RAND_2676 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_ctrl_is_std = _RAND_2676[0:0];
  _RAND_2677 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_ctrl_op3_sel = _RAND_2677[1:0];
  _RAND_2678 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_iw_state = _RAND_2678[1:0];
  _RAND_2679 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_iw_p1_poisoned = _RAND_2679[0:0];
  _RAND_2680 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_iw_p2_poisoned = _RAND_2680[0:0];
  _RAND_2681 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_is_br = _RAND_2681[0:0];
  _RAND_2682 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_is_jalr = _RAND_2682[0:0];
  _RAND_2683 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_is_jal = _RAND_2683[0:0];
  _RAND_2684 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_is_sfb = _RAND_2684[0:0];
  _RAND_2685 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_br_mask = _RAND_2685[11:0];
  _RAND_2686 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_br_tag = _RAND_2686[3:0];
  _RAND_2687 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_ftq_idx = _RAND_2687[4:0];
  _RAND_2688 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_edge_inst = _RAND_2688[0:0];
  _RAND_2689 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_pc_lob = _RAND_2689[5:0];
  _RAND_2690 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_taken = _RAND_2690[0:0];
  _RAND_2691 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_imm_packed = _RAND_2691[19:0];
  _RAND_2692 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_csr_addr = _RAND_2692[11:0];
  _RAND_2693 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_rob_idx = _RAND_2693[5:0];
  _RAND_2694 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_ldq_idx = _RAND_2694[4:0];
  _RAND_2695 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_stq_idx = _RAND_2695[4:0];
  _RAND_2696 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_rxq_idx = _RAND_2696[1:0];
  _RAND_2697 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_pdst = _RAND_2697[6:0];
  _RAND_2698 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_prs1 = _RAND_2698[6:0];
  _RAND_2699 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_prs2 = _RAND_2699[6:0];
  _RAND_2700 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_prs3 = _RAND_2700[6:0];
  _RAND_2701 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_ppred = _RAND_2701[4:0];
  _RAND_2702 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_prs1_busy = _RAND_2702[0:0];
  _RAND_2703 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_prs2_busy = _RAND_2703[0:0];
  _RAND_2704 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_prs3_busy = _RAND_2704[0:0];
  _RAND_2705 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_ppred_busy = _RAND_2705[0:0];
  _RAND_2706 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_stale_pdst = _RAND_2706[6:0];
  _RAND_2707 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_exception = _RAND_2707[0:0];
  _RAND_2708 = {2{`RANDOM}};
  enq_buffer_6_dec_uops_3_exc_cause = _RAND_2708[63:0];
  _RAND_2709 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_bypassable = _RAND_2709[0:0];
  _RAND_2710 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_mem_cmd = _RAND_2710[4:0];
  _RAND_2711 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_mem_size = _RAND_2711[1:0];
  _RAND_2712 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_mem_signed = _RAND_2712[0:0];
  _RAND_2713 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_is_fence = _RAND_2713[0:0];
  _RAND_2714 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_is_fencei = _RAND_2714[0:0];
  _RAND_2715 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_is_amo = _RAND_2715[0:0];
  _RAND_2716 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_uses_ldq = _RAND_2716[0:0];
  _RAND_2717 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_uses_stq = _RAND_2717[0:0];
  _RAND_2718 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_is_sys_pc2epc = _RAND_2718[0:0];
  _RAND_2719 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_is_unique = _RAND_2719[0:0];
  _RAND_2720 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_flush_on_commit = _RAND_2720[0:0];
  _RAND_2721 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_ldst_is_rs1 = _RAND_2721[0:0];
  _RAND_2722 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_ldst = _RAND_2722[5:0];
  _RAND_2723 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_lrs1 = _RAND_2723[5:0];
  _RAND_2724 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_lrs2 = _RAND_2724[5:0];
  _RAND_2725 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_lrs3 = _RAND_2725[5:0];
  _RAND_2726 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_ldst_val = _RAND_2726[0:0];
  _RAND_2727 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_dst_rtype = _RAND_2727[1:0];
  _RAND_2728 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_lrs1_rtype = _RAND_2728[1:0];
  _RAND_2729 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_lrs2_rtype = _RAND_2729[1:0];
  _RAND_2730 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_frs3_en = _RAND_2730[0:0];
  _RAND_2731 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_fp_val = _RAND_2731[0:0];
  _RAND_2732 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_fp_single = _RAND_2732[0:0];
  _RAND_2733 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_xcpt_pf_if = _RAND_2733[0:0];
  _RAND_2734 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_xcpt_ae_if = _RAND_2734[0:0];
  _RAND_2735 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_xcpt_ma_if = _RAND_2735[0:0];
  _RAND_2736 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_bp_debug_if = _RAND_2736[0:0];
  _RAND_2737 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_bp_xcpt_if = _RAND_2737[0:0];
  _RAND_2738 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_debug_fsrc = _RAND_2738[1:0];
  _RAND_2739 = {1{`RANDOM}};
  enq_buffer_6_dec_uops_3_debug_tsrc = _RAND_2739[1:0];
  _RAND_2740 = {1{`RANDOM}};
  enq_buffer_6_val_mask_0 = _RAND_2740[0:0];
  _RAND_2741 = {1{`RANDOM}};
  enq_buffer_6_val_mask_1 = _RAND_2741[0:0];
  _RAND_2742 = {1{`RANDOM}};
  enq_buffer_6_val_mask_2 = _RAND_2742[0:0];
  _RAND_2743 = {1{`RANDOM}};
  enq_buffer_6_val_mask_3 = _RAND_2743[0:0];
  _RAND_2744 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_switch = _RAND_2744[0:0];
  _RAND_2745 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_switch_off = _RAND_2745[0:0];
  _RAND_2746 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_is_unicore = _RAND_2746[0:0];
  _RAND_2747 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_shift = _RAND_2747[2:0];
  _RAND_2748 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_lrs3_rtype = _RAND_2748[1:0];
  _RAND_2749 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_rflag = _RAND_2749[0:0];
  _RAND_2750 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_wflag = _RAND_2750[0:0];
  _RAND_2751 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_prflag = _RAND_2751[3:0];
  _RAND_2752 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_pwflag = _RAND_2752[3:0];
  _RAND_2753 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_pflag_busy = _RAND_2753[0:0];
  _RAND_2754 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_stale_pflag = _RAND_2754[3:0];
  _RAND_2755 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_op1_sel = _RAND_2755[3:0];
  _RAND_2756 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_op2_sel = _RAND_2756[3:0];
  _RAND_2757 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_split_num = _RAND_2757[5:0];
  _RAND_2758 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_self_index = _RAND_2758[5:0];
  _RAND_2759 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_rob_inst_idx = _RAND_2759[5:0];
  _RAND_2760 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_address_num = _RAND_2760[5:0];
  _RAND_2761 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_uopc = _RAND_2761[6:0];
  _RAND_2762 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_inst = _RAND_2762[31:0];
  _RAND_2763 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_debug_inst = _RAND_2763[31:0];
  _RAND_2764 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_is_rvc = _RAND_2764[0:0];
  _RAND_2765 = {2{`RANDOM}};
  enq_buffer_7_dec_uops_0_debug_pc = _RAND_2765[39:0];
  _RAND_2766 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_iq_type = _RAND_2766[2:0];
  _RAND_2767 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_fu_code = _RAND_2767[9:0];
  _RAND_2768 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_ctrl_br_type = _RAND_2768[3:0];
  _RAND_2769 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_ctrl_op1_sel = _RAND_2769[1:0];
  _RAND_2770 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_ctrl_op2_sel = _RAND_2770[2:0];
  _RAND_2771 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_ctrl_imm_sel = _RAND_2771[2:0];
  _RAND_2772 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_ctrl_op_fcn = _RAND_2772[3:0];
  _RAND_2773 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_ctrl_fcn_dw = _RAND_2773[0:0];
  _RAND_2774 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_ctrl_csr_cmd = _RAND_2774[2:0];
  _RAND_2775 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_ctrl_is_load = _RAND_2775[0:0];
  _RAND_2776 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_ctrl_is_sta = _RAND_2776[0:0];
  _RAND_2777 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_ctrl_is_std = _RAND_2777[0:0];
  _RAND_2778 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_ctrl_op3_sel = _RAND_2778[1:0];
  _RAND_2779 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_iw_state = _RAND_2779[1:0];
  _RAND_2780 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_iw_p1_poisoned = _RAND_2780[0:0];
  _RAND_2781 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_iw_p2_poisoned = _RAND_2781[0:0];
  _RAND_2782 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_is_br = _RAND_2782[0:0];
  _RAND_2783 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_is_jalr = _RAND_2783[0:0];
  _RAND_2784 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_is_jal = _RAND_2784[0:0];
  _RAND_2785 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_is_sfb = _RAND_2785[0:0];
  _RAND_2786 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_br_mask = _RAND_2786[11:0];
  _RAND_2787 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_br_tag = _RAND_2787[3:0];
  _RAND_2788 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_ftq_idx = _RAND_2788[4:0];
  _RAND_2789 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_edge_inst = _RAND_2789[0:0];
  _RAND_2790 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_pc_lob = _RAND_2790[5:0];
  _RAND_2791 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_taken = _RAND_2791[0:0];
  _RAND_2792 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_imm_packed = _RAND_2792[19:0];
  _RAND_2793 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_csr_addr = _RAND_2793[11:0];
  _RAND_2794 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_rob_idx = _RAND_2794[5:0];
  _RAND_2795 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_ldq_idx = _RAND_2795[4:0];
  _RAND_2796 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_stq_idx = _RAND_2796[4:0];
  _RAND_2797 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_rxq_idx = _RAND_2797[1:0];
  _RAND_2798 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_pdst = _RAND_2798[6:0];
  _RAND_2799 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_prs1 = _RAND_2799[6:0];
  _RAND_2800 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_prs2 = _RAND_2800[6:0];
  _RAND_2801 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_prs3 = _RAND_2801[6:0];
  _RAND_2802 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_ppred = _RAND_2802[4:0];
  _RAND_2803 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_prs1_busy = _RAND_2803[0:0];
  _RAND_2804 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_prs2_busy = _RAND_2804[0:0];
  _RAND_2805 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_prs3_busy = _RAND_2805[0:0];
  _RAND_2806 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_ppred_busy = _RAND_2806[0:0];
  _RAND_2807 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_stale_pdst = _RAND_2807[6:0];
  _RAND_2808 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_exception = _RAND_2808[0:0];
  _RAND_2809 = {2{`RANDOM}};
  enq_buffer_7_dec_uops_0_exc_cause = _RAND_2809[63:0];
  _RAND_2810 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_bypassable = _RAND_2810[0:0];
  _RAND_2811 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_mem_cmd = _RAND_2811[4:0];
  _RAND_2812 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_mem_size = _RAND_2812[1:0];
  _RAND_2813 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_mem_signed = _RAND_2813[0:0];
  _RAND_2814 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_is_fence = _RAND_2814[0:0];
  _RAND_2815 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_is_fencei = _RAND_2815[0:0];
  _RAND_2816 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_is_amo = _RAND_2816[0:0];
  _RAND_2817 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_uses_ldq = _RAND_2817[0:0];
  _RAND_2818 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_uses_stq = _RAND_2818[0:0];
  _RAND_2819 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_is_sys_pc2epc = _RAND_2819[0:0];
  _RAND_2820 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_is_unique = _RAND_2820[0:0];
  _RAND_2821 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_flush_on_commit = _RAND_2821[0:0];
  _RAND_2822 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_ldst_is_rs1 = _RAND_2822[0:0];
  _RAND_2823 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_ldst = _RAND_2823[5:0];
  _RAND_2824 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_lrs1 = _RAND_2824[5:0];
  _RAND_2825 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_lrs2 = _RAND_2825[5:0];
  _RAND_2826 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_lrs3 = _RAND_2826[5:0];
  _RAND_2827 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_ldst_val = _RAND_2827[0:0];
  _RAND_2828 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_dst_rtype = _RAND_2828[1:0];
  _RAND_2829 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_lrs1_rtype = _RAND_2829[1:0];
  _RAND_2830 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_lrs2_rtype = _RAND_2830[1:0];
  _RAND_2831 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_frs3_en = _RAND_2831[0:0];
  _RAND_2832 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_fp_val = _RAND_2832[0:0];
  _RAND_2833 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_fp_single = _RAND_2833[0:0];
  _RAND_2834 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_xcpt_pf_if = _RAND_2834[0:0];
  _RAND_2835 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_xcpt_ae_if = _RAND_2835[0:0];
  _RAND_2836 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_xcpt_ma_if = _RAND_2836[0:0];
  _RAND_2837 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_bp_debug_if = _RAND_2837[0:0];
  _RAND_2838 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_bp_xcpt_if = _RAND_2838[0:0];
  _RAND_2839 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_debug_fsrc = _RAND_2839[1:0];
  _RAND_2840 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_0_debug_tsrc = _RAND_2840[1:0];
  _RAND_2841 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_switch = _RAND_2841[0:0];
  _RAND_2842 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_switch_off = _RAND_2842[0:0];
  _RAND_2843 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_is_unicore = _RAND_2843[0:0];
  _RAND_2844 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_shift = _RAND_2844[2:0];
  _RAND_2845 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_lrs3_rtype = _RAND_2845[1:0];
  _RAND_2846 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_rflag = _RAND_2846[0:0];
  _RAND_2847 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_wflag = _RAND_2847[0:0];
  _RAND_2848 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_prflag = _RAND_2848[3:0];
  _RAND_2849 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_pwflag = _RAND_2849[3:0];
  _RAND_2850 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_pflag_busy = _RAND_2850[0:0];
  _RAND_2851 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_stale_pflag = _RAND_2851[3:0];
  _RAND_2852 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_op1_sel = _RAND_2852[3:0];
  _RAND_2853 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_op2_sel = _RAND_2853[3:0];
  _RAND_2854 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_split_num = _RAND_2854[5:0];
  _RAND_2855 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_self_index = _RAND_2855[5:0];
  _RAND_2856 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_rob_inst_idx = _RAND_2856[5:0];
  _RAND_2857 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_address_num = _RAND_2857[5:0];
  _RAND_2858 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_uopc = _RAND_2858[6:0];
  _RAND_2859 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_inst = _RAND_2859[31:0];
  _RAND_2860 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_debug_inst = _RAND_2860[31:0];
  _RAND_2861 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_is_rvc = _RAND_2861[0:0];
  _RAND_2862 = {2{`RANDOM}};
  enq_buffer_7_dec_uops_1_debug_pc = _RAND_2862[39:0];
  _RAND_2863 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_iq_type = _RAND_2863[2:0];
  _RAND_2864 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_fu_code = _RAND_2864[9:0];
  _RAND_2865 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_ctrl_br_type = _RAND_2865[3:0];
  _RAND_2866 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_ctrl_op1_sel = _RAND_2866[1:0];
  _RAND_2867 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_ctrl_op2_sel = _RAND_2867[2:0];
  _RAND_2868 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_ctrl_imm_sel = _RAND_2868[2:0];
  _RAND_2869 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_ctrl_op_fcn = _RAND_2869[3:0];
  _RAND_2870 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_ctrl_fcn_dw = _RAND_2870[0:0];
  _RAND_2871 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_ctrl_csr_cmd = _RAND_2871[2:0];
  _RAND_2872 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_ctrl_is_load = _RAND_2872[0:0];
  _RAND_2873 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_ctrl_is_sta = _RAND_2873[0:0];
  _RAND_2874 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_ctrl_is_std = _RAND_2874[0:0];
  _RAND_2875 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_ctrl_op3_sel = _RAND_2875[1:0];
  _RAND_2876 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_iw_state = _RAND_2876[1:0];
  _RAND_2877 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_iw_p1_poisoned = _RAND_2877[0:0];
  _RAND_2878 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_iw_p2_poisoned = _RAND_2878[0:0];
  _RAND_2879 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_is_br = _RAND_2879[0:0];
  _RAND_2880 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_is_jalr = _RAND_2880[0:0];
  _RAND_2881 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_is_jal = _RAND_2881[0:0];
  _RAND_2882 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_is_sfb = _RAND_2882[0:0];
  _RAND_2883 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_br_mask = _RAND_2883[11:0];
  _RAND_2884 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_br_tag = _RAND_2884[3:0];
  _RAND_2885 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_ftq_idx = _RAND_2885[4:0];
  _RAND_2886 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_edge_inst = _RAND_2886[0:0];
  _RAND_2887 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_pc_lob = _RAND_2887[5:0];
  _RAND_2888 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_taken = _RAND_2888[0:0];
  _RAND_2889 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_imm_packed = _RAND_2889[19:0];
  _RAND_2890 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_csr_addr = _RAND_2890[11:0];
  _RAND_2891 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_rob_idx = _RAND_2891[5:0];
  _RAND_2892 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_ldq_idx = _RAND_2892[4:0];
  _RAND_2893 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_stq_idx = _RAND_2893[4:0];
  _RAND_2894 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_rxq_idx = _RAND_2894[1:0];
  _RAND_2895 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_pdst = _RAND_2895[6:0];
  _RAND_2896 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_prs1 = _RAND_2896[6:0];
  _RAND_2897 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_prs2 = _RAND_2897[6:0];
  _RAND_2898 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_prs3 = _RAND_2898[6:0];
  _RAND_2899 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_ppred = _RAND_2899[4:0];
  _RAND_2900 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_prs1_busy = _RAND_2900[0:0];
  _RAND_2901 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_prs2_busy = _RAND_2901[0:0];
  _RAND_2902 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_prs3_busy = _RAND_2902[0:0];
  _RAND_2903 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_ppred_busy = _RAND_2903[0:0];
  _RAND_2904 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_stale_pdst = _RAND_2904[6:0];
  _RAND_2905 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_exception = _RAND_2905[0:0];
  _RAND_2906 = {2{`RANDOM}};
  enq_buffer_7_dec_uops_1_exc_cause = _RAND_2906[63:0];
  _RAND_2907 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_bypassable = _RAND_2907[0:0];
  _RAND_2908 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_mem_cmd = _RAND_2908[4:0];
  _RAND_2909 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_mem_size = _RAND_2909[1:0];
  _RAND_2910 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_mem_signed = _RAND_2910[0:0];
  _RAND_2911 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_is_fence = _RAND_2911[0:0];
  _RAND_2912 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_is_fencei = _RAND_2912[0:0];
  _RAND_2913 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_is_amo = _RAND_2913[0:0];
  _RAND_2914 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_uses_ldq = _RAND_2914[0:0];
  _RAND_2915 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_uses_stq = _RAND_2915[0:0];
  _RAND_2916 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_is_sys_pc2epc = _RAND_2916[0:0];
  _RAND_2917 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_is_unique = _RAND_2917[0:0];
  _RAND_2918 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_flush_on_commit = _RAND_2918[0:0];
  _RAND_2919 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_ldst_is_rs1 = _RAND_2919[0:0];
  _RAND_2920 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_ldst = _RAND_2920[5:0];
  _RAND_2921 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_lrs1 = _RAND_2921[5:0];
  _RAND_2922 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_lrs2 = _RAND_2922[5:0];
  _RAND_2923 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_lrs3 = _RAND_2923[5:0];
  _RAND_2924 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_ldst_val = _RAND_2924[0:0];
  _RAND_2925 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_dst_rtype = _RAND_2925[1:0];
  _RAND_2926 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_lrs1_rtype = _RAND_2926[1:0];
  _RAND_2927 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_lrs2_rtype = _RAND_2927[1:0];
  _RAND_2928 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_frs3_en = _RAND_2928[0:0];
  _RAND_2929 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_fp_val = _RAND_2929[0:0];
  _RAND_2930 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_fp_single = _RAND_2930[0:0];
  _RAND_2931 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_xcpt_pf_if = _RAND_2931[0:0];
  _RAND_2932 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_xcpt_ae_if = _RAND_2932[0:0];
  _RAND_2933 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_xcpt_ma_if = _RAND_2933[0:0];
  _RAND_2934 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_bp_debug_if = _RAND_2934[0:0];
  _RAND_2935 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_bp_xcpt_if = _RAND_2935[0:0];
  _RAND_2936 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_debug_fsrc = _RAND_2936[1:0];
  _RAND_2937 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_1_debug_tsrc = _RAND_2937[1:0];
  _RAND_2938 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_switch = _RAND_2938[0:0];
  _RAND_2939 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_switch_off = _RAND_2939[0:0];
  _RAND_2940 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_is_unicore = _RAND_2940[0:0];
  _RAND_2941 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_shift = _RAND_2941[2:0];
  _RAND_2942 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_lrs3_rtype = _RAND_2942[1:0];
  _RAND_2943 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_rflag = _RAND_2943[0:0];
  _RAND_2944 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_wflag = _RAND_2944[0:0];
  _RAND_2945 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_prflag = _RAND_2945[3:0];
  _RAND_2946 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_pwflag = _RAND_2946[3:0];
  _RAND_2947 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_pflag_busy = _RAND_2947[0:0];
  _RAND_2948 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_stale_pflag = _RAND_2948[3:0];
  _RAND_2949 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_op1_sel = _RAND_2949[3:0];
  _RAND_2950 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_op2_sel = _RAND_2950[3:0];
  _RAND_2951 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_split_num = _RAND_2951[5:0];
  _RAND_2952 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_self_index = _RAND_2952[5:0];
  _RAND_2953 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_rob_inst_idx = _RAND_2953[5:0];
  _RAND_2954 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_address_num = _RAND_2954[5:0];
  _RAND_2955 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_uopc = _RAND_2955[6:0];
  _RAND_2956 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_inst = _RAND_2956[31:0];
  _RAND_2957 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_debug_inst = _RAND_2957[31:0];
  _RAND_2958 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_is_rvc = _RAND_2958[0:0];
  _RAND_2959 = {2{`RANDOM}};
  enq_buffer_7_dec_uops_2_debug_pc = _RAND_2959[39:0];
  _RAND_2960 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_iq_type = _RAND_2960[2:0];
  _RAND_2961 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_fu_code = _RAND_2961[9:0];
  _RAND_2962 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_ctrl_br_type = _RAND_2962[3:0];
  _RAND_2963 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_ctrl_op1_sel = _RAND_2963[1:0];
  _RAND_2964 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_ctrl_op2_sel = _RAND_2964[2:0];
  _RAND_2965 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_ctrl_imm_sel = _RAND_2965[2:0];
  _RAND_2966 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_ctrl_op_fcn = _RAND_2966[3:0];
  _RAND_2967 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_ctrl_fcn_dw = _RAND_2967[0:0];
  _RAND_2968 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_ctrl_csr_cmd = _RAND_2968[2:0];
  _RAND_2969 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_ctrl_is_load = _RAND_2969[0:0];
  _RAND_2970 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_ctrl_is_sta = _RAND_2970[0:0];
  _RAND_2971 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_ctrl_is_std = _RAND_2971[0:0];
  _RAND_2972 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_ctrl_op3_sel = _RAND_2972[1:0];
  _RAND_2973 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_iw_state = _RAND_2973[1:0];
  _RAND_2974 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_iw_p1_poisoned = _RAND_2974[0:0];
  _RAND_2975 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_iw_p2_poisoned = _RAND_2975[0:0];
  _RAND_2976 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_is_br = _RAND_2976[0:0];
  _RAND_2977 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_is_jalr = _RAND_2977[0:0];
  _RAND_2978 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_is_jal = _RAND_2978[0:0];
  _RAND_2979 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_is_sfb = _RAND_2979[0:0];
  _RAND_2980 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_br_mask = _RAND_2980[11:0];
  _RAND_2981 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_br_tag = _RAND_2981[3:0];
  _RAND_2982 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_ftq_idx = _RAND_2982[4:0];
  _RAND_2983 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_edge_inst = _RAND_2983[0:0];
  _RAND_2984 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_pc_lob = _RAND_2984[5:0];
  _RAND_2985 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_taken = _RAND_2985[0:0];
  _RAND_2986 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_imm_packed = _RAND_2986[19:0];
  _RAND_2987 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_csr_addr = _RAND_2987[11:0];
  _RAND_2988 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_rob_idx = _RAND_2988[5:0];
  _RAND_2989 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_ldq_idx = _RAND_2989[4:0];
  _RAND_2990 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_stq_idx = _RAND_2990[4:0];
  _RAND_2991 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_rxq_idx = _RAND_2991[1:0];
  _RAND_2992 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_pdst = _RAND_2992[6:0];
  _RAND_2993 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_prs1 = _RAND_2993[6:0];
  _RAND_2994 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_prs2 = _RAND_2994[6:0];
  _RAND_2995 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_prs3 = _RAND_2995[6:0];
  _RAND_2996 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_ppred = _RAND_2996[4:0];
  _RAND_2997 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_prs1_busy = _RAND_2997[0:0];
  _RAND_2998 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_prs2_busy = _RAND_2998[0:0];
  _RAND_2999 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_prs3_busy = _RAND_2999[0:0];
  _RAND_3000 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_ppred_busy = _RAND_3000[0:0];
  _RAND_3001 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_stale_pdst = _RAND_3001[6:0];
  _RAND_3002 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_exception = _RAND_3002[0:0];
  _RAND_3003 = {2{`RANDOM}};
  enq_buffer_7_dec_uops_2_exc_cause = _RAND_3003[63:0];
  _RAND_3004 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_bypassable = _RAND_3004[0:0];
  _RAND_3005 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_mem_cmd = _RAND_3005[4:0];
  _RAND_3006 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_mem_size = _RAND_3006[1:0];
  _RAND_3007 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_mem_signed = _RAND_3007[0:0];
  _RAND_3008 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_is_fence = _RAND_3008[0:0];
  _RAND_3009 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_is_fencei = _RAND_3009[0:0];
  _RAND_3010 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_is_amo = _RAND_3010[0:0];
  _RAND_3011 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_uses_ldq = _RAND_3011[0:0];
  _RAND_3012 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_uses_stq = _RAND_3012[0:0];
  _RAND_3013 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_is_sys_pc2epc = _RAND_3013[0:0];
  _RAND_3014 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_is_unique = _RAND_3014[0:0];
  _RAND_3015 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_flush_on_commit = _RAND_3015[0:0];
  _RAND_3016 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_ldst_is_rs1 = _RAND_3016[0:0];
  _RAND_3017 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_ldst = _RAND_3017[5:0];
  _RAND_3018 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_lrs1 = _RAND_3018[5:0];
  _RAND_3019 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_lrs2 = _RAND_3019[5:0];
  _RAND_3020 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_lrs3 = _RAND_3020[5:0];
  _RAND_3021 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_ldst_val = _RAND_3021[0:0];
  _RAND_3022 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_dst_rtype = _RAND_3022[1:0];
  _RAND_3023 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_lrs1_rtype = _RAND_3023[1:0];
  _RAND_3024 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_lrs2_rtype = _RAND_3024[1:0];
  _RAND_3025 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_frs3_en = _RAND_3025[0:0];
  _RAND_3026 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_fp_val = _RAND_3026[0:0];
  _RAND_3027 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_fp_single = _RAND_3027[0:0];
  _RAND_3028 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_xcpt_pf_if = _RAND_3028[0:0];
  _RAND_3029 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_xcpt_ae_if = _RAND_3029[0:0];
  _RAND_3030 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_xcpt_ma_if = _RAND_3030[0:0];
  _RAND_3031 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_bp_debug_if = _RAND_3031[0:0];
  _RAND_3032 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_bp_xcpt_if = _RAND_3032[0:0];
  _RAND_3033 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_debug_fsrc = _RAND_3033[1:0];
  _RAND_3034 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_2_debug_tsrc = _RAND_3034[1:0];
  _RAND_3035 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_switch = _RAND_3035[0:0];
  _RAND_3036 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_switch_off = _RAND_3036[0:0];
  _RAND_3037 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_is_unicore = _RAND_3037[0:0];
  _RAND_3038 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_shift = _RAND_3038[2:0];
  _RAND_3039 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_lrs3_rtype = _RAND_3039[1:0];
  _RAND_3040 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_rflag = _RAND_3040[0:0];
  _RAND_3041 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_wflag = _RAND_3041[0:0];
  _RAND_3042 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_prflag = _RAND_3042[3:0];
  _RAND_3043 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_pwflag = _RAND_3043[3:0];
  _RAND_3044 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_pflag_busy = _RAND_3044[0:0];
  _RAND_3045 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_stale_pflag = _RAND_3045[3:0];
  _RAND_3046 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_op1_sel = _RAND_3046[3:0];
  _RAND_3047 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_op2_sel = _RAND_3047[3:0];
  _RAND_3048 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_split_num = _RAND_3048[5:0];
  _RAND_3049 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_self_index = _RAND_3049[5:0];
  _RAND_3050 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_rob_inst_idx = _RAND_3050[5:0];
  _RAND_3051 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_address_num = _RAND_3051[5:0];
  _RAND_3052 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_uopc = _RAND_3052[6:0];
  _RAND_3053 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_inst = _RAND_3053[31:0];
  _RAND_3054 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_debug_inst = _RAND_3054[31:0];
  _RAND_3055 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_is_rvc = _RAND_3055[0:0];
  _RAND_3056 = {2{`RANDOM}};
  enq_buffer_7_dec_uops_3_debug_pc = _RAND_3056[39:0];
  _RAND_3057 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_iq_type = _RAND_3057[2:0];
  _RAND_3058 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_fu_code = _RAND_3058[9:0];
  _RAND_3059 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_ctrl_br_type = _RAND_3059[3:0];
  _RAND_3060 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_ctrl_op1_sel = _RAND_3060[1:0];
  _RAND_3061 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_ctrl_op2_sel = _RAND_3061[2:0];
  _RAND_3062 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_ctrl_imm_sel = _RAND_3062[2:0];
  _RAND_3063 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_ctrl_op_fcn = _RAND_3063[3:0];
  _RAND_3064 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_ctrl_fcn_dw = _RAND_3064[0:0];
  _RAND_3065 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_ctrl_csr_cmd = _RAND_3065[2:0];
  _RAND_3066 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_ctrl_is_load = _RAND_3066[0:0];
  _RAND_3067 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_ctrl_is_sta = _RAND_3067[0:0];
  _RAND_3068 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_ctrl_is_std = _RAND_3068[0:0];
  _RAND_3069 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_ctrl_op3_sel = _RAND_3069[1:0];
  _RAND_3070 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_iw_state = _RAND_3070[1:0];
  _RAND_3071 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_iw_p1_poisoned = _RAND_3071[0:0];
  _RAND_3072 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_iw_p2_poisoned = _RAND_3072[0:0];
  _RAND_3073 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_is_br = _RAND_3073[0:0];
  _RAND_3074 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_is_jalr = _RAND_3074[0:0];
  _RAND_3075 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_is_jal = _RAND_3075[0:0];
  _RAND_3076 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_is_sfb = _RAND_3076[0:0];
  _RAND_3077 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_br_mask = _RAND_3077[11:0];
  _RAND_3078 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_br_tag = _RAND_3078[3:0];
  _RAND_3079 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_ftq_idx = _RAND_3079[4:0];
  _RAND_3080 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_edge_inst = _RAND_3080[0:0];
  _RAND_3081 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_pc_lob = _RAND_3081[5:0];
  _RAND_3082 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_taken = _RAND_3082[0:0];
  _RAND_3083 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_imm_packed = _RAND_3083[19:0];
  _RAND_3084 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_csr_addr = _RAND_3084[11:0];
  _RAND_3085 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_rob_idx = _RAND_3085[5:0];
  _RAND_3086 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_ldq_idx = _RAND_3086[4:0];
  _RAND_3087 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_stq_idx = _RAND_3087[4:0];
  _RAND_3088 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_rxq_idx = _RAND_3088[1:0];
  _RAND_3089 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_pdst = _RAND_3089[6:0];
  _RAND_3090 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_prs1 = _RAND_3090[6:0];
  _RAND_3091 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_prs2 = _RAND_3091[6:0];
  _RAND_3092 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_prs3 = _RAND_3092[6:0];
  _RAND_3093 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_ppred = _RAND_3093[4:0];
  _RAND_3094 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_prs1_busy = _RAND_3094[0:0];
  _RAND_3095 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_prs2_busy = _RAND_3095[0:0];
  _RAND_3096 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_prs3_busy = _RAND_3096[0:0];
  _RAND_3097 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_ppred_busy = _RAND_3097[0:0];
  _RAND_3098 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_stale_pdst = _RAND_3098[6:0];
  _RAND_3099 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_exception = _RAND_3099[0:0];
  _RAND_3100 = {2{`RANDOM}};
  enq_buffer_7_dec_uops_3_exc_cause = _RAND_3100[63:0];
  _RAND_3101 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_bypassable = _RAND_3101[0:0];
  _RAND_3102 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_mem_cmd = _RAND_3102[4:0];
  _RAND_3103 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_mem_size = _RAND_3103[1:0];
  _RAND_3104 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_mem_signed = _RAND_3104[0:0];
  _RAND_3105 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_is_fence = _RAND_3105[0:0];
  _RAND_3106 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_is_fencei = _RAND_3106[0:0];
  _RAND_3107 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_is_amo = _RAND_3107[0:0];
  _RAND_3108 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_uses_ldq = _RAND_3108[0:0];
  _RAND_3109 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_uses_stq = _RAND_3109[0:0];
  _RAND_3110 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_is_sys_pc2epc = _RAND_3110[0:0];
  _RAND_3111 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_is_unique = _RAND_3111[0:0];
  _RAND_3112 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_flush_on_commit = _RAND_3112[0:0];
  _RAND_3113 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_ldst_is_rs1 = _RAND_3113[0:0];
  _RAND_3114 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_ldst = _RAND_3114[5:0];
  _RAND_3115 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_lrs1 = _RAND_3115[5:0];
  _RAND_3116 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_lrs2 = _RAND_3116[5:0];
  _RAND_3117 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_lrs3 = _RAND_3117[5:0];
  _RAND_3118 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_ldst_val = _RAND_3118[0:0];
  _RAND_3119 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_dst_rtype = _RAND_3119[1:0];
  _RAND_3120 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_lrs1_rtype = _RAND_3120[1:0];
  _RAND_3121 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_lrs2_rtype = _RAND_3121[1:0];
  _RAND_3122 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_frs3_en = _RAND_3122[0:0];
  _RAND_3123 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_fp_val = _RAND_3123[0:0];
  _RAND_3124 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_fp_single = _RAND_3124[0:0];
  _RAND_3125 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_xcpt_pf_if = _RAND_3125[0:0];
  _RAND_3126 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_xcpt_ae_if = _RAND_3126[0:0];
  _RAND_3127 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_xcpt_ma_if = _RAND_3127[0:0];
  _RAND_3128 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_bp_debug_if = _RAND_3128[0:0];
  _RAND_3129 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_bp_xcpt_if = _RAND_3129[0:0];
  _RAND_3130 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_debug_fsrc = _RAND_3130[1:0];
  _RAND_3131 = {1{`RANDOM}};
  enq_buffer_7_dec_uops_3_debug_tsrc = _RAND_3131[1:0];
  _RAND_3132 = {1{`RANDOM}};
  enq_buffer_7_val_mask_0 = _RAND_3132[0:0];
  _RAND_3133 = {1{`RANDOM}};
  enq_buffer_7_val_mask_1 = _RAND_3133[0:0];
  _RAND_3134 = {1{`RANDOM}};
  enq_buffer_7_val_mask_2 = _RAND_3134[0:0];
  _RAND_3135 = {1{`RANDOM}};
  enq_buffer_7_val_mask_3 = _RAND_3135[0:0];
  _RAND_3136 = {1{`RANDOM}};
  enq_valid = _RAND_3136[0:0];
  _RAND_3137 = {1{`RANDOM}};
  set_idx = _RAND_3137[4:0];
  _RAND_3138 = {1{`RANDOM}};
  set_num = _RAND_3138[4:0];
  _RAND_3139 = {1{`RANDOM}};
  REG = _RAND_3139[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
