module BundleBridgeNexus_12(
  input   clock,
  input   reset
);
endmodule
