module ForwardingAgeLogic(
  input         clock,
  input         reset,
  input  [15:0] io_addr_matches,
  input  [3:0]  io_youngest_st_idx,
  output        io_forwarding_val,
  output [3:0]  io_forwarding_idx
);
  wire  _T = 4'h0 >= io_youngest_st_idx; // @[lsu.scala 1691:17]
  wire  age_mask_0 = _T ? 1'h0 : 1'h1; // @[lsu.scala 1692:7 lsu.scala 1693:22 lsu.scala 1690:19]
  wire  _T_1 = 4'h1 >= io_youngest_st_idx; // @[lsu.scala 1691:17]
  wire  age_mask_1 = _T_1 ? 1'h0 : 1'h1; // @[lsu.scala 1692:7 lsu.scala 1693:22 lsu.scala 1690:19]
  wire  _T_2 = 4'h2 >= io_youngest_st_idx; // @[lsu.scala 1691:17]
  wire  age_mask_2 = _T_2 ? 1'h0 : 1'h1; // @[lsu.scala 1692:7 lsu.scala 1693:22 lsu.scala 1690:19]
  wire  _T_3 = 4'h3 >= io_youngest_st_idx; // @[lsu.scala 1691:17]
  wire  age_mask_3 = _T_3 ? 1'h0 : 1'h1; // @[lsu.scala 1692:7 lsu.scala 1693:22 lsu.scala 1690:19]
  wire  _T_4 = 4'h4 >= io_youngest_st_idx; // @[lsu.scala 1691:17]
  wire  age_mask_4 = _T_4 ? 1'h0 : 1'h1; // @[lsu.scala 1692:7 lsu.scala 1693:22 lsu.scala 1690:19]
  wire  _T_5 = 4'h5 >= io_youngest_st_idx; // @[lsu.scala 1691:17]
  wire  age_mask_5 = _T_5 ? 1'h0 : 1'h1; // @[lsu.scala 1692:7 lsu.scala 1693:22 lsu.scala 1690:19]
  wire  _T_6 = 4'h6 >= io_youngest_st_idx; // @[lsu.scala 1691:17]
  wire  age_mask_6 = _T_6 ? 1'h0 : 1'h1; // @[lsu.scala 1692:7 lsu.scala 1693:22 lsu.scala 1690:19]
  wire  _T_7 = 4'h7 >= io_youngest_st_idx; // @[lsu.scala 1691:17]
  wire  age_mask_7 = _T_7 ? 1'h0 : 1'h1; // @[lsu.scala 1692:7 lsu.scala 1693:22 lsu.scala 1690:19]
  wire  _T_8 = 4'h8 >= io_youngest_st_idx; // @[lsu.scala 1691:17]
  wire  age_mask_8 = _T_8 ? 1'h0 : 1'h1; // @[lsu.scala 1692:7 lsu.scala 1693:22 lsu.scala 1690:19]
  wire  _T_9 = 4'h9 >= io_youngest_st_idx; // @[lsu.scala 1691:17]
  wire  age_mask_9 = _T_9 ? 1'h0 : 1'h1; // @[lsu.scala 1692:7 lsu.scala 1693:22 lsu.scala 1690:19]
  wire  _T_10 = 4'ha >= io_youngest_st_idx; // @[lsu.scala 1691:17]
  wire  age_mask_10 = _T_10 ? 1'h0 : 1'h1; // @[lsu.scala 1692:7 lsu.scala 1693:22 lsu.scala 1690:19]
  wire  _T_11 = 4'hb >= io_youngest_st_idx; // @[lsu.scala 1691:17]
  wire  age_mask_11 = _T_11 ? 1'h0 : 1'h1; // @[lsu.scala 1692:7 lsu.scala 1693:22 lsu.scala 1690:19]
  wire  _T_12 = 4'hc >= io_youngest_st_idx; // @[lsu.scala 1691:17]
  wire  age_mask_12 = _T_12 ? 1'h0 : 1'h1; // @[lsu.scala 1692:7 lsu.scala 1693:22 lsu.scala 1690:19]
  wire  _T_13 = 4'hd >= io_youngest_st_idx; // @[lsu.scala 1691:17]
  wire  age_mask_13 = _T_13 ? 1'h0 : 1'h1; // @[lsu.scala 1692:7 lsu.scala 1693:22 lsu.scala 1690:19]
  wire  _T_14 = 4'he >= io_youngest_st_idx; // @[lsu.scala 1691:17]
  wire  age_mask_14 = _T_14 ? 1'h0 : 1'h1; // @[lsu.scala 1692:7 lsu.scala 1693:22 lsu.scala 1690:19]
  wire [7:0] lo = {age_mask_7,age_mask_6,age_mask_5,age_mask_4,age_mask_3,age_mask_2,age_mask_1,age_mask_0}; // @[lsu.scala 1699:46]
  wire [15:0] _T_16 = {1'h0,age_mask_14,age_mask_13,age_mask_12,age_mask_11,age_mask_10,age_mask_9,age_mask_8,lo}; // @[lsu.scala 1699:46]
  wire [15:0] hi_1 = io_addr_matches & _T_16; // @[lsu.scala 1699:35]
  wire [31:0] matches_ = {hi_1,io_addr_matches}; // @[Cat.scala 30:58]
  wire [1:0] _GEN_21 = matches_[2] ? 2'h2 : {{1'd0}, matches_[1]}; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [1:0] _GEN_23 = matches_[3] ? 2'h3 : _GEN_21; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [2:0] _GEN_25 = matches_[4] ? 3'h4 : {{1'd0}, _GEN_23}; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [2:0] _GEN_27 = matches_[5] ? 3'h5 : _GEN_25; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [2:0] _GEN_29 = matches_[6] ? 3'h6 : _GEN_27; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [2:0] _GEN_31 = matches_[7] ? 3'h7 : _GEN_29; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_33 = matches_[8] ? 4'h8 : {{1'd0}, _GEN_31}; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_35 = matches_[9] ? 4'h9 : _GEN_33; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_37 = matches_[10] ? 4'ha : _GEN_35; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_39 = matches_[11] ? 4'hb : _GEN_37; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_41 = matches_[12] ? 4'hc : _GEN_39; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_43 = matches_[13] ? 4'hd : _GEN_41; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_45 = matches_[14] ? 4'he : _GEN_43; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_47 = matches_[15] ? 4'hf : _GEN_45; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_49 = matches_[16] ? 4'h0 : _GEN_47; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_51 = matches_[17] ? 4'h1 : _GEN_49; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_53 = matches_[18] ? 4'h2 : _GEN_51; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_55 = matches_[19] ? 4'h3 : _GEN_53; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_57 = matches_[20] ? 4'h4 : _GEN_55; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_59 = matches_[21] ? 4'h5 : _GEN_57; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_61 = matches_[22] ? 4'h6 : _GEN_59; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_63 = matches_[23] ? 4'h7 : _GEN_61; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_65 = matches_[24] ? 4'h8 : _GEN_63; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_67 = matches_[25] ? 4'h9 : _GEN_65; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_69 = matches_[26] ? 4'ha : _GEN_67; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_71 = matches_[27] ? 4'hb : _GEN_69; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_73 = matches_[28] ? 4'hc : _GEN_71; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire [3:0] _GEN_75 = matches_[29] ? 4'hd : _GEN_73; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  wire  _GEN_76 = matches_[30] | (matches_[29] | (matches_[28] | (matches_[27] | (matches_[26] | (matches_[25] | (
    matches_[24] | (matches_[23] | (matches_[22] | (matches_[21] | (matches_[20] | (matches_[19] | (matches_[18] | (
    matches_[17] | (matches_[16] | (matches_[15] | (matches_[14] | (matches_[13] | (matches_[12] | (matches_[11] | (
    matches_[10] | (matches_[9] | (matches_[8] | (matches_[7] | (matches_[6] | (matches_[5] | (matches_[4] | (matches_[3
    ] | (matches_[2] | (matches_[1] | matches_[0]))))))))))))))))))))))))))))); // @[lsu.scala 1710:7 lsu.scala 1711:22]
  wire [3:0] _GEN_77 = matches_[30] ? 4'he : _GEN_75; // @[lsu.scala 1710:7 lsu.scala 1712:28]
  assign io_forwarding_val = matches_[31] | _GEN_76; // @[lsu.scala 1710:7 lsu.scala 1711:22]
  assign io_forwarding_idx = matches_[31] ? 4'hf : _GEN_77; // @[lsu.scala 1710:7 lsu.scala 1712:28]
endmodule
