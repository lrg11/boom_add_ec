module BundleBridgeNexus_16(
  input   clock,
  input   reset,
  output  auto_out
);
  assign auto_out = 1'h0; // @[HasTiles.scala 162:32]
endmodule
